magic
tech sky130A
magscale 1 2
timestamp 1745609222
<< checkpaint >>
rect -3932 -3108 10832 14396
<< viali >>
rect 4997 9129 5031 9163
rect 5365 9061 5399 9095
rect 1409 8925 1443 8959
rect 1685 8925 1719 8959
rect 3893 8925 3927 8959
rect 4077 8925 4111 8959
rect 4813 8925 4847 8959
rect 5181 8925 5215 8959
rect 1593 8789 1627 8823
rect 1869 8789 1903 8823
rect 3985 8789 4019 8823
rect 2881 8449 2915 8483
rect 3065 8449 3099 8483
rect 4353 8449 4387 8483
rect 4813 8449 4847 8483
rect 4675 8381 4709 8415
rect 4445 8313 4479 8347
rect 4537 8313 4571 8347
rect 3065 8245 3099 8279
rect 4353 7905 4387 7939
rect 1409 7837 1443 7871
rect 4445 7837 4479 7871
rect 5181 7837 5215 7871
rect 1593 7701 1627 7735
rect 4813 7701 4847 7735
rect 5365 7701 5399 7735
rect 1685 7361 1719 7395
rect 1961 7361 1995 7395
rect 2513 7361 2547 7395
rect 1777 7293 1811 7327
rect 2605 7293 2639 7327
rect 1685 7157 1719 7191
rect 2145 7157 2179 7191
rect 2881 7157 2915 7191
rect 1593 6885 1627 6919
rect 1961 6817 1995 6851
rect 1501 6749 1535 6783
rect 1685 6749 1719 6783
rect 1777 6749 1811 6783
rect 2053 6749 2087 6783
rect 5181 6749 5215 6783
rect 2237 6613 2271 6647
rect 5365 6613 5399 6647
rect 1593 6409 1627 6443
rect 1409 6273 1443 6307
rect 2697 5661 2731 5695
rect 2881 5661 2915 5695
rect 3065 5661 3099 5695
rect 5365 5661 5399 5695
rect 5181 5525 5215 5559
rect 3341 5321 3375 5355
rect 2605 5253 2639 5287
rect 1409 5185 1443 5219
rect 2513 5185 2547 5219
rect 2697 5185 2731 5219
rect 3801 5185 3835 5219
rect 5181 5185 5215 5219
rect 3525 5049 3559 5083
rect 1593 4981 1627 5015
rect 5365 4981 5399 5015
rect 3157 4641 3191 4675
rect 3065 4573 3099 4607
rect 3433 4437 3467 4471
rect 1409 4097 1443 4131
rect 1777 4097 1811 4131
rect 1869 4097 1903 4131
rect 2145 4097 2179 4131
rect 3985 4097 4019 4131
rect 4169 4097 4203 4131
rect 5181 4097 5215 4131
rect 4353 4029 4387 4063
rect 2053 3961 2087 3995
rect 1593 3893 1627 3927
rect 2329 3893 2363 3927
rect 5365 3893 5399 3927
rect 2789 3689 2823 3723
rect 3249 3689 3283 3723
rect 2973 3485 3007 3519
rect 3065 3485 3099 3519
rect 3249 3485 3283 3519
rect 3433 3145 3467 3179
rect 3341 3009 3375 3043
rect 3525 3009 3559 3043
rect 1869 2601 1903 2635
rect 1593 2533 1627 2567
rect 1409 2397 1443 2431
rect 1685 2397 1719 2431
rect 4905 2397 4939 2431
rect 5089 2397 5123 2431
rect 5457 2329 5491 2363
rect 4721 2261 4755 2295
<< metal1 >>
rect 1104 9274 5796 9296
rect 1104 9222 1950 9274
rect 2002 9222 2014 9274
rect 2066 9222 2078 9274
rect 2130 9222 2142 9274
rect 2194 9222 2206 9274
rect 2258 9222 5796 9274
rect 1104 9200 5796 9222
rect 4982 9120 4988 9172
rect 5040 9120 5046 9172
rect 5350 9052 5356 9104
rect 5408 9052 5414 9104
rect 1394 8916 1400 8968
rect 1452 8916 1458 8968
rect 1673 8959 1731 8965
rect 1673 8925 1685 8959
rect 1719 8925 1731 8959
rect 1673 8919 1731 8925
rect 842 8848 848 8900
rect 900 8888 906 8900
rect 1688 8888 1716 8919
rect 3878 8916 3884 8968
rect 3936 8916 3942 8968
rect 4062 8916 4068 8968
rect 4120 8916 4126 8968
rect 4798 8916 4804 8968
rect 4856 8916 4862 8968
rect 4982 8916 4988 8968
rect 5040 8956 5046 8968
rect 5169 8959 5227 8965
rect 5169 8956 5181 8959
rect 5040 8928 5181 8956
rect 5040 8916 5046 8928
rect 5169 8925 5181 8928
rect 5215 8925 5227 8959
rect 5169 8919 5227 8925
rect 900 8860 1716 8888
rect 900 8848 906 8860
rect 1578 8780 1584 8832
rect 1636 8780 1642 8832
rect 1854 8780 1860 8832
rect 1912 8780 1918 8832
rect 3970 8780 3976 8832
rect 4028 8780 4034 8832
rect 1104 8730 5796 8752
rect 1104 8678 2610 8730
rect 2662 8678 2674 8730
rect 2726 8678 2738 8730
rect 2790 8678 2802 8730
rect 2854 8678 2866 8730
rect 2918 8678 5796 8730
rect 1104 8656 5796 8678
rect 1578 8508 1584 8560
rect 1636 8548 1642 8560
rect 1636 8520 3096 8548
rect 1636 8508 1642 8520
rect 1854 8440 1860 8492
rect 1912 8480 1918 8492
rect 3068 8489 3096 8520
rect 4062 8508 4068 8560
rect 4120 8548 4126 8560
rect 4120 8520 4844 8548
rect 4120 8508 4126 8520
rect 2869 8483 2927 8489
rect 2869 8480 2881 8483
rect 1912 8452 2881 8480
rect 1912 8440 1918 8452
rect 2869 8449 2881 8452
rect 2915 8449 2927 8483
rect 2869 8443 2927 8449
rect 3053 8483 3111 8489
rect 3053 8449 3065 8483
rect 3099 8449 3111 8483
rect 3053 8443 3111 8449
rect 4338 8440 4344 8492
rect 4396 8440 4402 8492
rect 4816 8489 4844 8520
rect 4801 8483 4859 8489
rect 4801 8449 4813 8483
rect 4847 8449 4859 8483
rect 4801 8443 4859 8449
rect 3234 8372 3240 8424
rect 3292 8412 3298 8424
rect 4663 8415 4721 8421
rect 4663 8412 4675 8415
rect 3292 8384 4675 8412
rect 3292 8372 3298 8384
rect 4663 8381 4675 8384
rect 4709 8381 4721 8415
rect 4663 8375 4721 8381
rect 4430 8304 4436 8356
rect 4488 8304 4494 8356
rect 4525 8347 4583 8353
rect 4525 8313 4537 8347
rect 4571 8313 4583 8347
rect 4525 8307 4583 8313
rect 3050 8236 3056 8288
rect 3108 8236 3114 8288
rect 3418 8236 3424 8288
rect 3476 8276 3482 8288
rect 3878 8276 3884 8288
rect 3476 8248 3884 8276
rect 3476 8236 3482 8248
rect 3878 8236 3884 8248
rect 3936 8276 3942 8288
rect 4540 8276 4568 8307
rect 3936 8248 4568 8276
rect 3936 8236 3942 8248
rect 1104 8186 5796 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 5796 8186
rect 1104 8112 5796 8134
rect 3050 7896 3056 7948
rect 3108 7936 3114 7948
rect 3510 7936 3516 7948
rect 3108 7908 3516 7936
rect 3108 7896 3114 7908
rect 3510 7896 3516 7908
rect 3568 7936 3574 7948
rect 4341 7939 4399 7945
rect 4341 7936 4353 7939
rect 3568 7908 4353 7936
rect 3568 7896 3574 7908
rect 4341 7905 4353 7908
rect 4387 7905 4399 7939
rect 4341 7899 4399 7905
rect 842 7828 848 7880
rect 900 7868 906 7880
rect 1397 7871 1455 7877
rect 1397 7868 1409 7871
rect 900 7840 1409 7868
rect 900 7828 906 7840
rect 1397 7837 1409 7840
rect 1443 7837 1455 7871
rect 1397 7831 1455 7837
rect 4433 7871 4491 7877
rect 4433 7837 4445 7871
rect 4479 7837 4491 7871
rect 5169 7871 5227 7877
rect 5169 7868 5181 7871
rect 4433 7831 4491 7837
rect 4816 7840 5181 7868
rect 1581 7735 1639 7741
rect 1581 7701 1593 7735
rect 1627 7732 1639 7735
rect 1762 7732 1768 7744
rect 1627 7704 1768 7732
rect 1627 7701 1639 7704
rect 1581 7695 1639 7701
rect 1762 7692 1768 7704
rect 1820 7732 1826 7744
rect 4448 7732 4476 7831
rect 4816 7741 4844 7840
rect 5169 7837 5181 7840
rect 5215 7837 5227 7871
rect 5169 7831 5227 7837
rect 1820 7704 4476 7732
rect 4801 7735 4859 7741
rect 1820 7692 1826 7704
rect 4801 7701 4813 7735
rect 4847 7701 4859 7735
rect 4801 7695 4859 7701
rect 5350 7692 5356 7744
rect 5408 7692 5414 7744
rect 1104 7642 5796 7664
rect 1104 7590 2610 7642
rect 2662 7590 2674 7642
rect 2726 7590 2738 7642
rect 2790 7590 2802 7642
rect 2854 7590 2866 7642
rect 2918 7590 5796 7642
rect 1104 7568 5796 7590
rect 1486 7352 1492 7404
rect 1544 7392 1550 7404
rect 1673 7395 1731 7401
rect 1673 7392 1685 7395
rect 1544 7364 1685 7392
rect 1544 7352 1550 7364
rect 1673 7361 1685 7364
rect 1719 7361 1731 7395
rect 1673 7355 1731 7361
rect 1854 7352 1860 7404
rect 1912 7392 1918 7404
rect 1949 7395 2007 7401
rect 1949 7392 1961 7395
rect 1912 7364 1961 7392
rect 1912 7352 1918 7364
rect 1949 7361 1961 7364
rect 1995 7361 2007 7395
rect 1949 7355 2007 7361
rect 2314 7352 2320 7404
rect 2372 7392 2378 7404
rect 2501 7395 2559 7401
rect 2501 7392 2513 7395
rect 2372 7364 2513 7392
rect 2372 7352 2378 7364
rect 2501 7361 2513 7364
rect 2547 7361 2559 7395
rect 2501 7355 2559 7361
rect 1762 7284 1768 7336
rect 1820 7284 1826 7336
rect 2593 7327 2651 7333
rect 2593 7324 2605 7327
rect 2516 7296 2605 7324
rect 2516 7268 2544 7296
rect 2593 7293 2605 7296
rect 2639 7293 2651 7327
rect 2593 7287 2651 7293
rect 2498 7216 2504 7268
rect 2556 7216 2562 7268
rect 3418 7256 3424 7268
rect 2792 7228 3424 7256
rect 1578 7148 1584 7200
rect 1636 7188 1642 7200
rect 1673 7191 1731 7197
rect 1673 7188 1685 7191
rect 1636 7160 1685 7188
rect 1636 7148 1642 7160
rect 1673 7157 1685 7160
rect 1719 7157 1731 7191
rect 1673 7151 1731 7157
rect 2133 7191 2191 7197
rect 2133 7157 2145 7191
rect 2179 7188 2191 7191
rect 2792 7188 2820 7228
rect 3418 7216 3424 7228
rect 3476 7216 3482 7268
rect 2179 7160 2820 7188
rect 2869 7191 2927 7197
rect 2179 7157 2191 7160
rect 2133 7151 2191 7157
rect 2869 7157 2881 7191
rect 2915 7188 2927 7191
rect 5074 7188 5080 7200
rect 2915 7160 5080 7188
rect 2915 7157 2927 7160
rect 2869 7151 2927 7157
rect 5074 7148 5080 7160
rect 5132 7148 5138 7200
rect 1104 7098 5796 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 5796 7098
rect 1104 7024 5796 7046
rect 1581 6919 1639 6925
rect 1581 6885 1593 6919
rect 1627 6916 1639 6919
rect 1670 6916 1676 6928
rect 1627 6888 1676 6916
rect 1627 6885 1639 6888
rect 1581 6879 1639 6885
rect 1670 6876 1676 6888
rect 1728 6876 1734 6928
rect 1949 6851 2007 6857
rect 1949 6817 1961 6851
rect 1995 6848 2007 6851
rect 3786 6848 3792 6860
rect 1995 6820 3792 6848
rect 1995 6817 2007 6820
rect 1949 6811 2007 6817
rect 3786 6808 3792 6820
rect 3844 6808 3850 6860
rect 1486 6740 1492 6792
rect 1544 6740 1550 6792
rect 1578 6740 1584 6792
rect 1636 6780 1642 6792
rect 1673 6783 1731 6789
rect 1673 6780 1685 6783
rect 1636 6752 1685 6780
rect 1636 6740 1642 6752
rect 1673 6749 1685 6752
rect 1719 6749 1731 6783
rect 1673 6743 1731 6749
rect 1762 6740 1768 6792
rect 1820 6740 1826 6792
rect 2041 6783 2099 6789
rect 2041 6749 2053 6783
rect 2087 6749 2099 6783
rect 2041 6743 2099 6749
rect 5169 6783 5227 6789
rect 5169 6749 5181 6783
rect 5215 6749 5227 6783
rect 5169 6743 5227 6749
rect 2056 6712 2084 6743
rect 3326 6712 3332 6724
rect 2056 6684 3332 6712
rect 3326 6672 3332 6684
rect 3384 6672 3390 6724
rect 2225 6647 2283 6653
rect 2225 6613 2237 6647
rect 2271 6644 2283 6647
rect 5184 6644 5212 6743
rect 2271 6616 5212 6644
rect 2271 6613 2283 6616
rect 2225 6607 2283 6613
rect 5350 6604 5356 6656
rect 5408 6604 5414 6656
rect 1104 6554 5796 6576
rect 1104 6502 2610 6554
rect 2662 6502 2674 6554
rect 2726 6502 2738 6554
rect 2790 6502 2802 6554
rect 2854 6502 2866 6554
rect 2918 6502 5796 6554
rect 1104 6480 5796 6502
rect 1486 6400 1492 6452
rect 1544 6440 1550 6452
rect 1581 6443 1639 6449
rect 1581 6440 1593 6443
rect 1544 6412 1593 6440
rect 1544 6400 1550 6412
rect 1581 6409 1593 6412
rect 1627 6409 1639 6443
rect 1581 6403 1639 6409
rect 842 6264 848 6316
rect 900 6304 906 6316
rect 1397 6307 1455 6313
rect 1397 6304 1409 6307
rect 900 6276 1409 6304
rect 900 6264 906 6276
rect 1397 6273 1409 6276
rect 1443 6273 1455 6307
rect 1397 6267 1455 6273
rect 1104 6010 5796 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 5796 6010
rect 1104 5936 5796 5958
rect 4430 5760 4436 5772
rect 2884 5732 4436 5760
rect 2498 5652 2504 5704
rect 2556 5692 2562 5704
rect 2884 5701 2912 5732
rect 4430 5720 4436 5732
rect 4488 5720 4494 5772
rect 2685 5695 2743 5701
rect 2685 5692 2697 5695
rect 2556 5664 2697 5692
rect 2556 5652 2562 5664
rect 2685 5661 2697 5664
rect 2731 5661 2743 5695
rect 2685 5655 2743 5661
rect 2869 5695 2927 5701
rect 2869 5661 2881 5695
rect 2915 5661 2927 5695
rect 2869 5655 2927 5661
rect 3053 5695 3111 5701
rect 3053 5661 3065 5695
rect 3099 5692 3111 5695
rect 5353 5695 5411 5701
rect 5353 5692 5365 5695
rect 3099 5664 5365 5692
rect 3099 5661 3111 5664
rect 3053 5655 3111 5661
rect 5353 5661 5365 5664
rect 5399 5661 5411 5695
rect 5353 5655 5411 5661
rect 4890 5516 4896 5568
rect 4948 5556 4954 5568
rect 5169 5559 5227 5565
rect 5169 5556 5181 5559
rect 4948 5528 5181 5556
rect 4948 5516 4954 5528
rect 5169 5525 5181 5528
rect 5215 5525 5227 5559
rect 5169 5519 5227 5525
rect 1104 5466 5796 5488
rect 1104 5414 2610 5466
rect 2662 5414 2674 5466
rect 2726 5414 2738 5466
rect 2790 5414 2802 5466
rect 2854 5414 2866 5466
rect 2918 5414 5796 5466
rect 1104 5392 5796 5414
rect 3326 5312 3332 5364
rect 3384 5312 3390 5364
rect 3418 5312 3424 5364
rect 3476 5352 3482 5364
rect 3602 5352 3608 5364
rect 3476 5324 3608 5352
rect 3476 5312 3482 5324
rect 3602 5312 3608 5324
rect 3660 5312 3666 5364
rect 2593 5287 2651 5293
rect 2593 5253 2605 5287
rect 2639 5284 2651 5287
rect 2639 5256 5212 5284
rect 2639 5253 2651 5256
rect 2593 5247 2651 5253
rect 842 5176 848 5228
rect 900 5216 906 5228
rect 1397 5219 1455 5225
rect 1397 5216 1409 5219
rect 900 5188 1409 5216
rect 900 5176 906 5188
rect 1397 5185 1409 5188
rect 1443 5185 1455 5219
rect 1397 5179 1455 5185
rect 2501 5219 2559 5225
rect 2501 5185 2513 5219
rect 2547 5185 2559 5219
rect 2501 5179 2559 5185
rect 2685 5219 2743 5225
rect 2685 5185 2697 5219
rect 2731 5216 2743 5219
rect 3418 5216 3424 5228
rect 2731 5188 3424 5216
rect 2731 5185 2743 5188
rect 2685 5179 2743 5185
rect 2516 5148 2544 5179
rect 3418 5176 3424 5188
rect 3476 5176 3482 5228
rect 3786 5176 3792 5228
rect 3844 5176 3850 5228
rect 5184 5225 5212 5256
rect 5169 5219 5227 5225
rect 5169 5185 5181 5219
rect 5215 5185 5227 5219
rect 5169 5179 5227 5185
rect 3970 5148 3976 5160
rect 2516 5120 3976 5148
rect 3970 5108 3976 5120
rect 4028 5108 4034 5160
rect 3513 5083 3571 5089
rect 3513 5049 3525 5083
rect 3559 5080 3571 5083
rect 3602 5080 3608 5092
rect 3559 5052 3608 5080
rect 3559 5049 3571 5052
rect 3513 5043 3571 5049
rect 3602 5040 3608 5052
rect 3660 5040 3666 5092
rect 1581 5015 1639 5021
rect 1581 4981 1593 5015
rect 1627 5012 1639 5015
rect 4062 5012 4068 5024
rect 1627 4984 4068 5012
rect 1627 4981 1639 4984
rect 1581 4975 1639 4981
rect 4062 4972 4068 4984
rect 4120 4972 4126 5024
rect 5350 4972 5356 5024
rect 5408 4972 5414 5024
rect 1104 4922 5796 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 5796 4922
rect 1104 4848 5796 4870
rect 3145 4675 3203 4681
rect 3145 4641 3157 4675
rect 3191 4672 3203 4675
rect 3970 4672 3976 4684
rect 3191 4644 3976 4672
rect 3191 4641 3203 4644
rect 3145 4635 3203 4641
rect 3970 4632 3976 4644
rect 4028 4632 4034 4684
rect 3053 4607 3111 4613
rect 3053 4573 3065 4607
rect 3099 4604 3111 4607
rect 3234 4604 3240 4616
rect 3099 4576 3240 4604
rect 3099 4573 3111 4576
rect 3053 4567 3111 4573
rect 3234 4564 3240 4576
rect 3292 4564 3298 4616
rect 3421 4471 3479 4477
rect 3421 4437 3433 4471
rect 3467 4468 3479 4471
rect 5166 4468 5172 4480
rect 3467 4440 5172 4468
rect 3467 4437 3479 4440
rect 3421 4431 3479 4437
rect 5166 4428 5172 4440
rect 5224 4428 5230 4480
rect 1104 4378 5796 4400
rect 1104 4326 2610 4378
rect 2662 4326 2674 4378
rect 2726 4326 2738 4378
rect 2790 4326 2802 4378
rect 2854 4326 2866 4378
rect 2918 4326 5796 4378
rect 1104 4304 5796 4326
rect 3602 4156 3608 4208
rect 3660 4196 3666 4208
rect 3660 4168 4108 4196
rect 3660 4156 3666 4168
rect 842 4088 848 4140
rect 900 4128 906 4140
rect 1397 4131 1455 4137
rect 1397 4128 1409 4131
rect 900 4100 1409 4128
rect 900 4088 906 4100
rect 1397 4097 1409 4100
rect 1443 4097 1455 4131
rect 1397 4091 1455 4097
rect 1762 4088 1768 4140
rect 1820 4088 1826 4140
rect 1857 4131 1915 4137
rect 1857 4097 1869 4131
rect 1903 4128 1915 4131
rect 2133 4131 2191 4137
rect 2133 4128 2145 4131
rect 1903 4100 2145 4128
rect 1903 4097 1915 4100
rect 1857 4091 1915 4097
rect 2133 4097 2145 4100
rect 2179 4097 2191 4131
rect 2133 4091 2191 4097
rect 1578 4020 1584 4072
rect 1636 4060 1642 4072
rect 1872 4060 1900 4091
rect 3418 4088 3424 4140
rect 3476 4128 3482 4140
rect 3973 4131 4031 4137
rect 3973 4128 3985 4131
rect 3476 4100 3985 4128
rect 3476 4088 3482 4100
rect 3973 4097 3985 4100
rect 4019 4097 4031 4131
rect 4080 4128 4108 4168
rect 4157 4131 4215 4137
rect 4157 4128 4169 4131
rect 4080 4100 4169 4128
rect 3973 4091 4031 4097
rect 4157 4097 4169 4100
rect 4203 4097 4215 4131
rect 4157 4091 4215 4097
rect 5166 4088 5172 4140
rect 5224 4088 5230 4140
rect 3234 4060 3240 4072
rect 1636 4032 1900 4060
rect 1964 4032 3240 4060
rect 1636 4020 1642 4032
rect 1581 3927 1639 3933
rect 1581 3893 1593 3927
rect 1627 3924 1639 3927
rect 1964 3924 1992 4032
rect 3234 4020 3240 4032
rect 3292 4020 3298 4072
rect 4062 4020 4068 4072
rect 4120 4060 4126 4072
rect 4341 4063 4399 4069
rect 4341 4060 4353 4063
rect 4120 4032 4353 4060
rect 4120 4020 4126 4032
rect 4341 4029 4353 4032
rect 4387 4029 4399 4063
rect 4341 4023 4399 4029
rect 2041 3995 2099 4001
rect 2041 3961 2053 3995
rect 2087 3992 2099 3995
rect 3326 3992 3332 4004
rect 2087 3964 3332 3992
rect 2087 3961 2099 3964
rect 2041 3955 2099 3961
rect 3326 3952 3332 3964
rect 3384 3952 3390 4004
rect 1627 3896 1992 3924
rect 2317 3927 2375 3933
rect 1627 3893 1639 3896
rect 1581 3887 1639 3893
rect 2317 3893 2329 3927
rect 2363 3924 2375 3927
rect 4798 3924 4804 3936
rect 2363 3896 4804 3924
rect 2363 3893 2375 3896
rect 2317 3887 2375 3893
rect 4798 3884 4804 3896
rect 4856 3884 4862 3936
rect 5350 3884 5356 3936
rect 5408 3884 5414 3936
rect 1104 3834 5796 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 5796 3834
rect 1104 3760 5796 3782
rect 2498 3680 2504 3732
rect 2556 3720 2562 3732
rect 2777 3723 2835 3729
rect 2777 3720 2789 3723
rect 2556 3692 2789 3720
rect 2556 3680 2562 3692
rect 2777 3689 2789 3692
rect 2823 3689 2835 3723
rect 2777 3683 2835 3689
rect 3234 3680 3240 3732
rect 3292 3680 3298 3732
rect 4062 3584 4068 3596
rect 2976 3556 4068 3584
rect 2976 3525 3004 3556
rect 4062 3544 4068 3556
rect 4120 3544 4126 3596
rect 2961 3519 3019 3525
rect 2961 3485 2973 3519
rect 3007 3485 3019 3519
rect 2961 3479 3019 3485
rect 3050 3476 3056 3528
rect 3108 3516 3114 3528
rect 3237 3519 3295 3525
rect 3108 3488 3188 3516
rect 3108 3476 3114 3488
rect 3160 3448 3188 3488
rect 3237 3485 3249 3519
rect 3283 3516 3295 3519
rect 3602 3516 3608 3528
rect 3283 3488 3608 3516
rect 3283 3485 3295 3488
rect 3237 3479 3295 3485
rect 3602 3476 3608 3488
rect 3660 3476 3666 3528
rect 4338 3448 4344 3460
rect 3160 3420 4344 3448
rect 4338 3408 4344 3420
rect 4396 3408 4402 3460
rect 1104 3290 5796 3312
rect 1104 3238 2610 3290
rect 2662 3238 2674 3290
rect 2726 3238 2738 3290
rect 2790 3238 2802 3290
rect 2854 3238 2866 3290
rect 2918 3238 5796 3290
rect 1104 3216 5796 3238
rect 3421 3179 3479 3185
rect 3421 3145 3433 3179
rect 3467 3176 3479 3179
rect 4982 3176 4988 3188
rect 3467 3148 4988 3176
rect 3467 3145 3479 3148
rect 3421 3139 3479 3145
rect 4982 3136 4988 3148
rect 5040 3136 5046 3188
rect 3326 3000 3332 3052
rect 3384 3000 3390 3052
rect 3510 3000 3516 3052
rect 3568 3000 3574 3052
rect 1104 2746 5796 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 5796 2746
rect 1104 2672 5796 2694
rect 1857 2635 1915 2641
rect 1857 2601 1869 2635
rect 1903 2632 1915 2635
rect 2314 2632 2320 2644
rect 1903 2604 2320 2632
rect 1903 2601 1915 2604
rect 1857 2595 1915 2601
rect 2314 2592 2320 2604
rect 2372 2592 2378 2644
rect 1581 2567 1639 2573
rect 1581 2533 1593 2567
rect 1627 2564 1639 2567
rect 3050 2564 3056 2576
rect 1627 2536 3056 2564
rect 1627 2533 1639 2536
rect 1581 2527 1639 2533
rect 3050 2524 3056 2536
rect 3108 2524 3114 2576
rect 842 2388 848 2440
rect 900 2428 906 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 900 2400 1409 2428
rect 900 2388 906 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 1670 2388 1676 2440
rect 1728 2388 1734 2440
rect 4890 2388 4896 2440
rect 4948 2388 4954 2440
rect 5074 2388 5080 2440
rect 5132 2388 5138 2440
rect 5442 2320 5448 2372
rect 5500 2320 5506 2372
rect 4706 2252 4712 2304
rect 4764 2252 4770 2304
rect 1104 2202 5796 2224
rect 1104 2150 2610 2202
rect 2662 2150 2674 2202
rect 2726 2150 2738 2202
rect 2790 2150 2802 2202
rect 2854 2150 2866 2202
rect 2918 2150 5796 2202
rect 1104 2128 5796 2150
<< via1 >>
rect 1950 9222 2002 9274
rect 2014 9222 2066 9274
rect 2078 9222 2130 9274
rect 2142 9222 2194 9274
rect 2206 9222 2258 9274
rect 4988 9163 5040 9172
rect 4988 9129 4997 9163
rect 4997 9129 5031 9163
rect 5031 9129 5040 9163
rect 4988 9120 5040 9129
rect 5356 9095 5408 9104
rect 5356 9061 5365 9095
rect 5365 9061 5399 9095
rect 5399 9061 5408 9095
rect 5356 9052 5408 9061
rect 1400 8959 1452 8968
rect 1400 8925 1409 8959
rect 1409 8925 1443 8959
rect 1443 8925 1452 8959
rect 1400 8916 1452 8925
rect 848 8848 900 8900
rect 3884 8959 3936 8968
rect 3884 8925 3893 8959
rect 3893 8925 3927 8959
rect 3927 8925 3936 8959
rect 3884 8916 3936 8925
rect 4068 8959 4120 8968
rect 4068 8925 4077 8959
rect 4077 8925 4111 8959
rect 4111 8925 4120 8959
rect 4068 8916 4120 8925
rect 4804 8959 4856 8968
rect 4804 8925 4813 8959
rect 4813 8925 4847 8959
rect 4847 8925 4856 8959
rect 4804 8916 4856 8925
rect 4988 8916 5040 8968
rect 1584 8823 1636 8832
rect 1584 8789 1593 8823
rect 1593 8789 1627 8823
rect 1627 8789 1636 8823
rect 1584 8780 1636 8789
rect 1860 8823 1912 8832
rect 1860 8789 1869 8823
rect 1869 8789 1903 8823
rect 1903 8789 1912 8823
rect 1860 8780 1912 8789
rect 3976 8823 4028 8832
rect 3976 8789 3985 8823
rect 3985 8789 4019 8823
rect 4019 8789 4028 8823
rect 3976 8780 4028 8789
rect 2610 8678 2662 8730
rect 2674 8678 2726 8730
rect 2738 8678 2790 8730
rect 2802 8678 2854 8730
rect 2866 8678 2918 8730
rect 1584 8508 1636 8560
rect 1860 8440 1912 8492
rect 4068 8508 4120 8560
rect 4344 8483 4396 8492
rect 4344 8449 4353 8483
rect 4353 8449 4387 8483
rect 4387 8449 4396 8483
rect 4344 8440 4396 8449
rect 3240 8372 3292 8424
rect 4436 8347 4488 8356
rect 4436 8313 4445 8347
rect 4445 8313 4479 8347
rect 4479 8313 4488 8347
rect 4436 8304 4488 8313
rect 3056 8279 3108 8288
rect 3056 8245 3065 8279
rect 3065 8245 3099 8279
rect 3099 8245 3108 8279
rect 3056 8236 3108 8245
rect 3424 8236 3476 8288
rect 3884 8236 3936 8288
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 3056 7896 3108 7948
rect 3516 7896 3568 7948
rect 848 7828 900 7880
rect 1768 7692 1820 7744
rect 5356 7735 5408 7744
rect 5356 7701 5365 7735
rect 5365 7701 5399 7735
rect 5399 7701 5408 7735
rect 5356 7692 5408 7701
rect 2610 7590 2662 7642
rect 2674 7590 2726 7642
rect 2738 7590 2790 7642
rect 2802 7590 2854 7642
rect 2866 7590 2918 7642
rect 1492 7352 1544 7404
rect 1860 7352 1912 7404
rect 2320 7352 2372 7404
rect 1768 7327 1820 7336
rect 1768 7293 1777 7327
rect 1777 7293 1811 7327
rect 1811 7293 1820 7327
rect 1768 7284 1820 7293
rect 2504 7216 2556 7268
rect 1584 7148 1636 7200
rect 3424 7216 3476 7268
rect 5080 7148 5132 7200
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 1676 6876 1728 6928
rect 3792 6808 3844 6860
rect 1492 6783 1544 6792
rect 1492 6749 1501 6783
rect 1501 6749 1535 6783
rect 1535 6749 1544 6783
rect 1492 6740 1544 6749
rect 1584 6740 1636 6792
rect 1768 6783 1820 6792
rect 1768 6749 1777 6783
rect 1777 6749 1811 6783
rect 1811 6749 1820 6783
rect 1768 6740 1820 6749
rect 3332 6672 3384 6724
rect 5356 6647 5408 6656
rect 5356 6613 5365 6647
rect 5365 6613 5399 6647
rect 5399 6613 5408 6647
rect 5356 6604 5408 6613
rect 2610 6502 2662 6554
rect 2674 6502 2726 6554
rect 2738 6502 2790 6554
rect 2802 6502 2854 6554
rect 2866 6502 2918 6554
rect 1492 6400 1544 6452
rect 848 6264 900 6316
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 2504 5652 2556 5704
rect 4436 5720 4488 5772
rect 4896 5516 4948 5568
rect 2610 5414 2662 5466
rect 2674 5414 2726 5466
rect 2738 5414 2790 5466
rect 2802 5414 2854 5466
rect 2866 5414 2918 5466
rect 3332 5355 3384 5364
rect 3332 5321 3341 5355
rect 3341 5321 3375 5355
rect 3375 5321 3384 5355
rect 3332 5312 3384 5321
rect 3424 5312 3476 5364
rect 3608 5312 3660 5364
rect 848 5176 900 5228
rect 3424 5176 3476 5228
rect 3792 5219 3844 5228
rect 3792 5185 3801 5219
rect 3801 5185 3835 5219
rect 3835 5185 3844 5219
rect 3792 5176 3844 5185
rect 3976 5108 4028 5160
rect 3608 5040 3660 5092
rect 4068 4972 4120 5024
rect 5356 5015 5408 5024
rect 5356 4981 5365 5015
rect 5365 4981 5399 5015
rect 5399 4981 5408 5015
rect 5356 4972 5408 4981
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 3976 4632 4028 4684
rect 3240 4564 3292 4616
rect 5172 4428 5224 4480
rect 2610 4326 2662 4378
rect 2674 4326 2726 4378
rect 2738 4326 2790 4378
rect 2802 4326 2854 4378
rect 2866 4326 2918 4378
rect 3608 4156 3660 4208
rect 848 4088 900 4140
rect 1768 4131 1820 4140
rect 1768 4097 1777 4131
rect 1777 4097 1811 4131
rect 1811 4097 1820 4131
rect 1768 4088 1820 4097
rect 1584 4020 1636 4072
rect 3424 4088 3476 4140
rect 5172 4131 5224 4140
rect 5172 4097 5181 4131
rect 5181 4097 5215 4131
rect 5215 4097 5224 4131
rect 5172 4088 5224 4097
rect 3240 4020 3292 4072
rect 4068 4020 4120 4072
rect 3332 3952 3384 4004
rect 4804 3884 4856 3936
rect 5356 3927 5408 3936
rect 5356 3893 5365 3927
rect 5365 3893 5399 3927
rect 5399 3893 5408 3927
rect 5356 3884 5408 3893
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 2504 3680 2556 3732
rect 3240 3723 3292 3732
rect 3240 3689 3249 3723
rect 3249 3689 3283 3723
rect 3283 3689 3292 3723
rect 3240 3680 3292 3689
rect 4068 3544 4120 3596
rect 3056 3519 3108 3528
rect 3056 3485 3065 3519
rect 3065 3485 3099 3519
rect 3099 3485 3108 3519
rect 3056 3476 3108 3485
rect 3608 3476 3660 3528
rect 4344 3408 4396 3460
rect 2610 3238 2662 3290
rect 2674 3238 2726 3290
rect 2738 3238 2790 3290
rect 2802 3238 2854 3290
rect 2866 3238 2918 3290
rect 4988 3136 5040 3188
rect 3332 3043 3384 3052
rect 3332 3009 3341 3043
rect 3341 3009 3375 3043
rect 3375 3009 3384 3043
rect 3332 3000 3384 3009
rect 3516 3043 3568 3052
rect 3516 3009 3525 3043
rect 3525 3009 3559 3043
rect 3559 3009 3568 3043
rect 3516 3000 3568 3009
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 2320 2592 2372 2644
rect 3056 2524 3108 2576
rect 848 2388 900 2440
rect 1676 2431 1728 2440
rect 1676 2397 1685 2431
rect 1685 2397 1719 2431
rect 1719 2397 1728 2431
rect 1676 2388 1728 2397
rect 4896 2431 4948 2440
rect 4896 2397 4905 2431
rect 4905 2397 4939 2431
rect 4939 2397 4948 2431
rect 4896 2388 4948 2397
rect 5080 2431 5132 2440
rect 5080 2397 5089 2431
rect 5089 2397 5123 2431
rect 5123 2397 5132 2431
rect 5080 2388 5132 2397
rect 5448 2363 5500 2372
rect 5448 2329 5457 2363
rect 5457 2329 5491 2363
rect 5491 2329 5500 2363
rect 5448 2320 5500 2329
rect 4712 2295 4764 2304
rect 4712 2261 4721 2295
rect 4721 2261 4755 2295
rect 4755 2261 4764 2295
rect 4712 2252 4764 2261
rect 2610 2150 2662 2202
rect 2674 2150 2726 2202
rect 2738 2150 2790 2202
rect 2802 2150 2854 2202
rect 2866 2150 2918 2202
<< metal2 >>
rect 1398 10432 1454 10441
rect 1398 10367 1454 10376
rect 4986 10432 5042 10441
rect 4986 10367 5042 10376
rect 1412 8974 1440 10367
rect 1950 9276 2258 9285
rect 1950 9274 1956 9276
rect 2012 9274 2036 9276
rect 2092 9274 2116 9276
rect 2172 9274 2196 9276
rect 2252 9274 2258 9276
rect 2012 9222 2014 9274
rect 2194 9222 2196 9274
rect 1950 9220 1956 9222
rect 2012 9220 2036 9222
rect 2092 9220 2116 9222
rect 2172 9220 2196 9222
rect 2252 9220 2258 9222
rect 1950 9211 2258 9220
rect 5000 9178 5028 10367
rect 4988 9172 5040 9178
rect 4988 9114 5040 9120
rect 5356 9104 5408 9110
rect 5354 9072 5356 9081
rect 5408 9072 5410 9081
rect 5354 9007 5410 9016
rect 1400 8968 1452 8974
rect 846 8936 902 8945
rect 1400 8910 1452 8916
rect 3884 8968 3936 8974
rect 3884 8910 3936 8916
rect 4068 8968 4120 8974
rect 4068 8910 4120 8916
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 4988 8968 5040 8974
rect 4988 8910 5040 8916
rect 846 8871 848 8880
rect 900 8871 902 8880
rect 848 8842 900 8848
rect 1584 8832 1636 8838
rect 1584 8774 1636 8780
rect 1860 8832 1912 8838
rect 1860 8774 1912 8780
rect 1596 8566 1624 8774
rect 1584 8560 1636 8566
rect 1584 8502 1636 8508
rect 848 7880 900 7886
rect 846 7848 848 7857
rect 900 7848 902 7857
rect 846 7783 902 7792
rect 1492 7404 1544 7410
rect 1492 7346 1544 7352
rect 1504 6798 1532 7346
rect 1596 7206 1624 8502
rect 1872 8498 1900 8774
rect 2610 8732 2918 8741
rect 2610 8730 2616 8732
rect 2672 8730 2696 8732
rect 2752 8730 2776 8732
rect 2832 8730 2856 8732
rect 2912 8730 2918 8732
rect 2672 8678 2674 8730
rect 2854 8678 2856 8730
rect 2610 8676 2616 8678
rect 2672 8676 2696 8678
rect 2752 8676 2776 8678
rect 2832 8676 2856 8678
rect 2912 8676 2918 8678
rect 2610 8667 2918 8676
rect 1860 8492 1912 8498
rect 1860 8434 1912 8440
rect 1768 7744 1820 7750
rect 1768 7686 1820 7692
rect 1780 7342 1808 7686
rect 1872 7410 1900 8434
rect 3240 8424 3292 8430
rect 3240 8366 3292 8372
rect 3056 8288 3108 8294
rect 3056 8230 3108 8236
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 3068 7954 3096 8230
rect 3056 7948 3108 7954
rect 3056 7890 3108 7896
rect 2610 7644 2918 7653
rect 2610 7642 2616 7644
rect 2672 7642 2696 7644
rect 2752 7642 2776 7644
rect 2832 7642 2856 7644
rect 2912 7642 2918 7644
rect 2672 7590 2674 7642
rect 2854 7590 2856 7642
rect 2610 7588 2616 7590
rect 2672 7588 2696 7590
rect 2752 7588 2776 7590
rect 2832 7588 2856 7590
rect 2912 7588 2918 7590
rect 2610 7579 2918 7588
rect 1860 7404 1912 7410
rect 1860 7346 1912 7352
rect 2320 7404 2372 7410
rect 2320 7346 2372 7352
rect 1768 7336 1820 7342
rect 1768 7278 1820 7284
rect 1584 7200 1636 7206
rect 1584 7142 1636 7148
rect 1596 6798 1624 7142
rect 1780 7018 1808 7278
rect 1688 6990 1808 7018
rect 1688 6934 1716 6990
rect 1676 6928 1728 6934
rect 1872 6914 1900 7346
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 1676 6870 1728 6876
rect 1780 6886 1900 6914
rect 1780 6798 1808 6886
rect 1492 6792 1544 6798
rect 1492 6734 1544 6740
rect 1584 6792 1636 6798
rect 1584 6734 1636 6740
rect 1768 6792 1820 6798
rect 1768 6734 1820 6740
rect 1504 6458 1532 6734
rect 1492 6452 1544 6458
rect 1492 6394 1544 6400
rect 848 6316 900 6322
rect 848 6258 900 6264
rect 860 6225 888 6258
rect 846 6216 902 6225
rect 846 6151 902 6160
rect 848 5228 900 5234
rect 848 5170 900 5176
rect 860 5137 888 5170
rect 846 5128 902 5137
rect 846 5063 902 5072
rect 848 4140 900 4146
rect 848 4082 900 4088
rect 860 3777 888 4082
rect 1596 4078 1624 6734
rect 1780 4146 1808 6734
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 1768 4140 1820 4146
rect 1768 4082 1820 4088
rect 1584 4072 1636 4078
rect 1584 4014 1636 4020
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 846 3768 902 3777
rect 1950 3771 2258 3780
rect 846 3703 902 3712
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 2332 2650 2360 7346
rect 2504 7268 2556 7274
rect 2504 7210 2556 7216
rect 2516 5710 2544 7210
rect 2610 6556 2918 6565
rect 2610 6554 2616 6556
rect 2672 6554 2696 6556
rect 2752 6554 2776 6556
rect 2832 6554 2856 6556
rect 2912 6554 2918 6556
rect 2672 6502 2674 6554
rect 2854 6502 2856 6554
rect 2610 6500 2616 6502
rect 2672 6500 2696 6502
rect 2752 6500 2776 6502
rect 2832 6500 2856 6502
rect 2912 6500 2918 6502
rect 2610 6491 2918 6500
rect 2504 5704 2556 5710
rect 2504 5646 2556 5652
rect 2516 3738 2544 5646
rect 2610 5468 2918 5477
rect 2610 5466 2616 5468
rect 2672 5466 2696 5468
rect 2752 5466 2776 5468
rect 2832 5466 2856 5468
rect 2912 5466 2918 5468
rect 2672 5414 2674 5466
rect 2854 5414 2856 5466
rect 2610 5412 2616 5414
rect 2672 5412 2696 5414
rect 2752 5412 2776 5414
rect 2832 5412 2856 5414
rect 2912 5412 2918 5414
rect 2610 5403 2918 5412
rect 3252 4622 3280 8366
rect 3896 8294 3924 8910
rect 3976 8832 4028 8838
rect 3976 8774 4028 8780
rect 3424 8288 3476 8294
rect 3424 8230 3476 8236
rect 3884 8288 3936 8294
rect 3884 8230 3936 8236
rect 3436 7274 3464 8230
rect 3516 7948 3568 7954
rect 3516 7890 3568 7896
rect 3424 7268 3476 7274
rect 3424 7210 3476 7216
rect 3332 6724 3384 6730
rect 3332 6666 3384 6672
rect 3344 5370 3372 6666
rect 3436 5370 3464 7210
rect 3332 5364 3384 5370
rect 3332 5306 3384 5312
rect 3424 5364 3476 5370
rect 3424 5306 3476 5312
rect 3424 5228 3476 5234
rect 3424 5170 3476 5176
rect 3240 4616 3292 4622
rect 3240 4558 3292 4564
rect 2610 4380 2918 4389
rect 2610 4378 2616 4380
rect 2672 4378 2696 4380
rect 2752 4378 2776 4380
rect 2832 4378 2856 4380
rect 2912 4378 2918 4380
rect 2672 4326 2674 4378
rect 2854 4326 2856 4378
rect 2610 4324 2616 4326
rect 2672 4324 2696 4326
rect 2752 4324 2776 4326
rect 2832 4324 2856 4326
rect 2912 4324 2918 4326
rect 2610 4315 2918 4324
rect 3252 4078 3280 4558
rect 3436 4146 3464 5170
rect 3424 4140 3476 4146
rect 3424 4082 3476 4088
rect 3240 4072 3292 4078
rect 3240 4014 3292 4020
rect 3252 3738 3280 4014
rect 3332 4004 3384 4010
rect 3332 3946 3384 3952
rect 2504 3732 2556 3738
rect 2504 3674 2556 3680
rect 3240 3732 3292 3738
rect 3240 3674 3292 3680
rect 3056 3528 3108 3534
rect 3056 3470 3108 3476
rect 2610 3292 2918 3301
rect 2610 3290 2616 3292
rect 2672 3290 2696 3292
rect 2752 3290 2776 3292
rect 2832 3290 2856 3292
rect 2912 3290 2918 3292
rect 2672 3238 2674 3290
rect 2854 3238 2856 3290
rect 2610 3236 2616 3238
rect 2672 3236 2696 3238
rect 2752 3236 2776 3238
rect 2832 3236 2856 3238
rect 2912 3236 2918 3238
rect 2610 3227 2918 3236
rect 2320 2644 2372 2650
rect 2320 2586 2372 2592
rect 3068 2582 3096 3470
rect 3344 3058 3372 3946
rect 3528 3058 3556 7890
rect 3792 6860 3844 6866
rect 3792 6802 3844 6808
rect 3608 5364 3660 5370
rect 3608 5306 3660 5312
rect 3620 5098 3648 5306
rect 3804 5234 3832 6802
rect 3792 5228 3844 5234
rect 3792 5170 3844 5176
rect 3988 5166 4016 8774
rect 4080 8566 4108 8910
rect 4068 8560 4120 8566
rect 4068 8502 4120 8508
rect 3976 5160 4028 5166
rect 3976 5102 4028 5108
rect 3608 5092 3660 5098
rect 3608 5034 3660 5040
rect 3620 4214 3648 5034
rect 3988 4690 4016 5102
rect 4080 5030 4108 8502
rect 4344 8492 4396 8498
rect 4344 8434 4396 8440
rect 4068 5024 4120 5030
rect 4068 4966 4120 4972
rect 3976 4684 4028 4690
rect 3976 4626 4028 4632
rect 3608 4208 3660 4214
rect 3608 4150 3660 4156
rect 3620 3534 3648 4150
rect 4080 4078 4108 4966
rect 4068 4072 4120 4078
rect 4068 4014 4120 4020
rect 4080 3602 4108 4014
rect 4068 3596 4120 3602
rect 4068 3538 4120 3544
rect 3608 3528 3660 3534
rect 3608 3470 3660 3476
rect 4356 3466 4384 8434
rect 4436 8356 4488 8362
rect 4436 8298 4488 8304
rect 4448 5778 4476 8298
rect 4436 5772 4488 5778
rect 4436 5714 4488 5720
rect 4816 3942 4844 8910
rect 4896 5568 4948 5574
rect 4896 5510 4948 5516
rect 4804 3936 4856 3942
rect 4804 3878 4856 3884
rect 4344 3460 4396 3466
rect 4344 3402 4396 3408
rect 3332 3052 3384 3058
rect 3332 2994 3384 3000
rect 3516 3052 3568 3058
rect 3516 2994 3568 3000
rect 3056 2576 3108 2582
rect 3056 2518 3108 2524
rect 4908 2446 4936 5510
rect 5000 3194 5028 8910
rect 5356 7744 5408 7750
rect 5354 7712 5356 7721
rect 5408 7712 5410 7721
rect 5354 7647 5410 7656
rect 5080 7200 5132 7206
rect 5080 7142 5132 7148
rect 4988 3188 5040 3194
rect 4988 3130 5040 3136
rect 5092 2446 5120 7142
rect 5356 6656 5408 6662
rect 5356 6598 5408 6604
rect 5368 6361 5396 6598
rect 5354 6352 5410 6361
rect 5354 6287 5410 6296
rect 5356 5024 5408 5030
rect 5354 4992 5356 5001
rect 5408 4992 5410 5001
rect 5354 4927 5410 4936
rect 5172 4480 5224 4486
rect 5172 4422 5224 4428
rect 5184 4146 5212 4422
rect 5172 4140 5224 4146
rect 5172 4082 5224 4088
rect 5356 3936 5408 3942
rect 5356 3878 5408 3884
rect 5368 3641 5396 3878
rect 5354 3632 5410 3641
rect 5354 3567 5410 3576
rect 848 2440 900 2446
rect 846 2408 848 2417
rect 1676 2440 1728 2446
rect 900 2408 902 2417
rect 1676 2382 1728 2388
rect 4896 2440 4948 2446
rect 4896 2382 4948 2388
rect 5080 2440 5132 2446
rect 5080 2382 5132 2388
rect 846 2343 902 2352
rect 1688 921 1716 2382
rect 5448 2372 5500 2378
rect 5448 2314 5500 2320
rect 4712 2304 4764 2310
rect 4710 2272 4712 2281
rect 4764 2272 4766 2281
rect 2610 2204 2918 2213
rect 4710 2207 4766 2216
rect 2610 2202 2616 2204
rect 2672 2202 2696 2204
rect 2752 2202 2776 2204
rect 2832 2202 2856 2204
rect 2912 2202 2918 2204
rect 2672 2150 2674 2202
rect 2854 2150 2856 2202
rect 2610 2148 2616 2150
rect 2672 2148 2696 2150
rect 2752 2148 2776 2150
rect 2832 2148 2856 2150
rect 2912 2148 2918 2150
rect 2610 2139 2918 2148
rect 5460 921 5488 2314
rect 1674 912 1730 921
rect 1674 847 1730 856
rect 5446 912 5502 921
rect 5446 847 5502 856
<< via2 >>
rect 1398 10376 1454 10432
rect 4986 10376 5042 10432
rect 1956 9274 2012 9276
rect 2036 9274 2092 9276
rect 2116 9274 2172 9276
rect 2196 9274 2252 9276
rect 1956 9222 2002 9274
rect 2002 9222 2012 9274
rect 2036 9222 2066 9274
rect 2066 9222 2078 9274
rect 2078 9222 2092 9274
rect 2116 9222 2130 9274
rect 2130 9222 2142 9274
rect 2142 9222 2172 9274
rect 2196 9222 2206 9274
rect 2206 9222 2252 9274
rect 1956 9220 2012 9222
rect 2036 9220 2092 9222
rect 2116 9220 2172 9222
rect 2196 9220 2252 9222
rect 5354 9052 5356 9072
rect 5356 9052 5408 9072
rect 5408 9052 5410 9072
rect 5354 9016 5410 9052
rect 846 8900 902 8936
rect 846 8880 848 8900
rect 848 8880 900 8900
rect 900 8880 902 8900
rect 846 7828 848 7848
rect 848 7828 900 7848
rect 900 7828 902 7848
rect 846 7792 902 7828
rect 2616 8730 2672 8732
rect 2696 8730 2752 8732
rect 2776 8730 2832 8732
rect 2856 8730 2912 8732
rect 2616 8678 2662 8730
rect 2662 8678 2672 8730
rect 2696 8678 2726 8730
rect 2726 8678 2738 8730
rect 2738 8678 2752 8730
rect 2776 8678 2790 8730
rect 2790 8678 2802 8730
rect 2802 8678 2832 8730
rect 2856 8678 2866 8730
rect 2866 8678 2912 8730
rect 2616 8676 2672 8678
rect 2696 8676 2752 8678
rect 2776 8676 2832 8678
rect 2856 8676 2912 8678
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 2616 7642 2672 7644
rect 2696 7642 2752 7644
rect 2776 7642 2832 7644
rect 2856 7642 2912 7644
rect 2616 7590 2662 7642
rect 2662 7590 2672 7642
rect 2696 7590 2726 7642
rect 2726 7590 2738 7642
rect 2738 7590 2752 7642
rect 2776 7590 2790 7642
rect 2790 7590 2802 7642
rect 2802 7590 2832 7642
rect 2856 7590 2866 7642
rect 2866 7590 2912 7642
rect 2616 7588 2672 7590
rect 2696 7588 2752 7590
rect 2776 7588 2832 7590
rect 2856 7588 2912 7590
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 846 6160 902 6216
rect 846 5072 902 5128
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 846 3712 902 3768
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 2616 6554 2672 6556
rect 2696 6554 2752 6556
rect 2776 6554 2832 6556
rect 2856 6554 2912 6556
rect 2616 6502 2662 6554
rect 2662 6502 2672 6554
rect 2696 6502 2726 6554
rect 2726 6502 2738 6554
rect 2738 6502 2752 6554
rect 2776 6502 2790 6554
rect 2790 6502 2802 6554
rect 2802 6502 2832 6554
rect 2856 6502 2866 6554
rect 2866 6502 2912 6554
rect 2616 6500 2672 6502
rect 2696 6500 2752 6502
rect 2776 6500 2832 6502
rect 2856 6500 2912 6502
rect 2616 5466 2672 5468
rect 2696 5466 2752 5468
rect 2776 5466 2832 5468
rect 2856 5466 2912 5468
rect 2616 5414 2662 5466
rect 2662 5414 2672 5466
rect 2696 5414 2726 5466
rect 2726 5414 2738 5466
rect 2738 5414 2752 5466
rect 2776 5414 2790 5466
rect 2790 5414 2802 5466
rect 2802 5414 2832 5466
rect 2856 5414 2866 5466
rect 2866 5414 2912 5466
rect 2616 5412 2672 5414
rect 2696 5412 2752 5414
rect 2776 5412 2832 5414
rect 2856 5412 2912 5414
rect 2616 4378 2672 4380
rect 2696 4378 2752 4380
rect 2776 4378 2832 4380
rect 2856 4378 2912 4380
rect 2616 4326 2662 4378
rect 2662 4326 2672 4378
rect 2696 4326 2726 4378
rect 2726 4326 2738 4378
rect 2738 4326 2752 4378
rect 2776 4326 2790 4378
rect 2790 4326 2802 4378
rect 2802 4326 2832 4378
rect 2856 4326 2866 4378
rect 2866 4326 2912 4378
rect 2616 4324 2672 4326
rect 2696 4324 2752 4326
rect 2776 4324 2832 4326
rect 2856 4324 2912 4326
rect 2616 3290 2672 3292
rect 2696 3290 2752 3292
rect 2776 3290 2832 3292
rect 2856 3290 2912 3292
rect 2616 3238 2662 3290
rect 2662 3238 2672 3290
rect 2696 3238 2726 3290
rect 2726 3238 2738 3290
rect 2738 3238 2752 3290
rect 2776 3238 2790 3290
rect 2790 3238 2802 3290
rect 2802 3238 2832 3290
rect 2856 3238 2866 3290
rect 2866 3238 2912 3290
rect 2616 3236 2672 3238
rect 2696 3236 2752 3238
rect 2776 3236 2832 3238
rect 2856 3236 2912 3238
rect 5354 7692 5356 7712
rect 5356 7692 5408 7712
rect 5408 7692 5410 7712
rect 5354 7656 5410 7692
rect 5354 6296 5410 6352
rect 5354 4972 5356 4992
rect 5356 4972 5408 4992
rect 5408 4972 5410 4992
rect 5354 4936 5410 4972
rect 5354 3576 5410 3632
rect 846 2388 848 2408
rect 848 2388 900 2408
rect 900 2388 902 2408
rect 846 2352 902 2388
rect 4710 2252 4712 2272
rect 4712 2252 4764 2272
rect 4764 2252 4766 2272
rect 4710 2216 4766 2252
rect 2616 2202 2672 2204
rect 2696 2202 2752 2204
rect 2776 2202 2832 2204
rect 2856 2202 2912 2204
rect 2616 2150 2662 2202
rect 2662 2150 2672 2202
rect 2696 2150 2726 2202
rect 2726 2150 2738 2202
rect 2738 2150 2752 2202
rect 2776 2150 2790 2202
rect 2790 2150 2802 2202
rect 2802 2150 2832 2202
rect 2856 2150 2866 2202
rect 2866 2150 2912 2202
rect 2616 2148 2672 2150
rect 2696 2148 2752 2150
rect 2776 2148 2832 2150
rect 2856 2148 2912 2150
rect 1674 856 1730 912
rect 5446 856 5502 912
<< metal3 >>
rect 0 10434 800 10464
rect 1393 10434 1459 10437
rect 0 10432 1459 10434
rect 0 10376 1398 10432
rect 1454 10376 1459 10432
rect 0 10374 1459 10376
rect 0 10344 800 10374
rect 1393 10371 1459 10374
rect 4981 10434 5047 10437
rect 6100 10434 6900 10464
rect 4981 10432 6900 10434
rect 4981 10376 4986 10432
rect 5042 10376 6900 10432
rect 4981 10374 6900 10376
rect 4981 10371 5047 10374
rect 6100 10344 6900 10374
rect 1946 9280 2262 9281
rect 1946 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2262 9280
rect 1946 9215 2262 9216
rect 0 9074 800 9104
rect 5349 9074 5415 9077
rect 6100 9074 6900 9104
rect 0 8984 858 9074
rect 5349 9072 6900 9074
rect 5349 9016 5354 9072
rect 5410 9016 6900 9072
rect 5349 9014 6900 9016
rect 5349 9011 5415 9014
rect 6100 8984 6900 9014
rect 798 8941 858 8984
rect 798 8936 907 8941
rect 798 8880 846 8936
rect 902 8880 907 8936
rect 798 8878 907 8880
rect 841 8875 907 8878
rect 2606 8736 2922 8737
rect 2606 8672 2612 8736
rect 2676 8672 2692 8736
rect 2756 8672 2772 8736
rect 2836 8672 2852 8736
rect 2916 8672 2922 8736
rect 2606 8671 2922 8672
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 841 7850 907 7853
rect 798 7848 907 7850
rect 798 7792 846 7848
rect 902 7792 907 7848
rect 798 7787 907 7792
rect 798 7744 858 7787
rect 0 7654 858 7744
rect 5349 7714 5415 7717
rect 6100 7714 6900 7744
rect 5349 7712 6900 7714
rect 5349 7656 5354 7712
rect 5410 7656 6900 7712
rect 5349 7654 6900 7656
rect 0 7624 800 7654
rect 5349 7651 5415 7654
rect 2606 7648 2922 7649
rect 2606 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2922 7648
rect 6100 7624 6900 7654
rect 2606 7583 2922 7584
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 2606 6560 2922 6561
rect 2606 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2922 6560
rect 2606 6495 2922 6496
rect 0 6354 800 6384
rect 5349 6354 5415 6357
rect 6100 6354 6900 6384
rect 0 6264 858 6354
rect 5349 6352 6900 6354
rect 5349 6296 5354 6352
rect 5410 6296 6900 6352
rect 5349 6294 6900 6296
rect 5349 6291 5415 6294
rect 6100 6264 6900 6294
rect 798 6221 858 6264
rect 798 6216 907 6221
rect 798 6160 846 6216
rect 902 6160 907 6216
rect 798 6158 907 6160
rect 841 6155 907 6158
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 2606 5472 2922 5473
rect 2606 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2922 5472
rect 2606 5407 2922 5408
rect 841 5130 907 5133
rect 798 5128 907 5130
rect 798 5072 846 5128
rect 902 5072 907 5128
rect 798 5067 907 5072
rect 798 5024 858 5067
rect 0 4934 858 5024
rect 5349 4994 5415 4997
rect 6100 4994 6900 5024
rect 5349 4992 6900 4994
rect 5349 4936 5354 4992
rect 5410 4936 6900 4992
rect 5349 4934 6900 4936
rect 0 4904 800 4934
rect 5349 4931 5415 4934
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 6100 4904 6900 4934
rect 1946 4863 2262 4864
rect 2606 4384 2922 4385
rect 2606 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2922 4384
rect 2606 4319 2922 4320
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 841 3770 907 3773
rect 798 3768 907 3770
rect 798 3712 846 3768
rect 902 3712 907 3768
rect 798 3707 907 3712
rect 798 3664 858 3707
rect 0 3574 858 3664
rect 5349 3634 5415 3637
rect 6100 3634 6900 3664
rect 5349 3632 6900 3634
rect 5349 3576 5354 3632
rect 5410 3576 6900 3632
rect 5349 3574 6900 3576
rect 0 3544 800 3574
rect 5349 3571 5415 3574
rect 6100 3544 6900 3574
rect 2606 3296 2922 3297
rect 2606 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2922 3296
rect 2606 3231 2922 3232
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 841 2410 907 2413
rect 798 2408 907 2410
rect 798 2352 846 2408
rect 902 2352 907 2408
rect 798 2347 907 2352
rect 798 2304 858 2347
rect 0 2214 858 2304
rect 4705 2274 4771 2277
rect 6100 2274 6900 2304
rect 4705 2272 6900 2274
rect 4705 2216 4710 2272
rect 4766 2216 6900 2272
rect 4705 2214 6900 2216
rect 0 2184 800 2214
rect 4705 2211 4771 2214
rect 2606 2208 2922 2209
rect 2606 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2922 2208
rect 6100 2184 6900 2214
rect 2606 2143 2922 2144
rect 0 914 800 944
rect 1669 914 1735 917
rect 0 912 1735 914
rect 0 856 1674 912
rect 1730 856 1735 912
rect 0 854 1735 856
rect 0 824 800 854
rect 1669 851 1735 854
rect 5441 914 5507 917
rect 6100 914 6900 944
rect 5441 912 6900 914
rect 5441 856 5446 912
rect 5502 856 6900 912
rect 5441 854 6900 856
rect 5441 851 5507 854
rect 6100 824 6900 854
<< via3 >>
rect 1952 9276 2016 9280
rect 1952 9220 1956 9276
rect 1956 9220 2012 9276
rect 2012 9220 2016 9276
rect 1952 9216 2016 9220
rect 2032 9276 2096 9280
rect 2032 9220 2036 9276
rect 2036 9220 2092 9276
rect 2092 9220 2096 9276
rect 2032 9216 2096 9220
rect 2112 9276 2176 9280
rect 2112 9220 2116 9276
rect 2116 9220 2172 9276
rect 2172 9220 2176 9276
rect 2112 9216 2176 9220
rect 2192 9276 2256 9280
rect 2192 9220 2196 9276
rect 2196 9220 2252 9276
rect 2252 9220 2256 9276
rect 2192 9216 2256 9220
rect 2612 8732 2676 8736
rect 2612 8676 2616 8732
rect 2616 8676 2672 8732
rect 2672 8676 2676 8732
rect 2612 8672 2676 8676
rect 2692 8732 2756 8736
rect 2692 8676 2696 8732
rect 2696 8676 2752 8732
rect 2752 8676 2756 8732
rect 2692 8672 2756 8676
rect 2772 8732 2836 8736
rect 2772 8676 2776 8732
rect 2776 8676 2832 8732
rect 2832 8676 2836 8732
rect 2772 8672 2836 8676
rect 2852 8732 2916 8736
rect 2852 8676 2856 8732
rect 2856 8676 2912 8732
rect 2912 8676 2916 8732
rect 2852 8672 2916 8676
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 2612 7644 2676 7648
rect 2612 7588 2616 7644
rect 2616 7588 2672 7644
rect 2672 7588 2676 7644
rect 2612 7584 2676 7588
rect 2692 7644 2756 7648
rect 2692 7588 2696 7644
rect 2696 7588 2752 7644
rect 2752 7588 2756 7644
rect 2692 7584 2756 7588
rect 2772 7644 2836 7648
rect 2772 7588 2776 7644
rect 2776 7588 2832 7644
rect 2832 7588 2836 7644
rect 2772 7584 2836 7588
rect 2852 7644 2916 7648
rect 2852 7588 2856 7644
rect 2856 7588 2912 7644
rect 2912 7588 2916 7644
rect 2852 7584 2916 7588
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 2612 6556 2676 6560
rect 2612 6500 2616 6556
rect 2616 6500 2672 6556
rect 2672 6500 2676 6556
rect 2612 6496 2676 6500
rect 2692 6556 2756 6560
rect 2692 6500 2696 6556
rect 2696 6500 2752 6556
rect 2752 6500 2756 6556
rect 2692 6496 2756 6500
rect 2772 6556 2836 6560
rect 2772 6500 2776 6556
rect 2776 6500 2832 6556
rect 2832 6500 2836 6556
rect 2772 6496 2836 6500
rect 2852 6556 2916 6560
rect 2852 6500 2856 6556
rect 2856 6500 2912 6556
rect 2912 6500 2916 6556
rect 2852 6496 2916 6500
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 2612 5468 2676 5472
rect 2612 5412 2616 5468
rect 2616 5412 2672 5468
rect 2672 5412 2676 5468
rect 2612 5408 2676 5412
rect 2692 5468 2756 5472
rect 2692 5412 2696 5468
rect 2696 5412 2752 5468
rect 2752 5412 2756 5468
rect 2692 5408 2756 5412
rect 2772 5468 2836 5472
rect 2772 5412 2776 5468
rect 2776 5412 2832 5468
rect 2832 5412 2836 5468
rect 2772 5408 2836 5412
rect 2852 5468 2916 5472
rect 2852 5412 2856 5468
rect 2856 5412 2912 5468
rect 2912 5412 2916 5468
rect 2852 5408 2916 5412
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 2612 4380 2676 4384
rect 2612 4324 2616 4380
rect 2616 4324 2672 4380
rect 2672 4324 2676 4380
rect 2612 4320 2676 4324
rect 2692 4380 2756 4384
rect 2692 4324 2696 4380
rect 2696 4324 2752 4380
rect 2752 4324 2756 4380
rect 2692 4320 2756 4324
rect 2772 4380 2836 4384
rect 2772 4324 2776 4380
rect 2776 4324 2832 4380
rect 2832 4324 2836 4380
rect 2772 4320 2836 4324
rect 2852 4380 2916 4384
rect 2852 4324 2856 4380
rect 2856 4324 2912 4380
rect 2912 4324 2916 4380
rect 2852 4320 2916 4324
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 2612 3292 2676 3296
rect 2612 3236 2616 3292
rect 2616 3236 2672 3292
rect 2672 3236 2676 3292
rect 2612 3232 2676 3236
rect 2692 3292 2756 3296
rect 2692 3236 2696 3292
rect 2696 3236 2752 3292
rect 2752 3236 2756 3292
rect 2692 3232 2756 3236
rect 2772 3292 2836 3296
rect 2772 3236 2776 3292
rect 2776 3236 2832 3292
rect 2832 3236 2836 3292
rect 2772 3232 2836 3236
rect 2852 3292 2916 3296
rect 2852 3236 2856 3292
rect 2856 3236 2912 3292
rect 2912 3236 2916 3292
rect 2852 3232 2916 3236
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 2612 2204 2676 2208
rect 2612 2148 2616 2204
rect 2616 2148 2672 2204
rect 2672 2148 2676 2204
rect 2612 2144 2676 2148
rect 2692 2204 2756 2208
rect 2692 2148 2696 2204
rect 2696 2148 2752 2204
rect 2752 2148 2756 2204
rect 2692 2144 2756 2148
rect 2772 2204 2836 2208
rect 2772 2148 2776 2204
rect 2776 2148 2832 2204
rect 2832 2148 2836 2204
rect 2772 2144 2836 2148
rect 2852 2204 2916 2208
rect 2852 2148 2856 2204
rect 2856 2148 2912 2204
rect 2912 2148 2916 2204
rect 2852 2144 2916 2148
<< metal4 >>
rect 1944 9280 2264 9296
rect 1944 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2264 9280
rect 1944 8192 2264 9216
rect 1944 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2264 8192
rect 1944 7104 2264 8128
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 2752 2264 3776
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 2128 2264 2688
rect 2604 8736 2924 9296
rect 2604 8672 2612 8736
rect 2676 8672 2692 8736
rect 2756 8672 2772 8736
rect 2836 8672 2852 8736
rect 2916 8672 2924 8736
rect 2604 7648 2924 8672
rect 2604 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2924 7648
rect 2604 6560 2924 7584
rect 2604 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2924 6560
rect 2604 5472 2924 6496
rect 2604 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2924 5472
rect 2604 4384 2924 5408
rect 2604 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2924 4384
rect 2604 3296 2924 4320
rect 2604 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2924 3296
rect 2604 2208 2924 3232
rect 2604 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2924 2208
rect 2604 2128 2924 2144
use sky130_fd_sc_hd__nor2_1  _10_
timestamp 0
transform -1 0 3128 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _11_
timestamp 0
transform 1 0 4232 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _12_
timestamp 0
transform -1 0 2024 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _13_
timestamp 0
transform 1 0 1656 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _14_
timestamp 0
transform -1 0 3864 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _15_
timestamp 0
transform -1 0 2300 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _16_
timestamp 0
transform 1 0 3864 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _17_
timestamp 0
transform -1 0 4416 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _18_
timestamp 0
transform -1 0 2760 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _19_
timestamp 0
transform 1 0 2852 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _20_
timestamp 0
transform -1 0 3312 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _21_
timestamp 0
transform -1 0 4876 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _22_
timestamp 0
transform 1 0 2668 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _23_
timestamp 0
transform 1 0 5152 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _24_
timestamp 0
transform 1 0 2300 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _25_
timestamp 0
transform 1 0 1656 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _26_
timestamp 0
transform 1 0 3312 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _27_
timestamp 0
transform -1 0 2392 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_9
timestamp 0
transform 1 0 1932 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_21
timestamp 0
transform 1 0 3036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 0
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_37
timestamp 0
transform 1 0 4508 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 0
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_15
timestamp 0
transform 1 0 2484 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_23
timestamp 0
transform 1 0 3220 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 0
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_39
timestamp 0
transform 1 0 4692 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_47
timestamp 0
transform 1 0 5428 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 0
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_15
timestamp 0
transform 1 0 2484 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_24
timestamp 0
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_41
timestamp 0
transform 1 0 4876 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_47
timestamp 0
transform 1 0 5428 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_14
timestamp 0
transform 1 0 2392 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_26
timestamp 0
transform 1 0 3496 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_30
timestamp 0
transform 1 0 3864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_36
timestamp 0
transform 1 0 4416 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_15
timestamp 0
transform 1 0 2484 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_26
timestamp 0
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 0
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_41
timestamp 0
transform 1 0 4876 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_47
timestamp 0
transform 1 0 5428 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_6
timestamp 0
transform 1 0 1656 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_14
timestamp 0
transform 1 0 2392 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_18
timestamp 0
transform 1 0 2760 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_30
timestamp 0
transform 1 0 3864 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_42
timestamp 0
transform 1 0 4968 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 0
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_15
timestamp 0
transform 1 0 2484 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_22
timestamp 0
transform 1 0 3128 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_41
timestamp 0
transform 1 0 4876 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_47
timestamp 0
transform 1 0 5428 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_6
timestamp 0
transform 1 0 1656 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_18
timestamp 0
transform 1 0 2760 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_30
timestamp 0
transform 1 0 3864 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_42
timestamp 0
transform 1 0 4968 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_13
timestamp 0
transform 1 0 2300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_25
timestamp 0
transform 1 0 3404 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_41
timestamp 0
transform 1 0 4876 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_3
timestamp 0
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_20
timestamp 0
transform 1 0 2944 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_32
timestamp 0
transform 1 0 4048 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_44
timestamp 0
transform 1 0 5152 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_6
timestamp 0
transform 1 0 1656 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_18
timestamp 0
transform 1 0 2760 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_26
timestamp 0
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_29
timestamp 0
transform 1 0 3772 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_33
timestamp 0
transform 1 0 4140 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_41
timestamp 0
transform 1 0 4876 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 0
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_15
timestamp 0
transform 1 0 2484 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_22
timestamp 0
transform 1 0 3128 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_34
timestamp 0
transform 1 0 4232 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_41
timestamp 0
transform 1 0 4876 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_47
timestamp 0
transform 1 0 5428 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_9
timestamp 0
transform 1 0 1932 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_21
timestamp 0
transform 1 0 3036 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 0
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_29
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_33
timestamp 0
transform 1 0 4140 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_39
timestamp 0
transform 1 0 4692 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 0
transform 1 0 1380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 0
transform 1 0 1656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 0
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 0
transform -1 0 1656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 0
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 0
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 0
transform 1 0 1656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 0
transform 1 0 4784 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 0
transform 1 0 5152 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 0
transform 1 0 5152 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 0
transform 1 0 5152 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 0
transform 1 0 5152 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 0
transform 1 0 5152 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 0
transform -1 0 4968 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output16
timestamp 0
transform 1 0 4968 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_13
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 0
transform -1 0 5796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_14
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 0
transform -1 0 5796 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_15
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 0
transform -1 0 5796 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_16
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 0
transform -1 0 5796 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_17
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 0
transform -1 0 5796 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_18
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 0
transform -1 0 5796 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_19
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 0
transform -1 0 5796 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_20
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 0
transform -1 0 5796 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_21
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 0
transform -1 0 5796 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_22
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 0
transform -1 0 5796 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_23
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 0
transform -1 0 5796 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_24
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 0
transform -1 0 5796 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_25
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 0
transform -1 0 5796 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_26
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_27
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_28
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_29
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_30
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_31
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_32
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
<< labels >>
rlabel metal1 s 3450 8704 3450 8704 4 VGND
rlabel metal1 s 3450 9248 3450 9248 4 VPWR
rlabel metal1 s 3726 7922 3726 7922 4 _00_
rlabel metal2 s 3818 6018 3818 6018 4 _01_
rlabel metal1 s 3588 5066 3588 5066 4 _02_
rlabel metal2 s 3358 6018 3358 6018 4 _03_
rlabel metal1 s 3588 4658 3588 4658 4 _04_
rlabel metal1 s 3726 4114 3726 4114 4 _05_
rlabel metal1 s 2622 5678 2622 5678 4 _06_
rlabel metal1 s 3680 5746 3680 5746 4 _07_
rlabel metal1 s 4232 5678 4232 5678 4 _08_
rlabel metal2 s 3358 3502 3358 3502 4 _09_
rlabel metal3 s 1050 10404 1050 10404 4 in[0]
rlabel metal3 s 0 8984 800 9104 4 in[1]
port 4 nsew
rlabel metal3 s 0 7624 800 7744 4 in[2]
port 5 nsew
rlabel metal3 s 0 6264 800 6384 4 in[3]
port 6 nsew
rlabel metal3 s 0 4904 800 5024 4 in[4]
port 7 nsew
rlabel metal3 s 0 3544 800 3664 4 in[5]
port 8 nsew
rlabel metal3 s 0 2184 800 2304 4 in[6]
port 9 nsew
rlabel metal3 s 1188 884 1188 884 4 in[7]
rlabel metal1 s 1656 6766 1656 6766 4 net1
rlabel metal1 s 4232 3162 4232 3162 4 net10
rlabel metal1 s 5014 7854 5014 7854 4 net11
rlabel metal1 s 3726 6630 3726 6630 4 net12
rlabel metal1 s 5198 5236 5198 5236 4 net13
rlabel metal2 s 5198 4284 5198 4284 4 net14
rlabel metal2 s 4922 3978 4922 3978 4 net15
rlabel metal1 s 4002 7174 4002 7174 4 net16
rlabel metal2 s 1794 5440 1794 5440 4 net2
rlabel metal1 s 3036 7718 3036 7718 4 net3
rlabel metal1 s 1564 6426 1564 6426 4 net4
rlabel metal1 s 4232 4046 4232 4046 4 net5
rlabel metal1 s 3174 4590 3174 4590 4 net6
rlabel metal1 s 3128 3502 3128 3502 4 net7
rlabel metal1 s 2116 2618 2116 2618 4 net8
rlabel metal1 s 3588 3910 3588 3910 4 net9
rlabel metal2 s 5014 9775 5014 9775 4 out[0]
rlabel metal3 s 5382 9061 5382 9061 4 out[1]
rlabel metal3 s 5382 7701 5382 7701 4 out[2]
rlabel metal2 s 5382 6477 5382 6477 4 out[3]
rlabel metal3 s 5382 4981 5382 4981 4 out[4]
rlabel metal2 s 5382 3757 5382 3757 4 out[5]
rlabel metal3 s 4738 2261 4738 2261 4 out[6]
rlabel metal2 s 5474 1615 5474 1615 4 out[7]
flabel metal4 s 2604 2128 2924 9296 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 1944 2128 2264 9296 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal3 s 0 10344 800 10464 0 FreeSans 600 0 0 0 in[0]
port 3 nsew
flabel metal3 s 400 9044 400 9044 0 FreeSans 600 0 0 0 in[1]
flabel metal3 s 400 7684 400 7684 0 FreeSans 600 0 0 0 in[2]
flabel metal3 s 400 6324 400 6324 0 FreeSans 600 0 0 0 in[3]
flabel metal3 s 400 4964 400 4964 0 FreeSans 600 0 0 0 in[4]
flabel metal3 s 400 3604 400 3604 0 FreeSans 600 0 0 0 in[5]
flabel metal3 s 400 2244 400 2244 0 FreeSans 600 0 0 0 in[6]
flabel metal3 s 0 824 800 944 0 FreeSans 600 0 0 0 in[7]
port 10 nsew
flabel metal3 s 6100 10344 6900 10464 0 FreeSans 600 0 0 0 out[0]
port 11 nsew
flabel metal3 s 6100 8984 6900 9104 0 FreeSans 600 0 0 0 out[1]
port 12 nsew
flabel metal3 s 6100 7624 6900 7744 0 FreeSans 600 0 0 0 out[2]
port 13 nsew
flabel metal3 s 6100 6264 6900 6384 0 FreeSans 600 0 0 0 out[3]
port 14 nsew
flabel metal3 s 6100 4904 6900 5024 0 FreeSans 600 0 0 0 out[4]
port 15 nsew
flabel metal3 s 6100 3544 6900 3664 0 FreeSans 600 0 0 0 out[5]
port 16 nsew
flabel metal3 s 6100 2184 6900 2304 0 FreeSans 600 0 0 0 out[6]
port 17 nsew
flabel metal3 s 6100 824 6900 944 0 FreeSans 600 0 0 0 out[7]
port 18 nsew
<< properties >>
string FIXED_BBOX 0 0 6900 11424
<< end >>
