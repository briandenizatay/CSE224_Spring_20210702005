magic
tech sky130A
magscale 1 2
timestamp 1748033116
<< nwell >>
rect 1066 2159 40886 69649
<< obsli1 >>
rect 1104 2159 40848 69649
<< obsm1 >>
rect 1104 2128 40848 69680
<< metal2 >>
rect 2962 71200 3018 72000
rect 8942 71200 8998 72000
rect 14922 71200 14978 72000
rect 20902 71200 20958 72000
rect 26882 71200 26938 72000
rect 32862 71200 32918 72000
rect 38842 71200 38898 72000
rect 2594 0 2650 800
rect 7838 0 7894 800
rect 13082 0 13138 800
rect 18326 0 18382 800
rect 23570 0 23626 800
rect 28814 0 28870 800
rect 34058 0 34114 800
rect 39302 0 39358 800
<< obsm2 >>
rect 1400 71144 2906 71346
rect 3074 71144 8886 71346
rect 9054 71144 14866 71346
rect 15034 71144 20846 71346
rect 21014 71144 26826 71346
rect 26994 71144 32806 71346
rect 32974 71144 38786 71346
rect 38954 71144 40554 71346
rect 1400 856 40554 71144
rect 1400 800 2538 856
rect 2706 800 7782 856
rect 7950 800 13026 856
rect 13194 800 18270 856
rect 18438 800 23514 856
rect 23682 800 28758 856
rect 28926 800 34002 856
rect 34170 800 39246 856
rect 39414 800 40554 856
<< metal3 >>
rect 0 35912 800 36032
rect 41200 35912 42000 36032
<< obsm3 >>
rect 800 36112 41200 69665
rect 880 35832 41120 36112
rect 800 2143 41200 35832
<< metal4 >>
rect 1944 2128 2264 69680
rect 2604 2128 2924 69680
rect 6944 2128 7264 69680
rect 7604 2128 7924 69680
rect 11944 2128 12264 69680
rect 12604 2128 12924 69680
rect 16944 2128 17264 69680
rect 17604 2128 17924 69680
rect 21944 2128 22264 69680
rect 22604 2128 22924 69680
rect 26944 2128 27264 69680
rect 27604 2128 27924 69680
rect 31944 2128 32264 69680
rect 32604 2128 32924 69680
rect 36944 2128 37264 69680
rect 37604 2128 37924 69680
<< obsm4 >>
rect 18091 7787 21864 67693
rect 22344 7787 22524 67693
rect 23004 7787 26864 67693
rect 27344 7787 27524 67693
rect 28004 7787 31864 67693
rect 32344 7787 32524 67693
rect 33004 7787 33981 67693
<< metal5 >>
rect 1056 68676 40896 68996
rect 1056 68016 40896 68336
rect 1056 63676 40896 63996
rect 1056 63016 40896 63336
rect 1056 58676 40896 58996
rect 1056 58016 40896 58336
rect 1056 53676 40896 53996
rect 1056 53016 40896 53336
rect 1056 48676 40896 48996
rect 1056 48016 40896 48336
rect 1056 43676 40896 43996
rect 1056 43016 40896 43336
rect 1056 38676 40896 38996
rect 1056 38016 40896 38336
rect 1056 33676 40896 33996
rect 1056 33016 40896 33336
rect 1056 28676 40896 28996
rect 1056 28016 40896 28336
rect 1056 23676 40896 23996
rect 1056 23016 40896 23336
rect 1056 18676 40896 18996
rect 1056 18016 40896 18336
rect 1056 13676 40896 13996
rect 1056 13016 40896 13336
rect 1056 8676 40896 8996
rect 1056 8016 40896 8336
rect 1056 3676 40896 3996
rect 1056 3016 40896 3336
<< labels >>
rlabel metal4 s 2604 2128 2924 69680 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 7604 2128 7924 69680 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 12604 2128 12924 69680 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 17604 2128 17924 69680 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 22604 2128 22924 69680 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 27604 2128 27924 69680 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 32604 2128 32924 69680 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 37604 2128 37924 69680 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 3676 40896 3996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 8676 40896 8996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 13676 40896 13996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 18676 40896 18996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 23676 40896 23996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 28676 40896 28996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 33676 40896 33996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 38676 40896 38996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 43676 40896 43996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 48676 40896 48996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 53676 40896 53996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 58676 40896 58996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 63676 40896 63996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 68676 40896 68996 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 1944 2128 2264 69680 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 6944 2128 7264 69680 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 11944 2128 12264 69680 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 16944 2128 17264 69680 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 21944 2128 22264 69680 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 26944 2128 27264 69680 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 31944 2128 32264 69680 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 36944 2128 37264 69680 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 3016 40896 3336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 8016 40896 8336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 13016 40896 13336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 18016 40896 18336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 23016 40896 23336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 28016 40896 28336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 33016 40896 33336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 38016 40896 38336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 43016 40896 43336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 48016 40896 48336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 53016 40896 53336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 58016 40896 58336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 63016 40896 63336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 68016 40896 68336 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 39302 0 39358 800 6 an[0]
port 3 nsew signal output
rlabel metal2 s 34058 0 34114 800 6 an[1]
port 4 nsew signal output
rlabel metal2 s 28814 0 28870 800 6 an[2]
port 5 nsew signal output
rlabel metal2 s 23570 0 23626 800 6 an[3]
port 6 nsew signal output
rlabel metal2 s 18326 0 18382 800 6 an[4]
port 7 nsew signal output
rlabel metal2 s 13082 0 13138 800 6 an[5]
port 8 nsew signal output
rlabel metal2 s 7838 0 7894 800 6 an[6]
port 9 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 an[7]
port 10 nsew signal output
rlabel metal3 s 0 35912 800 36032 6 clk
port 11 nsew signal input
rlabel metal3 s 41200 35912 42000 36032 6 rst
port 12 nsew signal input
rlabel metal2 s 38842 71200 38898 72000 6 seg[0]
port 13 nsew signal output
rlabel metal2 s 32862 71200 32918 72000 6 seg[1]
port 14 nsew signal output
rlabel metal2 s 26882 71200 26938 72000 6 seg[2]
port 15 nsew signal output
rlabel metal2 s 20902 71200 20958 72000 6 seg[3]
port 16 nsew signal output
rlabel metal2 s 14922 71200 14978 72000 6 seg[4]
port 17 nsew signal output
rlabel metal2 s 8942 71200 8998 72000 6 seg[5]
port 18 nsew signal output
rlabel metal2 s 2962 71200 3018 72000 6 seg[6]
port 19 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 42000 72000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2566902
string GDS_FILE /openlane/designs/ZeroToFiveCounter/runs/RUN_2025.05.23_20.44.41/results/signoff/ZeroToFiveCounter.magic.gds
string GDS_START 467154
<< end >>

