magic
tech sky130A
magscale 1 2
timestamp 1748033115
<< viali >>
rect 3065 69513 3099 69547
rect 9045 69513 9079 69547
rect 15025 69513 15059 69547
rect 21005 69513 21039 69547
rect 26985 69513 27019 69547
rect 32965 69513 32999 69547
rect 38945 69513 38979 69547
rect 3249 69377 3283 69411
rect 9229 69377 9263 69411
rect 15209 69377 15243 69411
rect 21189 69377 21223 69411
rect 27169 69377 27203 69411
rect 33149 69377 33183 69411
rect 39129 69377 39163 69411
rect 37841 68765 37875 68799
rect 36001 68697 36035 68731
rect 36461 68697 36495 68731
rect 37013 68697 37047 68731
rect 35633 68629 35667 68663
rect 36277 68629 36311 68663
rect 36369 68629 36403 68663
rect 36645 68629 36679 68663
rect 37933 68629 37967 68663
rect 8953 68357 8987 68391
rect 9137 68357 9171 68391
rect 6837 68289 6871 68323
rect 7297 68289 7331 68323
rect 32413 68289 32447 68323
rect 32689 68289 32723 68323
rect 32137 68221 32171 68255
rect 32321 68221 32355 68255
rect 7389 68085 7423 68119
rect 9137 68085 9171 68119
rect 9321 68085 9355 68119
rect 2237 67813 2271 67847
rect 2053 67677 2087 67711
rect 6469 67677 6503 67711
rect 25237 67677 25271 67711
rect 34345 67677 34379 67711
rect 6377 67609 6411 67643
rect 24869 67609 24903 67643
rect 25053 67609 25087 67643
rect 34161 67609 34195 67643
rect 34529 67609 34563 67643
rect 14289 67201 14323 67235
rect 14197 67133 14231 67167
rect 15025 67133 15059 67167
rect 15117 67133 15151 67167
rect 6469 66589 6503 66623
rect 6653 66453 6687 66487
rect 23029 66113 23063 66147
rect 23397 66113 23431 66147
rect 23581 66113 23615 66147
rect 23765 65977 23799 66011
rect 6469 65705 6503 65739
rect 22845 65093 22879 65127
rect 2237 65025 2271 65059
rect 10885 65025 10919 65059
rect 22937 65025 22971 65059
rect 10701 64957 10735 64991
rect 10793 64957 10827 64991
rect 10977 64957 11011 64991
rect 11161 64957 11195 64991
rect 23397 64957 23431 64991
rect 2421 64889 2455 64923
rect 22661 64889 22695 64923
rect 26709 64617 26743 64651
rect 11069 64413 11103 64447
rect 11345 64413 11379 64447
rect 11897 64413 11931 64447
rect 16865 64413 16899 64447
rect 26341 64413 26375 64447
rect 16497 64345 16531 64379
rect 25973 64345 26007 64379
rect 26709 64345 26743 64379
rect 11805 64277 11839 64311
rect 16221 64277 16255 64311
rect 16681 64277 16715 64311
rect 16773 64277 16807 64311
rect 17049 64277 17083 64311
rect 26893 64277 26927 64311
rect 14473 64005 14507 64039
rect 14289 63937 14323 63971
rect 15393 63937 15427 63971
rect 18429 63937 18463 63971
rect 18521 63937 18555 63971
rect 18613 63937 18647 63971
rect 18797 63937 18831 63971
rect 21005 63937 21039 63971
rect 32505 63937 32539 63971
rect 14565 63733 14599 63767
rect 15301 63733 15335 63767
rect 18153 63733 18187 63767
rect 20913 63733 20947 63767
rect 32597 63733 32631 63767
rect 3893 63529 3927 63563
rect 20177 63461 20211 63495
rect 3801 63325 3835 63359
rect 4077 63325 4111 63359
rect 20361 63325 20395 63359
rect 20545 63325 20579 63359
rect 19901 63257 19935 63291
rect 19993 62849 20027 62883
rect 20085 62645 20119 62679
rect 19993 62237 20027 62271
rect 39037 62237 39071 62271
rect 39405 62237 39439 62271
rect 40325 62237 40359 62271
rect 19625 62169 19659 62203
rect 38945 62169 38979 62203
rect 39497 62169 39531 62203
rect 19809 62101 19843 62135
rect 19901 62101 19935 62135
rect 20177 62101 20211 62135
rect 40417 62101 40451 62135
rect 26249 61761 26283 61795
rect 26157 61557 26191 61591
rect 37933 60265 37967 60299
rect 24869 60061 24903 60095
rect 37901 59993 37935 60027
rect 38117 59993 38151 60027
rect 24777 59925 24811 59959
rect 37749 59925 37783 59959
rect 7573 58973 7607 59007
rect 7665 58837 7699 58871
rect 39129 58497 39163 58531
rect 39589 58497 39623 58531
rect 39773 58293 39807 58327
rect 40049 57885 40083 57919
rect 40141 57885 40175 57919
rect 39865 57817 39899 57851
rect 39963 57749 39997 57783
rect 5641 57545 5675 57579
rect 29837 57545 29871 57579
rect 3249 57477 3283 57511
rect 5733 57477 5767 57511
rect 30389 57477 30423 57511
rect 34437 57477 34471 57511
rect 36185 57477 36219 57511
rect 5549 57409 5583 57443
rect 29837 57409 29871 57443
rect 36369 57409 36403 57443
rect 36461 57409 36495 57443
rect 4997 57341 5031 57375
rect 5273 57341 5307 57375
rect 5365 57341 5399 57375
rect 6101 57341 6135 57375
rect 29745 57341 29779 57375
rect 34161 57341 34195 57375
rect 6009 56865 6043 56899
rect 8033 56797 8067 56831
rect 6285 56729 6319 56763
rect 28825 56389 28859 56423
rect 29009 56389 29043 56423
rect 33701 56389 33735 56423
rect 33885 56389 33919 56423
rect 37289 56321 37323 56355
rect 37565 56253 37599 56287
rect 39313 56253 39347 56287
rect 28549 56117 28583 56151
rect 29009 56117 29043 56151
rect 29193 56117 29227 56151
rect 33517 56117 33551 56151
rect 33701 56117 33735 56151
rect 29561 55709 29595 55743
rect 28825 55573 28859 55607
rect 29653 55573 29687 55607
rect 30389 55369 30423 55403
rect 20545 55233 20579 55267
rect 20729 55233 20763 55267
rect 30389 55233 30423 55267
rect 30573 55233 30607 55267
rect 39865 55233 39899 55267
rect 39957 55233 39991 55267
rect 20637 55029 20671 55063
rect 38669 54689 38703 54723
rect 38945 54621 38979 54655
rect 39681 54621 39715 54655
rect 39589 54485 39623 54519
rect 8401 54145 8435 54179
rect 10425 54145 10459 54179
rect 17325 54145 17359 54179
rect 17693 54145 17727 54179
rect 8677 54077 8711 54111
rect 17877 54077 17911 54111
rect 17417 54009 17451 54043
rect 12725 53601 12759 53635
rect 13829 53601 13863 53635
rect 32137 53601 32171 53635
rect 13553 53533 13587 53567
rect 37657 53533 37691 53567
rect 30113 53465 30147 53499
rect 31861 53465 31895 53499
rect 37381 53465 37415 53499
rect 35909 53397 35943 53431
rect 22937 52989 22971 53023
rect 24685 52989 24719 53023
rect 24961 52989 24995 53023
rect 36461 52649 36495 52683
rect 37105 52649 37139 52683
rect 24133 52581 24167 52615
rect 5089 52445 5123 52479
rect 5273 52445 5307 52479
rect 5365 52445 5399 52479
rect 5641 52445 5675 52479
rect 23949 52445 23983 52479
rect 24133 52445 24167 52479
rect 36829 52445 36863 52479
rect 4353 52377 4387 52411
rect 4721 52377 4755 52411
rect 37105 52377 37139 52411
rect 37289 52377 37323 52411
rect 5457 52309 5491 52343
rect 4353 52105 4387 52139
rect 10425 51969 10459 52003
rect 10701 51969 10735 52003
rect 31493 51969 31527 52003
rect 31585 51969 31619 52003
rect 31769 51969 31803 52003
rect 33057 51969 33091 52003
rect 10241 51901 10275 51935
rect 10609 51833 10643 51867
rect 31677 51833 31711 51867
rect 31309 51765 31343 51799
rect 33241 51765 33275 51799
rect 11253 51357 11287 51391
rect 11529 51357 11563 51391
rect 16589 51357 16623 51391
rect 16773 51357 16807 51391
rect 16865 51357 16899 51391
rect 16957 51357 16991 51391
rect 10793 51289 10827 51323
rect 11345 51289 11379 51323
rect 17233 51221 17267 51255
rect 33149 51221 33183 51255
rect 13093 50881 13127 50915
rect 12817 50813 12851 50847
rect 13001 50745 13035 50779
rect 13093 50677 13127 50711
rect 33977 50473 34011 50507
rect 25329 50337 25363 50371
rect 37657 50337 37691 50371
rect 37933 50337 37967 50371
rect 24961 50269 24995 50303
rect 34161 50201 34195 50235
rect 39681 50201 39715 50235
rect 33793 50133 33827 50167
rect 33977 50133 34011 50167
rect 29285 49929 29319 49963
rect 29101 49793 29135 49827
rect 29285 49793 29319 49827
rect 24593 49385 24627 49419
rect 33149 49385 33183 49419
rect 24561 49113 24595 49147
rect 24777 49113 24811 49147
rect 33333 49113 33367 49147
rect 24409 49045 24443 49079
rect 25053 49045 25087 49079
rect 32965 49045 32999 49079
rect 33133 49045 33167 49079
rect 11161 48705 11195 48739
rect 11345 48705 11379 48739
rect 21649 48705 21683 48739
rect 11161 48501 11195 48535
rect 21465 48501 21499 48535
rect 34437 48161 34471 48195
rect 2421 48093 2455 48127
rect 2697 48093 2731 48127
rect 30389 48093 30423 48127
rect 33885 48093 33919 48127
rect 33977 48093 34011 48127
rect 2881 48025 2915 48059
rect 29745 48025 29779 48059
rect 33517 47957 33551 47991
rect 35265 47617 35299 47651
rect 35173 47413 35207 47447
rect 36737 47209 36771 47243
rect 37473 47209 37507 47243
rect 37013 47141 37047 47175
rect 10609 47073 10643 47107
rect 37749 47073 37783 47107
rect 1685 47005 1719 47039
rect 10977 47005 11011 47039
rect 37197 47005 37231 47039
rect 37289 47005 37323 47039
rect 36277 46937 36311 46971
rect 37473 46937 37507 46971
rect 1869 46869 1903 46903
rect 28825 46529 28859 46563
rect 30113 46325 30147 46359
rect 26341 46121 26375 46155
rect 14197 45917 14231 45951
rect 16129 45917 16163 45951
rect 18613 45917 18647 45951
rect 14565 45849 14599 45883
rect 26341 45849 26375 45883
rect 26525 45849 26559 45883
rect 28917 45849 28951 45883
rect 18705 45781 18739 45815
rect 26157 45781 26191 45815
rect 3433 45441 3467 45475
rect 25053 45441 25087 45475
rect 1409 45373 1443 45407
rect 3157 45373 3191 45407
rect 24961 45373 24995 45407
rect 3801 45237 3835 45271
rect 2973 44897 3007 44931
rect 3157 44897 3191 44931
rect 3341 44897 3375 44931
rect 2881 44829 2915 44863
rect 3249 44829 3283 44863
rect 22569 44829 22603 44863
rect 22845 44829 22879 44863
rect 2697 44761 2731 44795
rect 22753 44761 22787 44795
rect 22385 44693 22419 44727
rect 24869 43809 24903 43843
rect 25513 43809 25547 43843
rect 24685 43741 24719 43775
rect 25237 43741 25271 43775
rect 24777 43605 24811 43639
rect 36553 41769 36587 41803
rect 24777 41633 24811 41667
rect 37197 41633 37231 41667
rect 14381 41565 14415 41599
rect 15393 41565 15427 41599
rect 26801 41565 26835 41599
rect 36921 41565 36955 41599
rect 25053 41497 25087 41531
rect 38945 41497 38979 41531
rect 14289 41429 14323 41463
rect 15485 41429 15519 41463
rect 7205 41089 7239 41123
rect 7297 41089 7331 41123
rect 7481 41089 7515 41123
rect 7849 41089 7883 41123
rect 25605 41089 25639 41123
rect 8125 41021 8159 41055
rect 25513 40885 25547 40919
rect 3617 40545 3651 40579
rect 2697 40477 2731 40511
rect 3065 40477 3099 40511
rect 3433 40477 3467 40511
rect 30941 39389 30975 39423
rect 30849 39253 30883 39287
rect 14197 39049 14231 39083
rect 24133 39049 24167 39083
rect 14013 38981 14047 39015
rect 22109 38981 22143 39015
rect 14289 38913 14323 38947
rect 20913 38913 20947 38947
rect 21373 38913 21407 38947
rect 21833 38913 21867 38947
rect 21649 38845 21683 38879
rect 23857 38845 23891 38879
rect 14013 38777 14047 38811
rect 6101 38369 6135 38403
rect 6377 38301 6411 38335
rect 7021 37825 7055 37859
rect 28641 37825 28675 37859
rect 29193 37825 29227 37859
rect 29009 37757 29043 37791
rect 7113 37621 7147 37655
rect 27813 37213 27847 37247
rect 27721 37145 27755 37179
rect 27077 36873 27111 36907
rect 7849 36737 7883 36771
rect 26985 36737 27019 36771
rect 7573 36669 7607 36703
rect 8125 36669 8159 36703
rect 9873 36669 9907 36703
rect 9505 36329 9539 36363
rect 9229 36193 9263 36227
rect 40233 36193 40267 36227
rect 9137 36125 9171 36159
rect 32045 36125 32079 36159
rect 40509 36125 40543 36159
rect 32413 36057 32447 36091
rect 31953 35989 31987 36023
rect 32137 35989 32171 36023
rect 32229 35989 32263 36023
rect 34989 35785 35023 35819
rect 34987 35649 35021 35683
rect 35449 35581 35483 35615
rect 34805 35513 34839 35547
rect 34345 35445 34379 35479
rect 35357 35445 35391 35479
rect 32689 34561 32723 34595
rect 32965 34561 32999 34595
rect 32597 34493 32631 34527
rect 25145 34017 25179 34051
rect 19625 33949 19659 33983
rect 24409 33949 24443 33983
rect 24685 33949 24719 33983
rect 24777 33881 24811 33915
rect 21097 33813 21131 33847
rect 24593 33813 24627 33847
rect 10425 33609 10459 33643
rect 10517 33473 10551 33507
rect 33057 33473 33091 33507
rect 32873 33269 32907 33303
rect 31401 32453 31435 32487
rect 18521 32385 18555 32419
rect 31493 32385 31527 32419
rect 37289 32385 37323 32419
rect 18061 32317 18095 32351
rect 18613 32317 18647 32351
rect 37565 32317 37599 32351
rect 39313 32317 39347 32351
rect 29653 31977 29687 32011
rect 39865 31977 39899 32011
rect 40233 31977 40267 32011
rect 25421 31841 25455 31875
rect 39405 31841 39439 31875
rect 39957 31841 39991 31875
rect 25237 31773 25271 31807
rect 25789 31773 25823 31807
rect 29745 31773 29779 31807
rect 36185 31773 36219 31807
rect 36553 31773 36587 31807
rect 36645 31773 36679 31807
rect 39865 31773 39899 31807
rect 7573 31433 7607 31467
rect 33149 31433 33183 31467
rect 7389 31297 7423 31331
rect 7665 31297 7699 31331
rect 33517 31297 33551 31331
rect 33701 31297 33735 31331
rect 33793 31297 33827 31331
rect 18889 31229 18923 31263
rect 19165 31229 19199 31263
rect 20913 31229 20947 31263
rect 18521 31161 18555 31195
rect 7205 31093 7239 31127
rect 33977 31093 34011 31127
rect 39037 30889 39071 30923
rect 40049 30889 40083 30923
rect 9045 30821 9079 30855
rect 11897 30753 11931 30787
rect 9229 30685 9263 30719
rect 39405 30685 39439 30719
rect 9873 30617 9907 30651
rect 11621 30617 11655 30651
rect 39865 30617 39899 30651
rect 40049 30617 40083 30651
rect 40233 30549 40267 30583
rect 11897 30277 11931 30311
rect 11713 30209 11747 30243
rect 18245 30209 18279 30243
rect 18153 30141 18187 30175
rect 12081 30073 12115 30107
rect 18429 30005 18463 30039
rect 8217 29801 8251 29835
rect 8033 29665 8067 29699
rect 14473 29665 14507 29699
rect 6009 29597 6043 29631
rect 8309 29597 8343 29631
rect 14105 29597 14139 29631
rect 7757 29529 7791 29563
rect 5917 29189 5951 29223
rect 17417 29189 17451 29223
rect 18521 29189 18555 29223
rect 3893 29121 3927 29155
rect 7297 29121 7331 29155
rect 17049 29121 17083 29155
rect 17325 29121 17359 29155
rect 20269 29121 20303 29155
rect 40325 29121 40359 29155
rect 3617 29053 3651 29087
rect 4169 29053 4203 29087
rect 6469 29053 6503 29087
rect 18245 29053 18279 29087
rect 39681 29053 39715 29087
rect 30573 28645 30607 28679
rect 19257 28577 19291 28611
rect 29837 28577 29871 28611
rect 4629 28509 4663 28543
rect 19625 28509 19659 28543
rect 19809 28509 19843 28543
rect 30113 28509 30147 28543
rect 30665 28509 30699 28543
rect 4721 28373 4755 28407
rect 19349 28373 19383 28407
rect 22017 28169 22051 28203
rect 29561 28169 29595 28203
rect 29377 28101 29411 28135
rect 29837 28101 29871 28135
rect 21833 28033 21867 28067
rect 22017 28033 22051 28067
rect 22293 28033 22327 28067
rect 29193 28033 29227 28067
rect 28825 27829 28859 27863
rect 17619 27625 17653 27659
rect 20453 27489 20487 27523
rect 17877 27421 17911 27455
rect 19993 27421 20027 27455
rect 20269 27421 20303 27455
rect 15853 27353 15887 27387
rect 15577 27285 15611 27319
rect 20545 27285 20579 27319
rect 8953 27013 8987 27047
rect 9137 26945 9171 26979
rect 9229 26741 9263 26775
rect 32413 25993 32447 26027
rect 32296 25925 32330 25959
rect 32781 25857 32815 25891
rect 32505 25789 32539 25823
rect 32137 25721 32171 25755
rect 11897 25313 11931 25347
rect 13921 25313 13955 25347
rect 28641 25313 28675 25347
rect 28825 25245 28859 25279
rect 11621 25177 11655 25211
rect 12173 25177 12207 25211
rect 29101 25177 29135 25211
rect 29009 25109 29043 25143
rect 23489 24769 23523 24803
rect 23765 24701 23799 24735
rect 25513 24701 25547 24735
rect 34989 24293 35023 24327
rect 35725 24225 35759 24259
rect 34897 24157 34931 24191
rect 35449 24157 35483 24191
rect 33425 23749 33459 23783
rect 33609 23749 33643 23783
rect 33885 23749 33919 23783
rect 22017 23681 22051 23715
rect 33241 23545 33275 23579
rect 21925 23477 21959 23511
rect 32873 23477 32907 23511
rect 33425 23477 33459 23511
rect 10333 23205 10367 23239
rect 10241 23069 10275 23103
rect 16497 23069 16531 23103
rect 16589 22933 16623 22967
rect 3249 22729 3283 22763
rect 6737 22661 6771 22695
rect 7113 22661 7147 22695
rect 24593 22661 24627 22695
rect 3249 22593 3283 22627
rect 3525 22593 3559 22627
rect 6561 22593 6595 22627
rect 6653 22593 6687 22627
rect 3065 22525 3099 22559
rect 6377 22525 6411 22559
rect 7481 22457 7515 22491
rect 25881 22389 25915 22423
rect 9781 22185 9815 22219
rect 11069 21913 11103 21947
rect 24685 21913 24719 21947
rect 22845 21573 22879 21607
rect 22569 21505 22603 21539
rect 32689 21505 32723 21539
rect 33517 21505 33551 21539
rect 24593 21437 24627 21471
rect 33885 21437 33919 21471
rect 32505 21369 32539 21403
rect 2697 20553 2731 20587
rect 2973 20485 3007 20519
rect 4721 20349 4755 20383
rect 4997 20349 5031 20383
rect 5365 20213 5399 20247
rect 22017 20009 22051 20043
rect 19257 19873 19291 19907
rect 21005 19873 21039 19907
rect 21281 19873 21315 19907
rect 21833 19805 21867 19839
rect 6653 19329 6687 19363
rect 8677 19329 8711 19363
rect 6929 19261 6963 19295
rect 9597 18785 9631 18819
rect 3157 18717 3191 18751
rect 3433 18717 3467 18751
rect 9873 18649 9907 18683
rect 11621 18649 11655 18683
rect 3617 18581 3651 18615
rect 9321 18581 9355 18615
rect 36645 18377 36679 18411
rect 36461 18309 36495 18343
rect 36921 18241 36955 18275
rect 36185 18037 36219 18071
rect 36645 18037 36679 18071
rect 3341 17289 3375 17323
rect 18705 17289 18739 17323
rect 18797 17289 18831 17323
rect 31585 17289 31619 17323
rect 2881 17221 2915 17255
rect 3249 17221 3283 17255
rect 3617 17221 3651 17255
rect 4537 17221 4571 17255
rect 4721 17221 4755 17255
rect 18521 17221 18555 17255
rect 18889 17221 18923 17255
rect 19257 17221 19291 17255
rect 28733 17221 28767 17255
rect 28917 17221 28951 17255
rect 3433 17153 3467 17187
rect 19533 17153 19567 17187
rect 31401 17153 31435 17187
rect 31585 17153 31619 17187
rect 4353 17017 4387 17051
rect 3893 16949 3927 16983
rect 4537 16949 4571 16983
rect 19441 16949 19475 16983
rect 28549 16949 28583 16983
rect 14289 16609 14323 16643
rect 15761 16609 15795 16643
rect 30849 16609 30883 16643
rect 31125 16609 31159 16643
rect 14749 16541 14783 16575
rect 15025 16541 15059 16575
rect 15209 16541 15243 16575
rect 15577 16541 15611 16575
rect 32873 16541 32907 16575
rect 14105 15453 14139 15487
rect 14381 15453 14415 15487
rect 14197 15317 14231 15351
rect 14565 15317 14599 15351
rect 32321 15045 32355 15079
rect 32505 15045 32539 15079
rect 38025 14977 38059 15011
rect 38209 14977 38243 15011
rect 38117 14841 38151 14875
rect 32229 14773 32263 14807
rect 38577 14365 38611 14399
rect 38945 14365 38979 14399
rect 38761 14297 38795 14331
rect 28549 14025 28583 14059
rect 14657 13957 14691 13991
rect 28641 13889 28675 13923
rect 12633 13821 12667 13855
rect 12896 13685 12930 13719
rect 27997 13481 28031 13515
rect 36553 13345 36587 13379
rect 28089 13277 28123 13311
rect 36737 13277 36771 13311
rect 36829 13277 36863 13311
rect 4813 12189 4847 12223
rect 23581 12189 23615 12223
rect 23765 12189 23799 12223
rect 23949 12121 23983 12155
rect 4721 12053 4755 12087
rect 31125 11169 31159 11203
rect 33149 11169 33183 11203
rect 30757 11033 30791 11067
rect 31401 11033 31435 11067
rect 24685 10693 24719 10727
rect 5457 10625 5491 10659
rect 5733 10625 5767 10659
rect 32965 10625 32999 10659
rect 33609 10625 33643 10659
rect 32137 10557 32171 10591
rect 5917 10489 5951 10523
rect 24869 10489 24903 10523
rect 7021 9605 7055 9639
rect 7573 9605 7607 9639
rect 9321 9537 9355 9571
rect 14565 9537 14599 9571
rect 7297 9469 7331 9503
rect 14657 9333 14691 9367
rect 7389 9129 7423 9163
rect 22753 9129 22787 9163
rect 37289 9129 37323 9163
rect 22937 8925 22971 8959
rect 36921 8925 36955 8959
rect 37565 8925 37599 8959
rect 37381 8857 37415 8891
rect 9045 8041 9079 8075
rect 18705 8041 18739 8075
rect 8953 7837 8987 7871
rect 18429 7837 18463 7871
rect 18889 7837 18923 7871
rect 21189 5185 21223 5219
rect 21097 4981 21131 5015
rect 25605 4777 25639 4811
rect 26065 4777 26099 4811
rect 1869 4573 1903 4607
rect 6285 4573 6319 4607
rect 25789 4573 25823 4607
rect 1777 4505 1811 4539
rect 25881 4505 25915 4539
rect 6193 4437 6227 4471
rect 3065 3621 3099 3655
rect 7113 3621 7147 3655
rect 1685 3553 1719 3587
rect 2237 3485 2271 3519
rect 2881 3485 2915 3519
rect 7205 3485 7239 3519
rect 14841 3145 14875 3179
rect 14657 3077 14691 3111
rect 7573 3009 7607 3043
rect 8125 3009 8159 3043
rect 8493 3009 8527 3043
rect 8769 3009 8803 3043
rect 9045 3009 9079 3043
rect 9505 3009 9539 3043
rect 9873 3009 9907 3043
rect 10149 3009 10183 3043
rect 14289 3009 14323 3043
rect 30665 3009 30699 3043
rect 30941 3009 30975 3043
rect 8309 2941 8343 2975
rect 9781 2941 9815 2975
rect 14841 2805 14875 2839
rect 15025 2805 15059 2839
rect 36829 2601 36863 2635
rect 39405 2533 39439 2567
rect 2697 2397 2731 2431
rect 36737 2397 36771 2431
rect 36921 2397 36955 2431
rect 39865 2397 39899 2431
rect 39221 2329 39255 2363
rect 7941 2261 7975 2295
rect 13185 2261 13219 2295
rect 18429 2261 18463 2295
rect 23673 2261 23707 2295
rect 28917 2261 28951 2295
rect 34161 2261 34195 2295
rect 38761 2261 38795 2295
<< metal1 >>
rect 1104 69658 40848 69680
rect 1104 69606 2610 69658
rect 2662 69606 2674 69658
rect 2726 69606 2738 69658
rect 2790 69606 2802 69658
rect 2854 69606 2866 69658
rect 2918 69606 7610 69658
rect 7662 69606 7674 69658
rect 7726 69606 7738 69658
rect 7790 69606 7802 69658
rect 7854 69606 7866 69658
rect 7918 69606 12610 69658
rect 12662 69606 12674 69658
rect 12726 69606 12738 69658
rect 12790 69606 12802 69658
rect 12854 69606 12866 69658
rect 12918 69606 17610 69658
rect 17662 69606 17674 69658
rect 17726 69606 17738 69658
rect 17790 69606 17802 69658
rect 17854 69606 17866 69658
rect 17918 69606 22610 69658
rect 22662 69606 22674 69658
rect 22726 69606 22738 69658
rect 22790 69606 22802 69658
rect 22854 69606 22866 69658
rect 22918 69606 27610 69658
rect 27662 69606 27674 69658
rect 27726 69606 27738 69658
rect 27790 69606 27802 69658
rect 27854 69606 27866 69658
rect 27918 69606 32610 69658
rect 32662 69606 32674 69658
rect 32726 69606 32738 69658
rect 32790 69606 32802 69658
rect 32854 69606 32866 69658
rect 32918 69606 37610 69658
rect 37662 69606 37674 69658
rect 37726 69606 37738 69658
rect 37790 69606 37802 69658
rect 37854 69606 37866 69658
rect 37918 69606 40848 69658
rect 1104 69584 40848 69606
rect 3050 69504 3056 69556
rect 3108 69504 3114 69556
rect 8938 69504 8944 69556
rect 8996 69544 9002 69556
rect 9033 69547 9091 69553
rect 9033 69544 9045 69547
rect 8996 69516 9045 69544
rect 8996 69504 9002 69516
rect 9033 69513 9045 69516
rect 9079 69513 9091 69547
rect 9033 69507 9091 69513
rect 15010 69504 15016 69556
rect 15068 69504 15074 69556
rect 20990 69504 20996 69556
rect 21048 69504 21054 69556
rect 26970 69504 26976 69556
rect 27028 69504 27034 69556
rect 32950 69504 32956 69556
rect 33008 69504 33014 69556
rect 38930 69504 38936 69556
rect 38988 69504 38994 69556
rect 3237 69411 3295 69417
rect 3237 69377 3249 69411
rect 3283 69408 3295 69411
rect 3326 69408 3332 69420
rect 3283 69380 3332 69408
rect 3283 69377 3295 69380
rect 3237 69371 3295 69377
rect 3326 69368 3332 69380
rect 3384 69368 3390 69420
rect 9214 69368 9220 69420
rect 9272 69368 9278 69420
rect 15194 69368 15200 69420
rect 15252 69368 15258 69420
rect 21174 69368 21180 69420
rect 21232 69368 21238 69420
rect 27157 69411 27215 69417
rect 27157 69377 27169 69411
rect 27203 69408 27215 69411
rect 27338 69408 27344 69420
rect 27203 69380 27344 69408
rect 27203 69377 27215 69380
rect 27157 69371 27215 69377
rect 27338 69368 27344 69380
rect 27396 69368 27402 69420
rect 33134 69368 33140 69420
rect 33192 69368 33198 69420
rect 39114 69368 39120 69420
rect 39172 69368 39178 69420
rect 1104 69114 40848 69136
rect 1104 69062 1950 69114
rect 2002 69062 2014 69114
rect 2066 69062 2078 69114
rect 2130 69062 2142 69114
rect 2194 69062 2206 69114
rect 2258 69062 6950 69114
rect 7002 69062 7014 69114
rect 7066 69062 7078 69114
rect 7130 69062 7142 69114
rect 7194 69062 7206 69114
rect 7258 69062 11950 69114
rect 12002 69062 12014 69114
rect 12066 69062 12078 69114
rect 12130 69062 12142 69114
rect 12194 69062 12206 69114
rect 12258 69062 16950 69114
rect 17002 69062 17014 69114
rect 17066 69062 17078 69114
rect 17130 69062 17142 69114
rect 17194 69062 17206 69114
rect 17258 69062 21950 69114
rect 22002 69062 22014 69114
rect 22066 69062 22078 69114
rect 22130 69062 22142 69114
rect 22194 69062 22206 69114
rect 22258 69062 26950 69114
rect 27002 69062 27014 69114
rect 27066 69062 27078 69114
rect 27130 69062 27142 69114
rect 27194 69062 27206 69114
rect 27258 69062 31950 69114
rect 32002 69062 32014 69114
rect 32066 69062 32078 69114
rect 32130 69062 32142 69114
rect 32194 69062 32206 69114
rect 32258 69062 36950 69114
rect 37002 69062 37014 69114
rect 37066 69062 37078 69114
rect 37130 69062 37142 69114
rect 37194 69062 37206 69114
rect 37258 69062 40848 69114
rect 1104 69040 40848 69062
rect 36170 68824 36176 68876
rect 36228 68864 36234 68876
rect 36228 68836 37872 68864
rect 36228 68824 36234 68836
rect 37844 68805 37872 68836
rect 37829 68799 37887 68805
rect 26206 68768 36492 68796
rect 16482 68688 16488 68740
rect 16540 68728 16546 68740
rect 26206 68728 26234 68768
rect 16540 68700 26234 68728
rect 16540 68688 16546 68700
rect 35986 68688 35992 68740
rect 36044 68688 36050 68740
rect 36464 68737 36492 68768
rect 37829 68765 37841 68799
rect 37875 68765 37887 68799
rect 37829 68759 37887 68765
rect 36449 68731 36507 68737
rect 36449 68697 36461 68731
rect 36495 68728 36507 68731
rect 37001 68731 37059 68737
rect 37001 68728 37013 68731
rect 36495 68700 37013 68728
rect 36495 68697 36507 68700
rect 36449 68691 36507 68697
rect 37001 68697 37013 68700
rect 37047 68697 37059 68731
rect 37001 68691 37059 68697
rect 16666 68620 16672 68672
rect 16724 68660 16730 68672
rect 35621 68663 35679 68669
rect 35621 68660 35633 68663
rect 16724 68632 35633 68660
rect 16724 68620 16730 68632
rect 35621 68629 35633 68632
rect 35667 68660 35679 68663
rect 36265 68663 36323 68669
rect 36265 68660 36277 68663
rect 35667 68632 36277 68660
rect 35667 68629 35679 68632
rect 35621 68623 35679 68629
rect 36265 68629 36277 68632
rect 36311 68629 36323 68663
rect 36265 68623 36323 68629
rect 36357 68663 36415 68669
rect 36357 68629 36369 68663
rect 36403 68660 36415 68663
rect 36538 68660 36544 68672
rect 36403 68632 36544 68660
rect 36403 68629 36415 68632
rect 36357 68623 36415 68629
rect 36538 68620 36544 68632
rect 36596 68620 36602 68672
rect 36630 68620 36636 68672
rect 36688 68620 36694 68672
rect 37366 68620 37372 68672
rect 37424 68660 37430 68672
rect 37921 68663 37979 68669
rect 37921 68660 37933 68663
rect 37424 68632 37933 68660
rect 37424 68620 37430 68632
rect 37921 68629 37933 68632
rect 37967 68629 37979 68663
rect 37921 68623 37979 68629
rect 1104 68570 40848 68592
rect 1104 68518 2610 68570
rect 2662 68518 2674 68570
rect 2726 68518 2738 68570
rect 2790 68518 2802 68570
rect 2854 68518 2866 68570
rect 2918 68518 7610 68570
rect 7662 68518 7674 68570
rect 7726 68518 7738 68570
rect 7790 68518 7802 68570
rect 7854 68518 7866 68570
rect 7918 68518 12610 68570
rect 12662 68518 12674 68570
rect 12726 68518 12738 68570
rect 12790 68518 12802 68570
rect 12854 68518 12866 68570
rect 12918 68518 17610 68570
rect 17662 68518 17674 68570
rect 17726 68518 17738 68570
rect 17790 68518 17802 68570
rect 17854 68518 17866 68570
rect 17918 68518 22610 68570
rect 22662 68518 22674 68570
rect 22726 68518 22738 68570
rect 22790 68518 22802 68570
rect 22854 68518 22866 68570
rect 22918 68518 27610 68570
rect 27662 68518 27674 68570
rect 27726 68518 27738 68570
rect 27790 68518 27802 68570
rect 27854 68518 27866 68570
rect 27918 68518 32610 68570
rect 32662 68518 32674 68570
rect 32726 68518 32738 68570
rect 32790 68518 32802 68570
rect 32854 68518 32866 68570
rect 32918 68518 37610 68570
rect 37662 68518 37674 68570
rect 37726 68518 37738 68570
rect 37790 68518 37802 68570
rect 37854 68518 37866 68570
rect 37918 68518 40848 68570
rect 1104 68496 40848 68518
rect 8941 68391 8999 68397
rect 8941 68357 8953 68391
rect 8987 68357 8999 68391
rect 8941 68351 8999 68357
rect 6822 68280 6828 68332
rect 6880 68280 6886 68332
rect 7282 68280 7288 68332
rect 7340 68280 7346 68332
rect 8956 68320 8984 68351
rect 9122 68348 9128 68400
rect 9180 68348 9186 68400
rect 18690 68388 18696 68400
rect 16546 68360 18696 68388
rect 16546 68320 16574 68360
rect 18690 68348 18696 68360
rect 18748 68348 18754 68400
rect 29086 68348 29092 68400
rect 29144 68388 29150 68400
rect 29144 68360 32720 68388
rect 29144 68348 29150 68360
rect 8956 68292 16574 68320
rect 32398 68280 32404 68332
rect 32456 68280 32462 68332
rect 32692 68329 32720 68360
rect 32677 68323 32735 68329
rect 32677 68289 32689 68323
rect 32723 68289 32735 68323
rect 32677 68283 32735 68289
rect 31846 68212 31852 68264
rect 31904 68252 31910 68264
rect 32125 68255 32183 68261
rect 32125 68252 32137 68255
rect 31904 68224 32137 68252
rect 31904 68212 31910 68224
rect 32125 68221 32137 68224
rect 32171 68221 32183 68255
rect 32125 68215 32183 68221
rect 32309 68255 32367 68261
rect 32309 68221 32321 68255
rect 32355 68252 32367 68255
rect 34146 68252 34152 68264
rect 32355 68224 34152 68252
rect 32355 68221 32367 68224
rect 32309 68215 32367 68221
rect 34146 68212 34152 68224
rect 34204 68212 34210 68264
rect 9582 68184 9588 68196
rect 9140 68156 9588 68184
rect 7377 68119 7435 68125
rect 7377 68085 7389 68119
rect 7423 68116 7435 68119
rect 9030 68116 9036 68128
rect 7423 68088 9036 68116
rect 7423 68085 7435 68088
rect 7377 68079 7435 68085
rect 9030 68076 9036 68088
rect 9088 68076 9094 68128
rect 9140 68125 9168 68156
rect 9582 68144 9588 68156
rect 9640 68144 9646 68196
rect 9125 68119 9183 68125
rect 9125 68085 9137 68119
rect 9171 68085 9183 68119
rect 9125 68079 9183 68085
rect 9306 68076 9312 68128
rect 9364 68076 9370 68128
rect 1104 68026 40848 68048
rect 1104 67974 1950 68026
rect 2002 67974 2014 68026
rect 2066 67974 2078 68026
rect 2130 67974 2142 68026
rect 2194 67974 2206 68026
rect 2258 67974 6950 68026
rect 7002 67974 7014 68026
rect 7066 67974 7078 68026
rect 7130 67974 7142 68026
rect 7194 67974 7206 68026
rect 7258 67974 11950 68026
rect 12002 67974 12014 68026
rect 12066 67974 12078 68026
rect 12130 67974 12142 68026
rect 12194 67974 12206 68026
rect 12258 67974 16950 68026
rect 17002 67974 17014 68026
rect 17066 67974 17078 68026
rect 17130 67974 17142 68026
rect 17194 67974 17206 68026
rect 17258 67974 21950 68026
rect 22002 67974 22014 68026
rect 22066 67974 22078 68026
rect 22130 67974 22142 68026
rect 22194 67974 22206 68026
rect 22258 67974 26950 68026
rect 27002 67974 27014 68026
rect 27066 67974 27078 68026
rect 27130 67974 27142 68026
rect 27194 67974 27206 68026
rect 27258 67974 31950 68026
rect 32002 67974 32014 68026
rect 32066 67974 32078 68026
rect 32130 67974 32142 68026
rect 32194 67974 32206 68026
rect 32258 67974 36950 68026
rect 37002 67974 37014 68026
rect 37066 67974 37078 68026
rect 37130 67974 37142 68026
rect 37194 67974 37206 68026
rect 37258 67974 40848 68026
rect 1104 67952 40848 67974
rect 2225 67847 2283 67853
rect 2225 67813 2237 67847
rect 2271 67844 2283 67847
rect 2498 67844 2504 67856
rect 2271 67816 2504 67844
rect 2271 67813 2283 67816
rect 2225 67807 2283 67813
rect 2498 67804 2504 67816
rect 2556 67804 2562 67856
rect 37458 67776 37464 67788
rect 26206 67748 37464 67776
rect 2041 67711 2099 67717
rect 2041 67677 2053 67711
rect 2087 67708 2099 67711
rect 2314 67708 2320 67720
rect 2087 67680 2320 67708
rect 2087 67677 2099 67680
rect 2041 67671 2099 67677
rect 2314 67668 2320 67680
rect 2372 67668 2378 67720
rect 6457 67711 6515 67717
rect 6457 67677 6469 67711
rect 6503 67708 6515 67711
rect 7466 67708 7472 67720
rect 6503 67680 7472 67708
rect 6503 67677 6515 67680
rect 6457 67671 6515 67677
rect 7466 67668 7472 67680
rect 7524 67668 7530 67720
rect 25225 67711 25283 67717
rect 25225 67677 25237 67711
rect 25271 67708 25283 67711
rect 26206 67708 26234 67748
rect 37458 67736 37464 67748
rect 37516 67736 37522 67788
rect 25271 67680 26234 67708
rect 25271 67677 25283 67680
rect 25225 67671 25283 67677
rect 29914 67668 29920 67720
rect 29972 67708 29978 67720
rect 34333 67711 34391 67717
rect 34333 67708 34345 67711
rect 29972 67680 34345 67708
rect 29972 67668 29978 67680
rect 34333 67677 34345 67680
rect 34379 67677 34391 67711
rect 34333 67671 34391 67677
rect 6362 67600 6368 67652
rect 6420 67600 6426 67652
rect 24854 67600 24860 67652
rect 24912 67600 24918 67652
rect 25038 67600 25044 67652
rect 25096 67600 25102 67652
rect 34146 67600 34152 67652
rect 34204 67600 34210 67652
rect 34514 67600 34520 67652
rect 34572 67600 34578 67652
rect 1104 67482 40848 67504
rect 1104 67430 2610 67482
rect 2662 67430 2674 67482
rect 2726 67430 2738 67482
rect 2790 67430 2802 67482
rect 2854 67430 2866 67482
rect 2918 67430 7610 67482
rect 7662 67430 7674 67482
rect 7726 67430 7738 67482
rect 7790 67430 7802 67482
rect 7854 67430 7866 67482
rect 7918 67430 12610 67482
rect 12662 67430 12674 67482
rect 12726 67430 12738 67482
rect 12790 67430 12802 67482
rect 12854 67430 12866 67482
rect 12918 67430 17610 67482
rect 17662 67430 17674 67482
rect 17726 67430 17738 67482
rect 17790 67430 17802 67482
rect 17854 67430 17866 67482
rect 17918 67430 22610 67482
rect 22662 67430 22674 67482
rect 22726 67430 22738 67482
rect 22790 67430 22802 67482
rect 22854 67430 22866 67482
rect 22918 67430 27610 67482
rect 27662 67430 27674 67482
rect 27726 67430 27738 67482
rect 27790 67430 27802 67482
rect 27854 67430 27866 67482
rect 27918 67430 32610 67482
rect 32662 67430 32674 67482
rect 32726 67430 32738 67482
rect 32790 67430 32802 67482
rect 32854 67430 32866 67482
rect 32918 67430 37610 67482
rect 37662 67430 37674 67482
rect 37726 67430 37738 67482
rect 37790 67430 37802 67482
rect 37854 67430 37866 67482
rect 37918 67430 40848 67482
rect 1104 67408 40848 67430
rect 14274 67192 14280 67244
rect 14332 67192 14338 67244
rect 14182 67124 14188 67176
rect 14240 67124 14246 67176
rect 15010 67124 15016 67176
rect 15068 67124 15074 67176
rect 15105 67167 15163 67173
rect 15105 67133 15117 67167
rect 15151 67164 15163 67167
rect 17310 67164 17316 67176
rect 15151 67136 17316 67164
rect 15151 67133 15163 67136
rect 15105 67127 15163 67133
rect 17310 67124 17316 67136
rect 17368 67124 17374 67176
rect 1104 66938 40848 66960
rect 1104 66886 1950 66938
rect 2002 66886 2014 66938
rect 2066 66886 2078 66938
rect 2130 66886 2142 66938
rect 2194 66886 2206 66938
rect 2258 66886 6950 66938
rect 7002 66886 7014 66938
rect 7066 66886 7078 66938
rect 7130 66886 7142 66938
rect 7194 66886 7206 66938
rect 7258 66886 11950 66938
rect 12002 66886 12014 66938
rect 12066 66886 12078 66938
rect 12130 66886 12142 66938
rect 12194 66886 12206 66938
rect 12258 66886 16950 66938
rect 17002 66886 17014 66938
rect 17066 66886 17078 66938
rect 17130 66886 17142 66938
rect 17194 66886 17206 66938
rect 17258 66886 21950 66938
rect 22002 66886 22014 66938
rect 22066 66886 22078 66938
rect 22130 66886 22142 66938
rect 22194 66886 22206 66938
rect 22258 66886 26950 66938
rect 27002 66886 27014 66938
rect 27066 66886 27078 66938
rect 27130 66886 27142 66938
rect 27194 66886 27206 66938
rect 27258 66886 31950 66938
rect 32002 66886 32014 66938
rect 32066 66886 32078 66938
rect 32130 66886 32142 66938
rect 32194 66886 32206 66938
rect 32258 66886 36950 66938
rect 37002 66886 37014 66938
rect 37066 66886 37078 66938
rect 37130 66886 37142 66938
rect 37194 66886 37206 66938
rect 37258 66886 40848 66938
rect 1104 66864 40848 66886
rect 6454 66580 6460 66632
rect 6512 66580 6518 66632
rect 6638 66444 6644 66496
rect 6696 66444 6702 66496
rect 1104 66394 40848 66416
rect 1104 66342 2610 66394
rect 2662 66342 2674 66394
rect 2726 66342 2738 66394
rect 2790 66342 2802 66394
rect 2854 66342 2866 66394
rect 2918 66342 7610 66394
rect 7662 66342 7674 66394
rect 7726 66342 7738 66394
rect 7790 66342 7802 66394
rect 7854 66342 7866 66394
rect 7918 66342 12610 66394
rect 12662 66342 12674 66394
rect 12726 66342 12738 66394
rect 12790 66342 12802 66394
rect 12854 66342 12866 66394
rect 12918 66342 17610 66394
rect 17662 66342 17674 66394
rect 17726 66342 17738 66394
rect 17790 66342 17802 66394
rect 17854 66342 17866 66394
rect 17918 66342 22610 66394
rect 22662 66342 22674 66394
rect 22726 66342 22738 66394
rect 22790 66342 22802 66394
rect 22854 66342 22866 66394
rect 22918 66342 27610 66394
rect 27662 66342 27674 66394
rect 27726 66342 27738 66394
rect 27790 66342 27802 66394
rect 27854 66342 27866 66394
rect 27918 66342 32610 66394
rect 32662 66342 32674 66394
rect 32726 66342 32738 66394
rect 32790 66342 32802 66394
rect 32854 66342 32866 66394
rect 32918 66342 37610 66394
rect 37662 66342 37674 66394
rect 37726 66342 37738 66394
rect 37790 66342 37802 66394
rect 37854 66342 37866 66394
rect 37918 66342 40848 66394
rect 1104 66320 40848 66342
rect 3602 66104 3608 66156
rect 3660 66144 3666 66156
rect 9122 66144 9128 66156
rect 3660 66116 9128 66144
rect 3660 66104 3666 66116
rect 9122 66104 9128 66116
rect 9180 66144 9186 66156
rect 23017 66147 23075 66153
rect 23017 66144 23029 66147
rect 9180 66116 23029 66144
rect 9180 66104 9186 66116
rect 23017 66113 23029 66116
rect 23063 66144 23075 66147
rect 23385 66147 23443 66153
rect 23385 66144 23397 66147
rect 23063 66116 23397 66144
rect 23063 66113 23075 66116
rect 23017 66107 23075 66113
rect 23385 66113 23397 66116
rect 23431 66113 23443 66147
rect 23385 66107 23443 66113
rect 23569 66147 23627 66153
rect 23569 66113 23581 66147
rect 23615 66144 23627 66147
rect 24210 66144 24216 66156
rect 23615 66116 24216 66144
rect 23615 66113 23627 66116
rect 23569 66107 23627 66113
rect 24210 66104 24216 66116
rect 24268 66104 24274 66156
rect 23753 66011 23811 66017
rect 23753 65977 23765 66011
rect 23799 66008 23811 66011
rect 25498 66008 25504 66020
rect 23799 65980 25504 66008
rect 23799 65977 23811 65980
rect 23753 65971 23811 65977
rect 25498 65968 25504 65980
rect 25556 65968 25562 66020
rect 1104 65850 40848 65872
rect 1104 65798 1950 65850
rect 2002 65798 2014 65850
rect 2066 65798 2078 65850
rect 2130 65798 2142 65850
rect 2194 65798 2206 65850
rect 2258 65798 6950 65850
rect 7002 65798 7014 65850
rect 7066 65798 7078 65850
rect 7130 65798 7142 65850
rect 7194 65798 7206 65850
rect 7258 65798 11950 65850
rect 12002 65798 12014 65850
rect 12066 65798 12078 65850
rect 12130 65798 12142 65850
rect 12194 65798 12206 65850
rect 12258 65798 16950 65850
rect 17002 65798 17014 65850
rect 17066 65798 17078 65850
rect 17130 65798 17142 65850
rect 17194 65798 17206 65850
rect 17258 65798 21950 65850
rect 22002 65798 22014 65850
rect 22066 65798 22078 65850
rect 22130 65798 22142 65850
rect 22194 65798 22206 65850
rect 22258 65798 26950 65850
rect 27002 65798 27014 65850
rect 27066 65798 27078 65850
rect 27130 65798 27142 65850
rect 27194 65798 27206 65850
rect 27258 65798 31950 65850
rect 32002 65798 32014 65850
rect 32066 65798 32078 65850
rect 32130 65798 32142 65850
rect 32194 65798 32206 65850
rect 32258 65798 36950 65850
rect 37002 65798 37014 65850
rect 37066 65798 37078 65850
rect 37130 65798 37142 65850
rect 37194 65798 37206 65850
rect 37258 65798 40848 65850
rect 1104 65776 40848 65798
rect 6454 65696 6460 65748
rect 6512 65696 6518 65748
rect 1104 65306 40848 65328
rect 1104 65254 2610 65306
rect 2662 65254 2674 65306
rect 2726 65254 2738 65306
rect 2790 65254 2802 65306
rect 2854 65254 2866 65306
rect 2918 65254 7610 65306
rect 7662 65254 7674 65306
rect 7726 65254 7738 65306
rect 7790 65254 7802 65306
rect 7854 65254 7866 65306
rect 7918 65254 12610 65306
rect 12662 65254 12674 65306
rect 12726 65254 12738 65306
rect 12790 65254 12802 65306
rect 12854 65254 12866 65306
rect 12918 65254 17610 65306
rect 17662 65254 17674 65306
rect 17726 65254 17738 65306
rect 17790 65254 17802 65306
rect 17854 65254 17866 65306
rect 17918 65254 22610 65306
rect 22662 65254 22674 65306
rect 22726 65254 22738 65306
rect 22790 65254 22802 65306
rect 22854 65254 22866 65306
rect 22918 65254 27610 65306
rect 27662 65254 27674 65306
rect 27726 65254 27738 65306
rect 27790 65254 27802 65306
rect 27854 65254 27866 65306
rect 27918 65254 32610 65306
rect 32662 65254 32674 65306
rect 32726 65254 32738 65306
rect 32790 65254 32802 65306
rect 32854 65254 32866 65306
rect 32918 65254 37610 65306
rect 37662 65254 37674 65306
rect 37726 65254 37738 65306
rect 37790 65254 37802 65306
rect 37854 65254 37866 65306
rect 37918 65254 40848 65306
rect 1104 65232 40848 65254
rect 17402 65124 17408 65136
rect 6886 65096 17408 65124
rect 2225 65059 2283 65065
rect 2225 65025 2237 65059
rect 2271 65056 2283 65059
rect 6886 65056 6914 65096
rect 17402 65084 17408 65096
rect 17460 65084 17466 65136
rect 22833 65127 22891 65133
rect 22833 65093 22845 65127
rect 22879 65124 22891 65127
rect 23106 65124 23112 65136
rect 22879 65096 23112 65124
rect 22879 65093 22891 65096
rect 22833 65087 22891 65093
rect 23106 65084 23112 65096
rect 23164 65084 23170 65136
rect 2271 65028 6914 65056
rect 10873 65059 10931 65065
rect 2271 65025 2283 65028
rect 2225 65019 2283 65025
rect 10873 65025 10885 65059
rect 10919 65056 10931 65059
rect 22925 65059 22983 65065
rect 10919 65028 22876 65056
rect 10919 65025 10931 65028
rect 10873 65019 10931 65025
rect 10686 64948 10692 65000
rect 10744 64948 10750 65000
rect 10778 64948 10784 65000
rect 10836 64948 10842 65000
rect 10962 64948 10968 65000
rect 11020 64948 11026 65000
rect 11149 64991 11207 64997
rect 11149 64957 11161 64991
rect 11195 64988 11207 64991
rect 22848 64988 22876 65028
rect 22925 65025 22937 65059
rect 22971 65056 22983 65059
rect 23014 65056 23020 65068
rect 22971 65028 23020 65056
rect 22971 65025 22983 65028
rect 22925 65019 22983 65025
rect 23014 65016 23020 65028
rect 23072 65016 23078 65068
rect 23290 64988 23296 65000
rect 11195 64960 22784 64988
rect 22848 64960 23296 64988
rect 11195 64957 11207 64960
rect 11149 64951 11207 64957
rect 2406 64880 2412 64932
rect 2464 64880 2470 64932
rect 22370 64880 22376 64932
rect 22428 64920 22434 64932
rect 22649 64923 22707 64929
rect 22649 64920 22661 64923
rect 22428 64892 22661 64920
rect 22428 64880 22434 64892
rect 22649 64889 22661 64892
rect 22695 64889 22707 64923
rect 22756 64920 22784 64960
rect 23290 64948 23296 64960
rect 23348 64948 23354 65000
rect 23385 64991 23443 64997
rect 23385 64957 23397 64991
rect 23431 64988 23443 64991
rect 35434 64988 35440 65000
rect 23431 64960 35440 64988
rect 23431 64957 23443 64960
rect 23385 64951 23443 64957
rect 35434 64948 35440 64960
rect 35492 64948 35498 65000
rect 26694 64920 26700 64932
rect 22756 64892 26700 64920
rect 22649 64883 22707 64889
rect 26694 64880 26700 64892
rect 26752 64880 26758 64932
rect 1104 64762 40848 64784
rect 1104 64710 1950 64762
rect 2002 64710 2014 64762
rect 2066 64710 2078 64762
rect 2130 64710 2142 64762
rect 2194 64710 2206 64762
rect 2258 64710 6950 64762
rect 7002 64710 7014 64762
rect 7066 64710 7078 64762
rect 7130 64710 7142 64762
rect 7194 64710 7206 64762
rect 7258 64710 11950 64762
rect 12002 64710 12014 64762
rect 12066 64710 12078 64762
rect 12130 64710 12142 64762
rect 12194 64710 12206 64762
rect 12258 64710 16950 64762
rect 17002 64710 17014 64762
rect 17066 64710 17078 64762
rect 17130 64710 17142 64762
rect 17194 64710 17206 64762
rect 17258 64710 21950 64762
rect 22002 64710 22014 64762
rect 22066 64710 22078 64762
rect 22130 64710 22142 64762
rect 22194 64710 22206 64762
rect 22258 64710 26950 64762
rect 27002 64710 27014 64762
rect 27066 64710 27078 64762
rect 27130 64710 27142 64762
rect 27194 64710 27206 64762
rect 27258 64710 31950 64762
rect 32002 64710 32014 64762
rect 32066 64710 32078 64762
rect 32130 64710 32142 64762
rect 32194 64710 32206 64762
rect 32258 64710 36950 64762
rect 37002 64710 37014 64762
rect 37066 64710 37078 64762
rect 37130 64710 37142 64762
rect 37194 64710 37206 64762
rect 37258 64710 40848 64762
rect 1104 64688 40848 64710
rect 26697 64651 26755 64657
rect 26697 64648 26709 64651
rect 26206 64620 26709 64648
rect 17494 64512 17500 64524
rect 11348 64484 17500 64512
rect 11054 64404 11060 64456
rect 11112 64404 11118 64456
rect 11348 64453 11376 64484
rect 17494 64472 17500 64484
rect 17552 64472 17558 64524
rect 11333 64447 11391 64453
rect 11333 64413 11345 64447
rect 11379 64413 11391 64447
rect 11333 64407 11391 64413
rect 11885 64447 11943 64453
rect 11885 64413 11897 64447
rect 11931 64444 11943 64447
rect 12342 64444 12348 64456
rect 11931 64416 12348 64444
rect 11931 64413 11943 64416
rect 11885 64407 11943 64413
rect 12342 64404 12348 64416
rect 12400 64404 12406 64456
rect 15010 64404 15016 64456
rect 15068 64444 15074 64456
rect 15068 64416 16620 64444
rect 15068 64404 15074 64416
rect 16482 64336 16488 64388
rect 16540 64336 16546 64388
rect 16592 64376 16620 64416
rect 16666 64404 16672 64456
rect 16724 64444 16730 64456
rect 16853 64447 16911 64453
rect 16853 64444 16865 64447
rect 16724 64416 16865 64444
rect 16724 64404 16730 64416
rect 16853 64413 16865 64416
rect 16899 64413 16911 64447
rect 16853 64407 16911 64413
rect 25961 64379 26019 64385
rect 25961 64376 25973 64379
rect 16592 64348 25973 64376
rect 25961 64345 25973 64348
rect 26007 64376 26019 64379
rect 26206 64376 26234 64620
rect 26697 64617 26709 64620
rect 26743 64617 26755 64651
rect 26697 64611 26755 64617
rect 26329 64447 26387 64453
rect 26329 64413 26341 64447
rect 26375 64413 26387 64447
rect 26329 64407 26387 64413
rect 26007 64348 26234 64376
rect 26007 64345 26019 64348
rect 25961 64339 26019 64345
rect 11790 64268 11796 64320
rect 11848 64268 11854 64320
rect 16209 64311 16267 64317
rect 16209 64277 16221 64311
rect 16255 64308 16267 64311
rect 16574 64308 16580 64320
rect 16255 64280 16580 64308
rect 16255 64277 16267 64280
rect 16209 64271 16267 64277
rect 16574 64268 16580 64280
rect 16632 64308 16638 64320
rect 16669 64311 16727 64317
rect 16669 64308 16681 64311
rect 16632 64280 16681 64308
rect 16632 64268 16638 64280
rect 16669 64277 16681 64280
rect 16715 64277 16727 64311
rect 16669 64271 16727 64277
rect 16758 64268 16764 64320
rect 16816 64268 16822 64320
rect 17037 64311 17095 64317
rect 17037 64277 17049 64311
rect 17083 64308 17095 64311
rect 19886 64308 19892 64320
rect 17083 64280 19892 64308
rect 17083 64277 17095 64280
rect 17037 64271 17095 64277
rect 19886 64268 19892 64280
rect 19944 64268 19950 64320
rect 24854 64268 24860 64320
rect 24912 64308 24918 64320
rect 26344 64308 26372 64407
rect 26694 64336 26700 64388
rect 26752 64336 26758 64388
rect 24912 64280 26372 64308
rect 26881 64311 26939 64317
rect 24912 64268 24918 64280
rect 26881 64277 26893 64311
rect 26927 64308 26939 64311
rect 27522 64308 27528 64320
rect 26927 64280 27528 64308
rect 26927 64277 26939 64280
rect 26881 64271 26939 64277
rect 27522 64268 27528 64280
rect 27580 64268 27586 64320
rect 1104 64218 40848 64240
rect 1104 64166 2610 64218
rect 2662 64166 2674 64218
rect 2726 64166 2738 64218
rect 2790 64166 2802 64218
rect 2854 64166 2866 64218
rect 2918 64166 7610 64218
rect 7662 64166 7674 64218
rect 7726 64166 7738 64218
rect 7790 64166 7802 64218
rect 7854 64166 7866 64218
rect 7918 64166 12610 64218
rect 12662 64166 12674 64218
rect 12726 64166 12738 64218
rect 12790 64166 12802 64218
rect 12854 64166 12866 64218
rect 12918 64166 17610 64218
rect 17662 64166 17674 64218
rect 17726 64166 17738 64218
rect 17790 64166 17802 64218
rect 17854 64166 17866 64218
rect 17918 64166 22610 64218
rect 22662 64166 22674 64218
rect 22726 64166 22738 64218
rect 22790 64166 22802 64218
rect 22854 64166 22866 64218
rect 22918 64166 27610 64218
rect 27662 64166 27674 64218
rect 27726 64166 27738 64218
rect 27790 64166 27802 64218
rect 27854 64166 27866 64218
rect 27918 64166 32610 64218
rect 32662 64166 32674 64218
rect 32726 64166 32738 64218
rect 32790 64166 32802 64218
rect 32854 64166 32866 64218
rect 32918 64166 37610 64218
rect 37662 64166 37674 64218
rect 37726 64166 37738 64218
rect 37790 64166 37802 64218
rect 37854 64166 37866 64218
rect 37918 64166 40848 64218
rect 1104 64144 40848 64166
rect 16574 64064 16580 64116
rect 16632 64104 16638 64116
rect 36538 64104 36544 64116
rect 16632 64076 36544 64104
rect 16632 64064 16638 64076
rect 36538 64064 36544 64076
rect 36596 64064 36602 64116
rect 14461 64039 14519 64045
rect 14461 64036 14473 64039
rect 6886 64008 14473 64036
rect 5718 63928 5724 63980
rect 5776 63968 5782 63980
rect 6886 63968 6914 64008
rect 14461 64005 14473 64008
rect 14507 64005 14519 64039
rect 18966 64036 18972 64048
rect 14461 63999 14519 64005
rect 18524 64008 18972 64036
rect 5776 63940 6914 63968
rect 14277 63971 14335 63977
rect 5776 63928 5782 63940
rect 14277 63937 14289 63971
rect 14323 63968 14335 63971
rect 14366 63968 14372 63980
rect 14323 63940 14372 63968
rect 14323 63937 14335 63940
rect 14277 63931 14335 63937
rect 14366 63928 14372 63940
rect 14424 63928 14430 63980
rect 15381 63971 15439 63977
rect 15381 63937 15393 63971
rect 15427 63968 15439 63971
rect 15654 63968 15660 63980
rect 15427 63940 15660 63968
rect 15427 63937 15439 63940
rect 15381 63931 15439 63937
rect 15654 63928 15660 63940
rect 15712 63928 15718 63980
rect 18524 63977 18552 64008
rect 18966 63996 18972 64008
rect 19024 63996 19030 64048
rect 18417 63971 18475 63977
rect 18417 63937 18429 63971
rect 18463 63937 18475 63971
rect 18417 63931 18475 63937
rect 18509 63971 18567 63977
rect 18509 63937 18521 63971
rect 18555 63937 18567 63971
rect 18509 63931 18567 63937
rect 18432 63900 18460 63931
rect 18598 63928 18604 63980
rect 18656 63928 18662 63980
rect 18690 63928 18696 63980
rect 18748 63968 18754 63980
rect 18785 63971 18843 63977
rect 18785 63968 18797 63971
rect 18748 63940 18797 63968
rect 18748 63928 18754 63940
rect 18785 63937 18797 63940
rect 18831 63937 18843 63971
rect 18785 63931 18843 63937
rect 20993 63971 21051 63977
rect 20993 63937 21005 63971
rect 21039 63968 21051 63971
rect 21818 63968 21824 63980
rect 21039 63940 21824 63968
rect 21039 63937 21051 63940
rect 20993 63931 21051 63937
rect 21818 63928 21824 63940
rect 21876 63968 21882 63980
rect 32493 63971 32551 63977
rect 32493 63968 32505 63971
rect 21876 63940 32505 63968
rect 21876 63928 21882 63940
rect 32493 63937 32505 63940
rect 32539 63937 32551 63971
rect 32493 63931 32551 63937
rect 27430 63900 27436 63912
rect 18432 63872 27436 63900
rect 27430 63860 27436 63872
rect 27488 63860 27494 63912
rect 14090 63724 14096 63776
rect 14148 63764 14154 63776
rect 14553 63767 14611 63773
rect 14553 63764 14565 63767
rect 14148 63736 14565 63764
rect 14148 63724 14154 63736
rect 14553 63733 14565 63736
rect 14599 63733 14611 63767
rect 14553 63727 14611 63733
rect 15286 63724 15292 63776
rect 15344 63724 15350 63776
rect 18141 63767 18199 63773
rect 18141 63733 18153 63767
rect 18187 63764 18199 63767
rect 18506 63764 18512 63776
rect 18187 63736 18512 63764
rect 18187 63733 18199 63736
rect 18141 63727 18199 63733
rect 18506 63724 18512 63736
rect 18564 63724 18570 63776
rect 20714 63724 20720 63776
rect 20772 63764 20778 63776
rect 20901 63767 20959 63773
rect 20901 63764 20913 63767
rect 20772 63736 20913 63764
rect 20772 63724 20778 63736
rect 20901 63733 20913 63736
rect 20947 63733 20959 63767
rect 20901 63727 20959 63733
rect 32490 63724 32496 63776
rect 32548 63764 32554 63776
rect 32585 63767 32643 63773
rect 32585 63764 32597 63767
rect 32548 63736 32597 63764
rect 32548 63724 32554 63736
rect 32585 63733 32597 63736
rect 32631 63733 32643 63767
rect 32585 63727 32643 63733
rect 1104 63674 40848 63696
rect 1104 63622 1950 63674
rect 2002 63622 2014 63674
rect 2066 63622 2078 63674
rect 2130 63622 2142 63674
rect 2194 63622 2206 63674
rect 2258 63622 6950 63674
rect 7002 63622 7014 63674
rect 7066 63622 7078 63674
rect 7130 63622 7142 63674
rect 7194 63622 7206 63674
rect 7258 63622 11950 63674
rect 12002 63622 12014 63674
rect 12066 63622 12078 63674
rect 12130 63622 12142 63674
rect 12194 63622 12206 63674
rect 12258 63622 16950 63674
rect 17002 63622 17014 63674
rect 17066 63622 17078 63674
rect 17130 63622 17142 63674
rect 17194 63622 17206 63674
rect 17258 63622 21950 63674
rect 22002 63622 22014 63674
rect 22066 63622 22078 63674
rect 22130 63622 22142 63674
rect 22194 63622 22206 63674
rect 22258 63622 26950 63674
rect 27002 63622 27014 63674
rect 27066 63622 27078 63674
rect 27130 63622 27142 63674
rect 27194 63622 27206 63674
rect 27258 63622 31950 63674
rect 32002 63622 32014 63674
rect 32066 63622 32078 63674
rect 32130 63622 32142 63674
rect 32194 63622 32206 63674
rect 32258 63622 36950 63674
rect 37002 63622 37014 63674
rect 37066 63622 37078 63674
rect 37130 63622 37142 63674
rect 37194 63622 37206 63674
rect 37258 63622 40848 63674
rect 1104 63600 40848 63622
rect 3881 63563 3939 63569
rect 3881 63529 3893 63563
rect 3927 63560 3939 63563
rect 4062 63560 4068 63572
rect 3927 63532 4068 63560
rect 3927 63529 3939 63532
rect 3881 63523 3939 63529
rect 4062 63520 4068 63532
rect 4120 63520 4126 63572
rect 24854 63520 24860 63572
rect 24912 63560 24918 63572
rect 25130 63560 25136 63572
rect 24912 63532 25136 63560
rect 24912 63520 24918 63532
rect 25130 63520 25136 63532
rect 25188 63520 25194 63572
rect 17402 63452 17408 63504
rect 17460 63492 17466 63504
rect 20165 63495 20223 63501
rect 20165 63492 20177 63495
rect 17460 63464 20177 63492
rect 17460 63452 17466 63464
rect 20165 63461 20177 63464
rect 20211 63461 20223 63495
rect 20165 63455 20223 63461
rect 3602 63316 3608 63368
rect 3660 63356 3666 63368
rect 3789 63359 3847 63365
rect 3789 63356 3801 63359
rect 3660 63328 3801 63356
rect 3660 63316 3666 63328
rect 3789 63325 3801 63328
rect 3835 63325 3847 63359
rect 3789 63319 3847 63325
rect 4065 63359 4123 63365
rect 4065 63325 4077 63359
rect 4111 63356 4123 63359
rect 4111 63328 6914 63356
rect 4111 63325 4123 63328
rect 4065 63319 4123 63325
rect 6886 63220 6914 63328
rect 20346 63316 20352 63368
rect 20404 63316 20410 63368
rect 20533 63359 20591 63365
rect 20533 63325 20545 63359
rect 20579 63356 20591 63359
rect 33226 63356 33232 63368
rect 20579 63328 33232 63356
rect 20579 63325 20591 63328
rect 20533 63319 20591 63325
rect 19889 63291 19947 63297
rect 19889 63257 19901 63291
rect 19935 63288 19947 63291
rect 20548 63288 20576 63319
rect 33226 63316 33232 63328
rect 33284 63316 33290 63368
rect 19935 63260 20576 63288
rect 19935 63257 19947 63260
rect 19889 63251 19947 63257
rect 24210 63220 24216 63232
rect 6886 63192 24216 63220
rect 24210 63180 24216 63192
rect 24268 63180 24274 63232
rect 1104 63130 40848 63152
rect 1104 63078 2610 63130
rect 2662 63078 2674 63130
rect 2726 63078 2738 63130
rect 2790 63078 2802 63130
rect 2854 63078 2866 63130
rect 2918 63078 7610 63130
rect 7662 63078 7674 63130
rect 7726 63078 7738 63130
rect 7790 63078 7802 63130
rect 7854 63078 7866 63130
rect 7918 63078 12610 63130
rect 12662 63078 12674 63130
rect 12726 63078 12738 63130
rect 12790 63078 12802 63130
rect 12854 63078 12866 63130
rect 12918 63078 17610 63130
rect 17662 63078 17674 63130
rect 17726 63078 17738 63130
rect 17790 63078 17802 63130
rect 17854 63078 17866 63130
rect 17918 63078 22610 63130
rect 22662 63078 22674 63130
rect 22726 63078 22738 63130
rect 22790 63078 22802 63130
rect 22854 63078 22866 63130
rect 22918 63078 27610 63130
rect 27662 63078 27674 63130
rect 27726 63078 27738 63130
rect 27790 63078 27802 63130
rect 27854 63078 27866 63130
rect 27918 63078 32610 63130
rect 32662 63078 32674 63130
rect 32726 63078 32738 63130
rect 32790 63078 32802 63130
rect 32854 63078 32866 63130
rect 32918 63078 37610 63130
rect 37662 63078 37674 63130
rect 37726 63078 37738 63130
rect 37790 63078 37802 63130
rect 37854 63078 37866 63130
rect 37918 63078 40848 63130
rect 1104 63056 40848 63078
rect 19981 62883 20039 62889
rect 19981 62849 19993 62883
rect 20027 62880 20039 62883
rect 24854 62880 24860 62892
rect 20027 62852 24860 62880
rect 20027 62849 20039 62852
rect 19981 62843 20039 62849
rect 24854 62840 24860 62852
rect 24912 62840 24918 62892
rect 20073 62679 20131 62685
rect 20073 62645 20085 62679
rect 20119 62676 20131 62679
rect 36078 62676 36084 62688
rect 20119 62648 36084 62676
rect 20119 62645 20131 62648
rect 20073 62639 20131 62645
rect 36078 62636 36084 62648
rect 36136 62636 36142 62688
rect 1104 62586 40848 62608
rect 1104 62534 1950 62586
rect 2002 62534 2014 62586
rect 2066 62534 2078 62586
rect 2130 62534 2142 62586
rect 2194 62534 2206 62586
rect 2258 62534 6950 62586
rect 7002 62534 7014 62586
rect 7066 62534 7078 62586
rect 7130 62534 7142 62586
rect 7194 62534 7206 62586
rect 7258 62534 11950 62586
rect 12002 62534 12014 62586
rect 12066 62534 12078 62586
rect 12130 62534 12142 62586
rect 12194 62534 12206 62586
rect 12258 62534 16950 62586
rect 17002 62534 17014 62586
rect 17066 62534 17078 62586
rect 17130 62534 17142 62586
rect 17194 62534 17206 62586
rect 17258 62534 21950 62586
rect 22002 62534 22014 62586
rect 22066 62534 22078 62586
rect 22130 62534 22142 62586
rect 22194 62534 22206 62586
rect 22258 62534 26950 62586
rect 27002 62534 27014 62586
rect 27066 62534 27078 62586
rect 27130 62534 27142 62586
rect 27194 62534 27206 62586
rect 27258 62534 31950 62586
rect 32002 62534 32014 62586
rect 32066 62534 32078 62586
rect 32130 62534 32142 62586
rect 32194 62534 32206 62586
rect 32258 62534 36950 62586
rect 37002 62534 37014 62586
rect 37066 62534 37078 62586
rect 37130 62534 37142 62586
rect 37194 62534 37206 62586
rect 37258 62534 40848 62586
rect 1104 62512 40848 62534
rect 11238 62296 11244 62348
rect 11296 62336 11302 62348
rect 11296 62308 20024 62336
rect 11296 62296 11302 62308
rect 19996 62277 20024 62308
rect 19981 62271 20039 62277
rect 19981 62237 19993 62271
rect 20027 62237 20039 62271
rect 19981 62231 20039 62237
rect 36814 62228 36820 62280
rect 36872 62268 36878 62280
rect 39025 62271 39083 62277
rect 39025 62268 39037 62271
rect 36872 62240 39037 62268
rect 36872 62228 36878 62240
rect 39025 62237 39037 62240
rect 39071 62237 39083 62271
rect 39025 62231 39083 62237
rect 39393 62271 39451 62277
rect 39393 62237 39405 62271
rect 39439 62268 39451 62271
rect 39758 62268 39764 62280
rect 39439 62240 39764 62268
rect 39439 62237 39451 62240
rect 39393 62231 39451 62237
rect 39758 62228 39764 62240
rect 39816 62228 39822 62280
rect 39942 62228 39948 62280
rect 40000 62268 40006 62280
rect 40313 62271 40371 62277
rect 40313 62268 40325 62271
rect 40000 62240 40325 62268
rect 40000 62228 40006 62240
rect 40313 62237 40325 62240
rect 40359 62237 40371 62271
rect 40313 62231 40371 62237
rect 19610 62160 19616 62212
rect 19668 62160 19674 62212
rect 38933 62203 38991 62209
rect 38933 62169 38945 62203
rect 38979 62200 38991 62203
rect 39298 62200 39304 62212
rect 38979 62172 39304 62200
rect 38979 62169 38991 62172
rect 38933 62163 38991 62169
rect 39298 62160 39304 62172
rect 39356 62160 39362 62212
rect 39482 62160 39488 62212
rect 39540 62160 39546 62212
rect 11330 62092 11336 62144
rect 11388 62132 11394 62144
rect 19797 62135 19855 62141
rect 19797 62132 19809 62135
rect 11388 62104 19809 62132
rect 11388 62092 11394 62104
rect 19797 62101 19809 62104
rect 19843 62101 19855 62135
rect 19797 62095 19855 62101
rect 19886 62092 19892 62144
rect 19944 62092 19950 62144
rect 20165 62135 20223 62141
rect 20165 62101 20177 62135
rect 20211 62132 20223 62135
rect 24946 62132 24952 62144
rect 20211 62104 24952 62132
rect 20211 62101 20223 62104
rect 20165 62095 20223 62101
rect 24946 62092 24952 62104
rect 25004 62092 25010 62144
rect 40402 62092 40408 62144
rect 40460 62092 40466 62144
rect 1104 62042 40848 62064
rect 1104 61990 2610 62042
rect 2662 61990 2674 62042
rect 2726 61990 2738 62042
rect 2790 61990 2802 62042
rect 2854 61990 2866 62042
rect 2918 61990 7610 62042
rect 7662 61990 7674 62042
rect 7726 61990 7738 62042
rect 7790 61990 7802 62042
rect 7854 61990 7866 62042
rect 7918 61990 12610 62042
rect 12662 61990 12674 62042
rect 12726 61990 12738 62042
rect 12790 61990 12802 62042
rect 12854 61990 12866 62042
rect 12918 61990 17610 62042
rect 17662 61990 17674 62042
rect 17726 61990 17738 62042
rect 17790 61990 17802 62042
rect 17854 61990 17866 62042
rect 17918 61990 22610 62042
rect 22662 61990 22674 62042
rect 22726 61990 22738 62042
rect 22790 61990 22802 62042
rect 22854 61990 22866 62042
rect 22918 61990 27610 62042
rect 27662 61990 27674 62042
rect 27726 61990 27738 62042
rect 27790 61990 27802 62042
rect 27854 61990 27866 62042
rect 27918 61990 32610 62042
rect 32662 61990 32674 62042
rect 32726 61990 32738 62042
rect 32790 61990 32802 62042
rect 32854 61990 32866 62042
rect 32918 61990 37610 62042
rect 37662 61990 37674 62042
rect 37726 61990 37738 62042
rect 37790 61990 37802 62042
rect 37854 61990 37866 62042
rect 37918 61990 40848 62042
rect 1104 61968 40848 61990
rect 25222 61752 25228 61804
rect 25280 61792 25286 61804
rect 26237 61795 26295 61801
rect 26237 61792 26249 61795
rect 25280 61764 26249 61792
rect 25280 61752 25286 61764
rect 26237 61761 26249 61764
rect 26283 61761 26295 61795
rect 26237 61755 26295 61761
rect 26142 61548 26148 61600
rect 26200 61548 26206 61600
rect 1104 61498 40848 61520
rect 1104 61446 1950 61498
rect 2002 61446 2014 61498
rect 2066 61446 2078 61498
rect 2130 61446 2142 61498
rect 2194 61446 2206 61498
rect 2258 61446 6950 61498
rect 7002 61446 7014 61498
rect 7066 61446 7078 61498
rect 7130 61446 7142 61498
rect 7194 61446 7206 61498
rect 7258 61446 11950 61498
rect 12002 61446 12014 61498
rect 12066 61446 12078 61498
rect 12130 61446 12142 61498
rect 12194 61446 12206 61498
rect 12258 61446 16950 61498
rect 17002 61446 17014 61498
rect 17066 61446 17078 61498
rect 17130 61446 17142 61498
rect 17194 61446 17206 61498
rect 17258 61446 21950 61498
rect 22002 61446 22014 61498
rect 22066 61446 22078 61498
rect 22130 61446 22142 61498
rect 22194 61446 22206 61498
rect 22258 61446 26950 61498
rect 27002 61446 27014 61498
rect 27066 61446 27078 61498
rect 27130 61446 27142 61498
rect 27194 61446 27206 61498
rect 27258 61446 31950 61498
rect 32002 61446 32014 61498
rect 32066 61446 32078 61498
rect 32130 61446 32142 61498
rect 32194 61446 32206 61498
rect 32258 61446 36950 61498
rect 37002 61446 37014 61498
rect 37066 61446 37078 61498
rect 37130 61446 37142 61498
rect 37194 61446 37206 61498
rect 37258 61446 40848 61498
rect 1104 61424 40848 61446
rect 1104 60954 40848 60976
rect 1104 60902 2610 60954
rect 2662 60902 2674 60954
rect 2726 60902 2738 60954
rect 2790 60902 2802 60954
rect 2854 60902 2866 60954
rect 2918 60902 7610 60954
rect 7662 60902 7674 60954
rect 7726 60902 7738 60954
rect 7790 60902 7802 60954
rect 7854 60902 7866 60954
rect 7918 60902 12610 60954
rect 12662 60902 12674 60954
rect 12726 60902 12738 60954
rect 12790 60902 12802 60954
rect 12854 60902 12866 60954
rect 12918 60902 17610 60954
rect 17662 60902 17674 60954
rect 17726 60902 17738 60954
rect 17790 60902 17802 60954
rect 17854 60902 17866 60954
rect 17918 60902 22610 60954
rect 22662 60902 22674 60954
rect 22726 60902 22738 60954
rect 22790 60902 22802 60954
rect 22854 60902 22866 60954
rect 22918 60902 27610 60954
rect 27662 60902 27674 60954
rect 27726 60902 27738 60954
rect 27790 60902 27802 60954
rect 27854 60902 27866 60954
rect 27918 60902 32610 60954
rect 32662 60902 32674 60954
rect 32726 60902 32738 60954
rect 32790 60902 32802 60954
rect 32854 60902 32866 60954
rect 32918 60902 37610 60954
rect 37662 60902 37674 60954
rect 37726 60902 37738 60954
rect 37790 60902 37802 60954
rect 37854 60902 37866 60954
rect 37918 60902 40848 60954
rect 1104 60880 40848 60902
rect 1104 60410 40848 60432
rect 1104 60358 1950 60410
rect 2002 60358 2014 60410
rect 2066 60358 2078 60410
rect 2130 60358 2142 60410
rect 2194 60358 2206 60410
rect 2258 60358 6950 60410
rect 7002 60358 7014 60410
rect 7066 60358 7078 60410
rect 7130 60358 7142 60410
rect 7194 60358 7206 60410
rect 7258 60358 11950 60410
rect 12002 60358 12014 60410
rect 12066 60358 12078 60410
rect 12130 60358 12142 60410
rect 12194 60358 12206 60410
rect 12258 60358 16950 60410
rect 17002 60358 17014 60410
rect 17066 60358 17078 60410
rect 17130 60358 17142 60410
rect 17194 60358 17206 60410
rect 17258 60358 21950 60410
rect 22002 60358 22014 60410
rect 22066 60358 22078 60410
rect 22130 60358 22142 60410
rect 22194 60358 22206 60410
rect 22258 60358 26950 60410
rect 27002 60358 27014 60410
rect 27066 60358 27078 60410
rect 27130 60358 27142 60410
rect 27194 60358 27206 60410
rect 27258 60358 31950 60410
rect 32002 60358 32014 60410
rect 32066 60358 32078 60410
rect 32130 60358 32142 60410
rect 32194 60358 32206 60410
rect 32258 60358 36950 60410
rect 37002 60358 37014 60410
rect 37066 60358 37078 60410
rect 37130 60358 37142 60410
rect 37194 60358 37206 60410
rect 37258 60358 40848 60410
rect 1104 60336 40848 60358
rect 37921 60299 37979 60305
rect 37921 60265 37933 60299
rect 37967 60296 37979 60299
rect 38470 60296 38476 60308
rect 37967 60268 38476 60296
rect 37967 60265 37979 60268
rect 37921 60259 37979 60265
rect 38470 60256 38476 60268
rect 38528 60256 38534 60308
rect 24854 60052 24860 60104
rect 24912 60092 24918 60104
rect 29638 60092 29644 60104
rect 24912 60064 29644 60092
rect 24912 60052 24918 60064
rect 29638 60052 29644 60064
rect 29696 60052 29702 60104
rect 23014 59984 23020 60036
rect 23072 60024 23078 60036
rect 23382 60024 23388 60036
rect 23072 59996 23388 60024
rect 23072 59984 23078 59996
rect 23382 59984 23388 59996
rect 23440 59984 23446 60036
rect 37458 59984 37464 60036
rect 37516 60024 37522 60036
rect 37889 60027 37947 60033
rect 37889 60024 37901 60027
rect 37516 59996 37901 60024
rect 37516 59984 37522 59996
rect 37889 59993 37901 59996
rect 37935 59993 37947 60027
rect 37889 59987 37947 59993
rect 38105 60027 38163 60033
rect 38105 59993 38117 60027
rect 38151 60024 38163 60027
rect 38194 60024 38200 60036
rect 38151 59996 38200 60024
rect 38151 59993 38163 59996
rect 38105 59987 38163 59993
rect 38194 59984 38200 59996
rect 38252 59984 38258 60036
rect 23198 59916 23204 59968
rect 23256 59956 23262 59968
rect 24765 59959 24823 59965
rect 24765 59956 24777 59959
rect 23256 59928 24777 59956
rect 23256 59916 23262 59928
rect 24765 59925 24777 59928
rect 24811 59925 24823 59959
rect 24765 59919 24823 59925
rect 37737 59959 37795 59965
rect 37737 59925 37749 59959
rect 37783 59956 37795 59959
rect 38286 59956 38292 59968
rect 37783 59928 38292 59956
rect 37783 59925 37795 59928
rect 37737 59919 37795 59925
rect 38286 59916 38292 59928
rect 38344 59916 38350 59968
rect 1104 59866 40848 59888
rect 1104 59814 2610 59866
rect 2662 59814 2674 59866
rect 2726 59814 2738 59866
rect 2790 59814 2802 59866
rect 2854 59814 2866 59866
rect 2918 59814 7610 59866
rect 7662 59814 7674 59866
rect 7726 59814 7738 59866
rect 7790 59814 7802 59866
rect 7854 59814 7866 59866
rect 7918 59814 12610 59866
rect 12662 59814 12674 59866
rect 12726 59814 12738 59866
rect 12790 59814 12802 59866
rect 12854 59814 12866 59866
rect 12918 59814 17610 59866
rect 17662 59814 17674 59866
rect 17726 59814 17738 59866
rect 17790 59814 17802 59866
rect 17854 59814 17866 59866
rect 17918 59814 22610 59866
rect 22662 59814 22674 59866
rect 22726 59814 22738 59866
rect 22790 59814 22802 59866
rect 22854 59814 22866 59866
rect 22918 59814 27610 59866
rect 27662 59814 27674 59866
rect 27726 59814 27738 59866
rect 27790 59814 27802 59866
rect 27854 59814 27866 59866
rect 27918 59814 32610 59866
rect 32662 59814 32674 59866
rect 32726 59814 32738 59866
rect 32790 59814 32802 59866
rect 32854 59814 32866 59866
rect 32918 59814 37610 59866
rect 37662 59814 37674 59866
rect 37726 59814 37738 59866
rect 37790 59814 37802 59866
rect 37854 59814 37866 59866
rect 37918 59814 40848 59866
rect 1104 59792 40848 59814
rect 1104 59322 40848 59344
rect 1104 59270 1950 59322
rect 2002 59270 2014 59322
rect 2066 59270 2078 59322
rect 2130 59270 2142 59322
rect 2194 59270 2206 59322
rect 2258 59270 6950 59322
rect 7002 59270 7014 59322
rect 7066 59270 7078 59322
rect 7130 59270 7142 59322
rect 7194 59270 7206 59322
rect 7258 59270 11950 59322
rect 12002 59270 12014 59322
rect 12066 59270 12078 59322
rect 12130 59270 12142 59322
rect 12194 59270 12206 59322
rect 12258 59270 16950 59322
rect 17002 59270 17014 59322
rect 17066 59270 17078 59322
rect 17130 59270 17142 59322
rect 17194 59270 17206 59322
rect 17258 59270 21950 59322
rect 22002 59270 22014 59322
rect 22066 59270 22078 59322
rect 22130 59270 22142 59322
rect 22194 59270 22206 59322
rect 22258 59270 26950 59322
rect 27002 59270 27014 59322
rect 27066 59270 27078 59322
rect 27130 59270 27142 59322
rect 27194 59270 27206 59322
rect 27258 59270 31950 59322
rect 32002 59270 32014 59322
rect 32066 59270 32078 59322
rect 32130 59270 32142 59322
rect 32194 59270 32206 59322
rect 32258 59270 36950 59322
rect 37002 59270 37014 59322
rect 37066 59270 37078 59322
rect 37130 59270 37142 59322
rect 37194 59270 37206 59322
rect 37258 59270 40848 59322
rect 1104 59248 40848 59270
rect 7466 58964 7472 59016
rect 7524 59004 7530 59016
rect 7561 59007 7619 59013
rect 7561 59004 7573 59007
rect 7524 58976 7573 59004
rect 7524 58964 7530 58976
rect 7561 58973 7573 58976
rect 7607 59004 7619 59007
rect 25222 59004 25228 59016
rect 7607 58976 25228 59004
rect 7607 58973 7619 58976
rect 7561 58967 7619 58973
rect 25222 58964 25228 58976
rect 25280 59004 25286 59016
rect 25590 59004 25596 59016
rect 25280 58976 25596 59004
rect 25280 58964 25286 58976
rect 25590 58964 25596 58976
rect 25648 58964 25654 59016
rect 7653 58871 7711 58877
rect 7653 58837 7665 58871
rect 7699 58868 7711 58871
rect 8018 58868 8024 58880
rect 7699 58840 8024 58868
rect 7699 58837 7711 58840
rect 7653 58831 7711 58837
rect 8018 58828 8024 58840
rect 8076 58828 8082 58880
rect 1104 58778 40848 58800
rect 1104 58726 2610 58778
rect 2662 58726 2674 58778
rect 2726 58726 2738 58778
rect 2790 58726 2802 58778
rect 2854 58726 2866 58778
rect 2918 58726 7610 58778
rect 7662 58726 7674 58778
rect 7726 58726 7738 58778
rect 7790 58726 7802 58778
rect 7854 58726 7866 58778
rect 7918 58726 12610 58778
rect 12662 58726 12674 58778
rect 12726 58726 12738 58778
rect 12790 58726 12802 58778
rect 12854 58726 12866 58778
rect 12918 58726 17610 58778
rect 17662 58726 17674 58778
rect 17726 58726 17738 58778
rect 17790 58726 17802 58778
rect 17854 58726 17866 58778
rect 17918 58726 22610 58778
rect 22662 58726 22674 58778
rect 22726 58726 22738 58778
rect 22790 58726 22802 58778
rect 22854 58726 22866 58778
rect 22918 58726 27610 58778
rect 27662 58726 27674 58778
rect 27726 58726 27738 58778
rect 27790 58726 27802 58778
rect 27854 58726 27866 58778
rect 27918 58726 32610 58778
rect 32662 58726 32674 58778
rect 32726 58726 32738 58778
rect 32790 58726 32802 58778
rect 32854 58726 32866 58778
rect 32918 58726 37610 58778
rect 37662 58726 37674 58778
rect 37726 58726 37738 58778
rect 37790 58726 37802 58778
rect 37854 58726 37866 58778
rect 37918 58726 40848 58778
rect 1104 58704 40848 58726
rect 38930 58488 38936 58540
rect 38988 58528 38994 58540
rect 39117 58531 39175 58537
rect 39117 58528 39129 58531
rect 38988 58500 39129 58528
rect 38988 58488 38994 58500
rect 39117 58497 39129 58500
rect 39163 58497 39175 58531
rect 39117 58491 39175 58497
rect 39577 58531 39635 58537
rect 39577 58497 39589 58531
rect 39623 58497 39635 58531
rect 39577 58491 39635 58497
rect 35434 58420 35440 58472
rect 35492 58460 35498 58472
rect 39592 58460 39620 58491
rect 35492 58432 39620 58460
rect 35492 58420 35498 58432
rect 33226 58284 33232 58336
rect 33284 58324 33290 58336
rect 39761 58327 39819 58333
rect 39761 58324 39773 58327
rect 33284 58296 39773 58324
rect 33284 58284 33290 58296
rect 39761 58293 39773 58296
rect 39807 58293 39819 58327
rect 39761 58287 39819 58293
rect 1104 58234 40848 58256
rect 1104 58182 1950 58234
rect 2002 58182 2014 58234
rect 2066 58182 2078 58234
rect 2130 58182 2142 58234
rect 2194 58182 2206 58234
rect 2258 58182 6950 58234
rect 7002 58182 7014 58234
rect 7066 58182 7078 58234
rect 7130 58182 7142 58234
rect 7194 58182 7206 58234
rect 7258 58182 11950 58234
rect 12002 58182 12014 58234
rect 12066 58182 12078 58234
rect 12130 58182 12142 58234
rect 12194 58182 12206 58234
rect 12258 58182 16950 58234
rect 17002 58182 17014 58234
rect 17066 58182 17078 58234
rect 17130 58182 17142 58234
rect 17194 58182 17206 58234
rect 17258 58182 21950 58234
rect 22002 58182 22014 58234
rect 22066 58182 22078 58234
rect 22130 58182 22142 58234
rect 22194 58182 22206 58234
rect 22258 58182 26950 58234
rect 27002 58182 27014 58234
rect 27066 58182 27078 58234
rect 27130 58182 27142 58234
rect 27194 58182 27206 58234
rect 27258 58182 31950 58234
rect 32002 58182 32014 58234
rect 32066 58182 32078 58234
rect 32130 58182 32142 58234
rect 32194 58182 32206 58234
rect 32258 58182 36950 58234
rect 37002 58182 37014 58234
rect 37066 58182 37078 58234
rect 37130 58182 37142 58234
rect 37194 58182 37206 58234
rect 37258 58182 40848 58234
rect 1104 58160 40848 58182
rect 10502 57876 10508 57928
rect 10560 57916 10566 57928
rect 10778 57916 10784 57928
rect 10560 57888 10784 57916
rect 10560 57876 10566 57888
rect 10778 57876 10784 57888
rect 10836 57876 10842 57928
rect 39206 57876 39212 57928
rect 39264 57916 39270 57928
rect 40037 57919 40095 57925
rect 40037 57916 40049 57919
rect 39264 57888 40049 57916
rect 39264 57876 39270 57888
rect 40037 57885 40049 57888
rect 40083 57885 40095 57919
rect 40037 57879 40095 57885
rect 40126 57876 40132 57928
rect 40184 57876 40190 57928
rect 3326 57808 3332 57860
rect 3384 57848 3390 57860
rect 29822 57848 29828 57860
rect 3384 57820 29828 57848
rect 3384 57808 3390 57820
rect 29822 57808 29828 57820
rect 29880 57808 29886 57860
rect 39022 57808 39028 57860
rect 39080 57848 39086 57860
rect 39298 57848 39304 57860
rect 39080 57820 39304 57848
rect 39080 57808 39086 57820
rect 39298 57808 39304 57820
rect 39356 57848 39362 57860
rect 39853 57851 39911 57857
rect 39853 57848 39865 57851
rect 39356 57820 39865 57848
rect 39356 57808 39362 57820
rect 39853 57817 39865 57820
rect 39899 57817 39911 57851
rect 39853 57811 39911 57817
rect 29730 57740 29736 57792
rect 29788 57780 29794 57792
rect 36814 57780 36820 57792
rect 29788 57752 36820 57780
rect 29788 57740 29794 57752
rect 36814 57740 36820 57752
rect 36872 57740 36878 57792
rect 39666 57740 39672 57792
rect 39724 57780 39730 57792
rect 39951 57783 40009 57789
rect 39951 57780 39963 57783
rect 39724 57752 39963 57780
rect 39724 57740 39730 57752
rect 39951 57749 39963 57752
rect 39997 57749 40009 57783
rect 39951 57743 40009 57749
rect 1104 57690 40848 57712
rect 1104 57638 2610 57690
rect 2662 57638 2674 57690
rect 2726 57638 2738 57690
rect 2790 57638 2802 57690
rect 2854 57638 2866 57690
rect 2918 57638 7610 57690
rect 7662 57638 7674 57690
rect 7726 57638 7738 57690
rect 7790 57638 7802 57690
rect 7854 57638 7866 57690
rect 7918 57638 12610 57690
rect 12662 57638 12674 57690
rect 12726 57638 12738 57690
rect 12790 57638 12802 57690
rect 12854 57638 12866 57690
rect 12918 57638 17610 57690
rect 17662 57638 17674 57690
rect 17726 57638 17738 57690
rect 17790 57638 17802 57690
rect 17854 57638 17866 57690
rect 17918 57638 22610 57690
rect 22662 57638 22674 57690
rect 22726 57638 22738 57690
rect 22790 57638 22802 57690
rect 22854 57638 22866 57690
rect 22918 57638 27610 57690
rect 27662 57638 27674 57690
rect 27726 57638 27738 57690
rect 27790 57638 27802 57690
rect 27854 57638 27866 57690
rect 27918 57638 32610 57690
rect 32662 57638 32674 57690
rect 32726 57638 32738 57690
rect 32790 57638 32802 57690
rect 32854 57638 32866 57690
rect 32918 57638 37610 57690
rect 37662 57638 37674 57690
rect 37726 57638 37738 57690
rect 37790 57638 37802 57690
rect 37854 57638 37866 57690
rect 37918 57638 40848 57690
rect 1104 57616 40848 57638
rect 5629 57579 5687 57585
rect 5629 57576 5641 57579
rect 3252 57548 5641 57576
rect 3252 57517 3280 57548
rect 5629 57545 5641 57548
rect 5675 57576 5687 57579
rect 8294 57576 8300 57588
rect 5675 57548 8300 57576
rect 5675 57545 5687 57548
rect 5629 57539 5687 57545
rect 8294 57536 8300 57548
rect 8352 57536 8358 57588
rect 29822 57536 29828 57588
rect 29880 57536 29886 57588
rect 40126 57576 40132 57588
rect 30392 57548 40132 57576
rect 3237 57511 3295 57517
rect 3237 57477 3249 57511
rect 3283 57477 3295 57511
rect 3237 57471 3295 57477
rect 5718 57468 5724 57520
rect 5776 57468 5782 57520
rect 30392 57517 30420 57548
rect 40126 57536 40132 57548
rect 40184 57536 40190 57588
rect 30377 57511 30435 57517
rect 30377 57477 30389 57511
rect 30423 57477 30435 57511
rect 30377 57471 30435 57477
rect 3878 57400 3884 57452
rect 3936 57400 3942 57452
rect 5534 57400 5540 57452
rect 5592 57400 5598 57452
rect 23106 57400 23112 57452
rect 23164 57440 23170 57452
rect 29822 57440 29828 57452
rect 23164 57412 29828 57440
rect 23164 57400 23170 57412
rect 29822 57400 29828 57412
rect 29880 57400 29886 57452
rect 4982 57332 4988 57384
rect 5040 57332 5046 57384
rect 5258 57332 5264 57384
rect 5316 57332 5322 57384
rect 5350 57332 5356 57384
rect 5408 57332 5414 57384
rect 6086 57332 6092 57384
rect 6144 57332 6150 57384
rect 24118 57332 24124 57384
rect 24176 57372 24182 57384
rect 29730 57372 29736 57384
rect 24176 57344 29736 57372
rect 24176 57332 24182 57344
rect 29730 57332 29736 57344
rect 29788 57332 29794 57384
rect 25774 57196 25780 57248
rect 25832 57236 25838 57248
rect 30392 57236 30420 57471
rect 31662 57468 31668 57520
rect 31720 57508 31726 57520
rect 34425 57511 34483 57517
rect 34425 57508 34437 57511
rect 31720 57480 34437 57508
rect 31720 57468 31726 57480
rect 34425 57477 34437 57480
rect 34471 57477 34483 57511
rect 34425 57471 34483 57477
rect 36170 57468 36176 57520
rect 36228 57468 36234 57520
rect 36357 57443 36415 57449
rect 36357 57440 36369 57443
rect 35558 57412 36369 57440
rect 36357 57409 36369 57412
rect 36403 57409 36415 57443
rect 36357 57403 36415 57409
rect 36446 57400 36452 57452
rect 36504 57440 36510 57452
rect 39942 57440 39948 57452
rect 36504 57412 39948 57440
rect 36504 57400 36510 57412
rect 39942 57400 39948 57412
rect 40000 57400 40006 57452
rect 34149 57375 34207 57381
rect 34149 57341 34161 57375
rect 34195 57341 34207 57375
rect 34149 57335 34207 57341
rect 25832 57208 30420 57236
rect 34164 57236 34192 57335
rect 37274 57304 37280 57316
rect 35866 57276 37280 57304
rect 35866 57236 35894 57276
rect 37274 57264 37280 57276
rect 37332 57264 37338 57316
rect 34164 57208 35894 57236
rect 25832 57196 25838 57208
rect 1104 57146 40848 57168
rect 1104 57094 1950 57146
rect 2002 57094 2014 57146
rect 2066 57094 2078 57146
rect 2130 57094 2142 57146
rect 2194 57094 2206 57146
rect 2258 57094 6950 57146
rect 7002 57094 7014 57146
rect 7066 57094 7078 57146
rect 7130 57094 7142 57146
rect 7194 57094 7206 57146
rect 7258 57094 11950 57146
rect 12002 57094 12014 57146
rect 12066 57094 12078 57146
rect 12130 57094 12142 57146
rect 12194 57094 12206 57146
rect 12258 57094 16950 57146
rect 17002 57094 17014 57146
rect 17066 57094 17078 57146
rect 17130 57094 17142 57146
rect 17194 57094 17206 57146
rect 17258 57094 21950 57146
rect 22002 57094 22014 57146
rect 22066 57094 22078 57146
rect 22130 57094 22142 57146
rect 22194 57094 22206 57146
rect 22258 57094 26950 57146
rect 27002 57094 27014 57146
rect 27066 57094 27078 57146
rect 27130 57094 27142 57146
rect 27194 57094 27206 57146
rect 27258 57094 31950 57146
rect 32002 57094 32014 57146
rect 32066 57094 32078 57146
rect 32130 57094 32142 57146
rect 32194 57094 32206 57146
rect 32258 57094 36950 57146
rect 37002 57094 37014 57146
rect 37066 57094 37078 57146
rect 37130 57094 37142 57146
rect 37194 57094 37206 57146
rect 37258 57094 40848 57146
rect 1104 57072 40848 57094
rect 29822 56992 29828 57044
rect 29880 57032 29886 57044
rect 39482 57032 39488 57044
rect 29880 57004 39488 57032
rect 29880 56992 29886 57004
rect 39482 56992 39488 57004
rect 39540 56992 39546 57044
rect 5258 56856 5264 56908
rect 5316 56896 5322 56908
rect 5997 56899 6055 56905
rect 5997 56896 6009 56899
rect 5316 56868 6009 56896
rect 5316 56856 5322 56868
rect 5997 56865 6009 56868
rect 6043 56896 6055 56899
rect 8386 56896 8392 56908
rect 6043 56868 8392 56896
rect 6043 56865 6055 56868
rect 5997 56859 6055 56865
rect 8386 56856 8392 56868
rect 8444 56856 8450 56908
rect 7374 56788 7380 56840
rect 7432 56788 7438 56840
rect 8021 56831 8079 56837
rect 8021 56797 8033 56831
rect 8067 56828 8079 56831
rect 10502 56828 10508 56840
rect 8067 56800 10508 56828
rect 8067 56797 8079 56800
rect 8021 56791 8079 56797
rect 10502 56788 10508 56800
rect 10560 56788 10566 56840
rect 2498 56720 2504 56772
rect 2556 56760 2562 56772
rect 6273 56763 6331 56769
rect 6273 56760 6285 56763
rect 2556 56732 6285 56760
rect 2556 56720 2562 56732
rect 6273 56729 6285 56732
rect 6319 56729 6331 56763
rect 6273 56723 6331 56729
rect 29822 56720 29828 56772
rect 29880 56760 29886 56772
rect 36446 56760 36452 56772
rect 29880 56732 36452 56760
rect 29880 56720 29886 56732
rect 36446 56720 36452 56732
rect 36504 56720 36510 56772
rect 8294 56652 8300 56704
rect 8352 56692 8358 56704
rect 30558 56692 30564 56704
rect 8352 56664 30564 56692
rect 8352 56652 8358 56664
rect 30558 56652 30564 56664
rect 30616 56652 30622 56704
rect 1104 56602 40848 56624
rect 1104 56550 2610 56602
rect 2662 56550 2674 56602
rect 2726 56550 2738 56602
rect 2790 56550 2802 56602
rect 2854 56550 2866 56602
rect 2918 56550 7610 56602
rect 7662 56550 7674 56602
rect 7726 56550 7738 56602
rect 7790 56550 7802 56602
rect 7854 56550 7866 56602
rect 7918 56550 12610 56602
rect 12662 56550 12674 56602
rect 12726 56550 12738 56602
rect 12790 56550 12802 56602
rect 12854 56550 12866 56602
rect 12918 56550 17610 56602
rect 17662 56550 17674 56602
rect 17726 56550 17738 56602
rect 17790 56550 17802 56602
rect 17854 56550 17866 56602
rect 17918 56550 22610 56602
rect 22662 56550 22674 56602
rect 22726 56550 22738 56602
rect 22790 56550 22802 56602
rect 22854 56550 22866 56602
rect 22918 56550 27610 56602
rect 27662 56550 27674 56602
rect 27726 56550 27738 56602
rect 27790 56550 27802 56602
rect 27854 56550 27866 56602
rect 27918 56550 32610 56602
rect 32662 56550 32674 56602
rect 32726 56550 32738 56602
rect 32790 56550 32802 56602
rect 32854 56550 32866 56602
rect 32918 56550 37610 56602
rect 37662 56550 37674 56602
rect 37726 56550 37738 56602
rect 37790 56550 37802 56602
rect 37854 56550 37866 56602
rect 37918 56550 40848 56602
rect 1104 56528 40848 56550
rect 33410 56448 33416 56500
rect 33468 56488 33474 56500
rect 34146 56488 34152 56500
rect 33468 56460 34152 56488
rect 33468 56448 33474 56460
rect 34146 56448 34152 56460
rect 34204 56448 34210 56500
rect 28534 56380 28540 56432
rect 28592 56420 28598 56432
rect 28813 56423 28871 56429
rect 28813 56420 28825 56423
rect 28592 56392 28825 56420
rect 28592 56380 28598 56392
rect 28813 56389 28825 56392
rect 28859 56389 28871 56423
rect 28813 56383 28871 56389
rect 28994 56380 29000 56432
rect 29052 56380 29058 56432
rect 33686 56380 33692 56432
rect 33744 56380 33750 56432
rect 33870 56380 33876 56432
rect 33928 56380 33934 56432
rect 37458 56420 37464 56432
rect 37292 56392 37464 56420
rect 37292 56364 37320 56392
rect 37458 56380 37464 56392
rect 37516 56380 37522 56432
rect 38838 56420 38844 56432
rect 38778 56392 38844 56420
rect 38838 56380 38844 56392
rect 38896 56380 38902 56432
rect 37274 56312 37280 56364
rect 37332 56312 37338 56364
rect 37553 56287 37611 56293
rect 37553 56253 37565 56287
rect 37599 56284 37611 56287
rect 38010 56284 38016 56296
rect 37599 56256 38016 56284
rect 37599 56253 37611 56256
rect 37553 56247 37611 56253
rect 38010 56244 38016 56256
rect 38068 56244 38074 56296
rect 38102 56244 38108 56296
rect 38160 56284 38166 56296
rect 39301 56287 39359 56293
rect 39301 56284 39313 56287
rect 38160 56256 39313 56284
rect 38160 56244 38166 56256
rect 39301 56253 39313 56256
rect 39347 56253 39359 56287
rect 39301 56247 39359 56253
rect 28534 56108 28540 56160
rect 28592 56108 28598 56160
rect 28626 56108 28632 56160
rect 28684 56148 28690 56160
rect 28997 56151 29055 56157
rect 28997 56148 29009 56151
rect 28684 56120 29009 56148
rect 28684 56108 28690 56120
rect 28997 56117 29009 56120
rect 29043 56117 29055 56151
rect 28997 56111 29055 56117
rect 29178 56108 29184 56160
rect 29236 56108 29242 56160
rect 33502 56108 33508 56160
rect 33560 56108 33566 56160
rect 33594 56108 33600 56160
rect 33652 56148 33658 56160
rect 33689 56151 33747 56157
rect 33689 56148 33701 56151
rect 33652 56120 33701 56148
rect 33652 56108 33658 56120
rect 33689 56117 33701 56120
rect 33735 56117 33747 56151
rect 33689 56111 33747 56117
rect 1104 56058 40848 56080
rect 1104 56006 1950 56058
rect 2002 56006 2014 56058
rect 2066 56006 2078 56058
rect 2130 56006 2142 56058
rect 2194 56006 2206 56058
rect 2258 56006 6950 56058
rect 7002 56006 7014 56058
rect 7066 56006 7078 56058
rect 7130 56006 7142 56058
rect 7194 56006 7206 56058
rect 7258 56006 11950 56058
rect 12002 56006 12014 56058
rect 12066 56006 12078 56058
rect 12130 56006 12142 56058
rect 12194 56006 12206 56058
rect 12258 56006 16950 56058
rect 17002 56006 17014 56058
rect 17066 56006 17078 56058
rect 17130 56006 17142 56058
rect 17194 56006 17206 56058
rect 17258 56006 21950 56058
rect 22002 56006 22014 56058
rect 22066 56006 22078 56058
rect 22130 56006 22142 56058
rect 22194 56006 22206 56058
rect 22258 56006 26950 56058
rect 27002 56006 27014 56058
rect 27066 56006 27078 56058
rect 27130 56006 27142 56058
rect 27194 56006 27206 56058
rect 27258 56006 31950 56058
rect 32002 56006 32014 56058
rect 32066 56006 32078 56058
rect 32130 56006 32142 56058
rect 32194 56006 32206 56058
rect 32258 56006 36950 56058
rect 37002 56006 37014 56058
rect 37066 56006 37078 56058
rect 37130 56006 37142 56058
rect 37194 56006 37206 56058
rect 37258 56006 40848 56058
rect 1104 55984 40848 56006
rect 12342 55836 12348 55888
rect 12400 55876 12406 55888
rect 38102 55876 38108 55888
rect 12400 55848 38108 55876
rect 12400 55836 12406 55848
rect 38102 55836 38108 55848
rect 38160 55836 38166 55888
rect 21450 55768 21456 55820
rect 21508 55808 21514 55820
rect 21818 55808 21824 55820
rect 21508 55780 21824 55808
rect 21508 55768 21514 55780
rect 21818 55768 21824 55780
rect 21876 55808 21882 55820
rect 21876 55780 26234 55808
rect 21876 55768 21882 55780
rect 26206 55740 26234 55780
rect 29549 55743 29607 55749
rect 29549 55740 29561 55743
rect 26206 55712 29561 55740
rect 29549 55709 29561 55712
rect 29595 55709 29607 55743
rect 29549 55703 29607 55709
rect 20530 55632 20536 55684
rect 20588 55672 20594 55684
rect 33410 55672 33416 55684
rect 20588 55644 33416 55672
rect 20588 55632 20594 55644
rect 33410 55632 33416 55644
rect 33468 55632 33474 55684
rect 28626 55564 28632 55616
rect 28684 55604 28690 55616
rect 28813 55607 28871 55613
rect 28813 55604 28825 55607
rect 28684 55576 28825 55604
rect 28684 55564 28690 55576
rect 28813 55573 28825 55576
rect 28859 55573 28871 55607
rect 28813 55567 28871 55573
rect 29638 55564 29644 55616
rect 29696 55564 29702 55616
rect 1104 55514 40848 55536
rect 1104 55462 2610 55514
rect 2662 55462 2674 55514
rect 2726 55462 2738 55514
rect 2790 55462 2802 55514
rect 2854 55462 2866 55514
rect 2918 55462 7610 55514
rect 7662 55462 7674 55514
rect 7726 55462 7738 55514
rect 7790 55462 7802 55514
rect 7854 55462 7866 55514
rect 7918 55462 12610 55514
rect 12662 55462 12674 55514
rect 12726 55462 12738 55514
rect 12790 55462 12802 55514
rect 12854 55462 12866 55514
rect 12918 55462 17610 55514
rect 17662 55462 17674 55514
rect 17726 55462 17738 55514
rect 17790 55462 17802 55514
rect 17854 55462 17866 55514
rect 17918 55462 22610 55514
rect 22662 55462 22674 55514
rect 22726 55462 22738 55514
rect 22790 55462 22802 55514
rect 22854 55462 22866 55514
rect 22918 55462 27610 55514
rect 27662 55462 27674 55514
rect 27726 55462 27738 55514
rect 27790 55462 27802 55514
rect 27854 55462 27866 55514
rect 27918 55462 32610 55514
rect 32662 55462 32674 55514
rect 32726 55462 32738 55514
rect 32790 55462 32802 55514
rect 32854 55462 32866 55514
rect 32918 55462 37610 55514
rect 37662 55462 37674 55514
rect 37726 55462 37738 55514
rect 37790 55462 37802 55514
rect 37854 55462 37866 55514
rect 37918 55462 40848 55514
rect 1104 55440 40848 55462
rect 20732 55372 27384 55400
rect 16850 55292 16856 55344
rect 16908 55332 16914 55344
rect 20732 55332 20760 55372
rect 16908 55304 20760 55332
rect 16908 55292 16914 55304
rect 20530 55224 20536 55276
rect 20588 55224 20594 55276
rect 20732 55273 20760 55304
rect 22278 55292 22284 55344
rect 22336 55332 22342 55344
rect 27356 55332 27384 55372
rect 27430 55360 27436 55412
rect 27488 55400 27494 55412
rect 30377 55403 30435 55409
rect 30377 55400 30389 55403
rect 27488 55372 30389 55400
rect 27488 55360 27494 55372
rect 30377 55369 30389 55372
rect 30423 55369 30435 55403
rect 30377 55363 30435 55369
rect 29914 55332 29920 55344
rect 22336 55304 26234 55332
rect 27356 55304 29920 55332
rect 22336 55292 22342 55304
rect 20717 55267 20775 55273
rect 20717 55233 20729 55267
rect 20763 55233 20775 55267
rect 26206 55264 26234 55304
rect 29914 55292 29920 55304
rect 29972 55292 29978 55344
rect 30377 55267 30435 55273
rect 30377 55264 30389 55267
rect 26206 55236 30389 55264
rect 20717 55227 20775 55233
rect 30377 55233 30389 55236
rect 30423 55233 30435 55267
rect 30377 55227 30435 55233
rect 30558 55224 30564 55276
rect 30616 55224 30622 55276
rect 39850 55224 39856 55276
rect 39908 55224 39914 55276
rect 39942 55224 39948 55276
rect 40000 55224 40006 55276
rect 20625 55063 20683 55069
rect 20625 55029 20637 55063
rect 20671 55060 20683 55063
rect 23014 55060 23020 55072
rect 20671 55032 23020 55060
rect 20671 55029 20683 55032
rect 20625 55023 20683 55029
rect 23014 55020 23020 55032
rect 23072 55020 23078 55072
rect 1104 54970 40848 54992
rect 1104 54918 1950 54970
rect 2002 54918 2014 54970
rect 2066 54918 2078 54970
rect 2130 54918 2142 54970
rect 2194 54918 2206 54970
rect 2258 54918 6950 54970
rect 7002 54918 7014 54970
rect 7066 54918 7078 54970
rect 7130 54918 7142 54970
rect 7194 54918 7206 54970
rect 7258 54918 11950 54970
rect 12002 54918 12014 54970
rect 12066 54918 12078 54970
rect 12130 54918 12142 54970
rect 12194 54918 12206 54970
rect 12258 54918 16950 54970
rect 17002 54918 17014 54970
rect 17066 54918 17078 54970
rect 17130 54918 17142 54970
rect 17194 54918 17206 54970
rect 17258 54918 21950 54970
rect 22002 54918 22014 54970
rect 22066 54918 22078 54970
rect 22130 54918 22142 54970
rect 22194 54918 22206 54970
rect 22258 54918 26950 54970
rect 27002 54918 27014 54970
rect 27066 54918 27078 54970
rect 27130 54918 27142 54970
rect 27194 54918 27206 54970
rect 27258 54918 31950 54970
rect 32002 54918 32014 54970
rect 32066 54918 32078 54970
rect 32130 54918 32142 54970
rect 32194 54918 32206 54970
rect 32258 54918 36950 54970
rect 37002 54918 37014 54970
rect 37066 54918 37078 54970
rect 37130 54918 37142 54970
rect 37194 54918 37206 54970
rect 37258 54918 40848 54970
rect 1104 54896 40848 54918
rect 23382 54680 23388 54732
rect 23440 54720 23446 54732
rect 38657 54723 38715 54729
rect 38657 54720 38669 54723
rect 23440 54692 38669 54720
rect 23440 54680 23446 54692
rect 38657 54689 38669 54692
rect 38703 54720 38715 54723
rect 39022 54720 39028 54732
rect 38703 54692 39028 54720
rect 38703 54689 38715 54692
rect 38657 54683 38715 54689
rect 39022 54680 39028 54692
rect 39080 54680 39086 54732
rect 38933 54655 38991 54661
rect 38933 54621 38945 54655
rect 38979 54652 38991 54655
rect 39206 54652 39212 54664
rect 38979 54624 39212 54652
rect 38979 54621 38991 54624
rect 38933 54615 38991 54621
rect 22370 54476 22376 54528
rect 22428 54516 22434 54528
rect 34974 54516 34980 54528
rect 22428 54488 34980 54516
rect 22428 54476 22434 54488
rect 34974 54476 34980 54488
rect 35032 54516 35038 54528
rect 38948 54516 38976 54615
rect 39206 54612 39212 54624
rect 39264 54612 39270 54664
rect 39666 54612 39672 54664
rect 39724 54612 39730 54664
rect 35032 54488 38976 54516
rect 35032 54476 35038 54488
rect 39574 54476 39580 54528
rect 39632 54476 39638 54528
rect 1104 54426 40848 54448
rect 1104 54374 2610 54426
rect 2662 54374 2674 54426
rect 2726 54374 2738 54426
rect 2790 54374 2802 54426
rect 2854 54374 2866 54426
rect 2918 54374 7610 54426
rect 7662 54374 7674 54426
rect 7726 54374 7738 54426
rect 7790 54374 7802 54426
rect 7854 54374 7866 54426
rect 7918 54374 12610 54426
rect 12662 54374 12674 54426
rect 12726 54374 12738 54426
rect 12790 54374 12802 54426
rect 12854 54374 12866 54426
rect 12918 54374 17610 54426
rect 17662 54374 17674 54426
rect 17726 54374 17738 54426
rect 17790 54374 17802 54426
rect 17854 54374 17866 54426
rect 17918 54374 22610 54426
rect 22662 54374 22674 54426
rect 22726 54374 22738 54426
rect 22790 54374 22802 54426
rect 22854 54374 22866 54426
rect 22918 54374 27610 54426
rect 27662 54374 27674 54426
rect 27726 54374 27738 54426
rect 27790 54374 27802 54426
rect 27854 54374 27866 54426
rect 27918 54374 32610 54426
rect 32662 54374 32674 54426
rect 32726 54374 32738 54426
rect 32790 54374 32802 54426
rect 32854 54374 32866 54426
rect 32918 54374 37610 54426
rect 37662 54374 37674 54426
rect 37726 54374 37738 54426
rect 37790 54374 37802 54426
rect 37854 54374 37866 54426
rect 37918 54374 40848 54426
rect 1104 54352 40848 54374
rect 23106 54244 23112 54256
rect 17328 54216 23112 54244
rect 8386 54136 8392 54188
rect 8444 54136 8450 54188
rect 9766 54136 9772 54188
rect 9824 54136 9830 54188
rect 10413 54179 10471 54185
rect 10413 54145 10425 54179
rect 10459 54176 10471 54179
rect 14734 54176 14740 54188
rect 10459 54148 14740 54176
rect 10459 54145 10471 54148
rect 10413 54139 10471 54145
rect 14734 54136 14740 54148
rect 14792 54176 14798 54188
rect 17328 54185 17356 54216
rect 23106 54204 23112 54216
rect 23164 54204 23170 54256
rect 17313 54179 17371 54185
rect 17313 54176 17325 54179
rect 14792 54148 17325 54176
rect 14792 54136 14798 54148
rect 17313 54145 17325 54148
rect 17359 54145 17371 54179
rect 17313 54139 17371 54145
rect 17681 54179 17739 54185
rect 17681 54145 17693 54179
rect 17727 54176 17739 54179
rect 22370 54176 22376 54188
rect 17727 54148 22376 54176
rect 17727 54145 17739 54148
rect 17681 54139 17739 54145
rect 22370 54136 22376 54148
rect 22428 54136 22434 54188
rect 8662 54068 8668 54120
rect 8720 54068 8726 54120
rect 17865 54111 17923 54117
rect 17865 54077 17877 54111
rect 17911 54108 17923 54111
rect 23382 54108 23388 54120
rect 17911 54080 23388 54108
rect 17911 54077 17923 54080
rect 17865 54071 17923 54077
rect 17402 54000 17408 54052
rect 17460 54000 17466 54052
rect 13814 53932 13820 53984
rect 13872 53972 13878 53984
rect 17880 53972 17908 54071
rect 23382 54068 23388 54080
rect 23440 54068 23446 54120
rect 13872 53944 17908 53972
rect 13872 53932 13878 53944
rect 1104 53882 40848 53904
rect 1104 53830 1950 53882
rect 2002 53830 2014 53882
rect 2066 53830 2078 53882
rect 2130 53830 2142 53882
rect 2194 53830 2206 53882
rect 2258 53830 6950 53882
rect 7002 53830 7014 53882
rect 7066 53830 7078 53882
rect 7130 53830 7142 53882
rect 7194 53830 7206 53882
rect 7258 53830 11950 53882
rect 12002 53830 12014 53882
rect 12066 53830 12078 53882
rect 12130 53830 12142 53882
rect 12194 53830 12206 53882
rect 12258 53830 16950 53882
rect 17002 53830 17014 53882
rect 17066 53830 17078 53882
rect 17130 53830 17142 53882
rect 17194 53830 17206 53882
rect 17258 53830 21950 53882
rect 22002 53830 22014 53882
rect 22066 53830 22078 53882
rect 22130 53830 22142 53882
rect 22194 53830 22206 53882
rect 22258 53830 26950 53882
rect 27002 53830 27014 53882
rect 27066 53830 27078 53882
rect 27130 53830 27142 53882
rect 27194 53830 27206 53882
rect 27258 53830 31950 53882
rect 32002 53830 32014 53882
rect 32066 53830 32078 53882
rect 32130 53830 32142 53882
rect 32194 53830 32206 53882
rect 32258 53830 36950 53882
rect 37002 53830 37014 53882
rect 37066 53830 37078 53882
rect 37130 53830 37142 53882
rect 37194 53830 37206 53882
rect 37258 53830 40848 53882
rect 1104 53808 40848 53830
rect 38286 53768 38292 53780
rect 26206 53740 38292 53768
rect 12713 53635 12771 53641
rect 12713 53601 12725 53635
rect 12759 53632 12771 53635
rect 13817 53635 13875 53641
rect 13817 53632 13829 53635
rect 12759 53604 13829 53632
rect 12759 53601 12771 53604
rect 12713 53595 12771 53601
rect 13817 53601 13829 53604
rect 13863 53632 13875 53635
rect 26206 53632 26234 53740
rect 38286 53728 38292 53740
rect 38344 53728 38350 53780
rect 13863 53604 26234 53632
rect 13863 53601 13875 53604
rect 13817 53595 13875 53601
rect 28902 53592 28908 53644
rect 28960 53632 28966 53644
rect 32125 53635 32183 53641
rect 32125 53632 32137 53635
rect 28960 53604 32137 53632
rect 28960 53592 28966 53604
rect 32125 53601 32137 53604
rect 32171 53632 32183 53635
rect 32171 53604 37688 53632
rect 32171 53601 32183 53604
rect 32125 53595 32183 53601
rect 13538 53524 13544 53576
rect 13596 53524 13602 53576
rect 27430 53524 27436 53576
rect 27488 53564 27494 53576
rect 27488 53536 30774 53564
rect 27488 53524 27494 53536
rect 36078 53524 36084 53576
rect 36136 53564 36142 53576
rect 37660 53573 37688 53604
rect 37645 53567 37703 53573
rect 36136 53536 36294 53564
rect 36136 53524 36142 53536
rect 37645 53533 37657 53567
rect 37691 53533 37703 53567
rect 37645 53527 37703 53533
rect 25314 53456 25320 53508
rect 25372 53496 25378 53508
rect 30101 53499 30159 53505
rect 30101 53496 30113 53499
rect 25372 53468 30113 53496
rect 25372 53456 25378 53468
rect 30101 53465 30113 53468
rect 30147 53465 30159 53499
rect 30101 53459 30159 53465
rect 31570 53456 31576 53508
rect 31628 53496 31634 53508
rect 31849 53499 31907 53505
rect 31849 53496 31861 53499
rect 31628 53468 31861 53496
rect 31628 53456 31634 53468
rect 31849 53465 31861 53468
rect 31895 53465 31907 53499
rect 31849 53459 31907 53465
rect 34514 53456 34520 53508
rect 34572 53496 34578 53508
rect 37369 53499 37427 53505
rect 34572 53468 36124 53496
rect 34572 53456 34578 53468
rect 17310 53388 17316 53440
rect 17368 53428 17374 53440
rect 35897 53431 35955 53437
rect 35897 53428 35909 53431
rect 17368 53400 35909 53428
rect 17368 53388 17374 53400
rect 35897 53397 35909 53400
rect 35943 53397 35955 53431
rect 36096 53428 36124 53468
rect 37369 53465 37381 53499
rect 37415 53465 37427 53499
rect 37369 53459 37427 53465
rect 37384 53428 37412 53459
rect 37458 53456 37464 53508
rect 37516 53496 37522 53508
rect 37660 53496 37688 53527
rect 37516 53468 37688 53496
rect 37516 53456 37522 53468
rect 36096 53400 37412 53428
rect 35897 53391 35955 53397
rect 1104 53338 40848 53360
rect 1104 53286 2610 53338
rect 2662 53286 2674 53338
rect 2726 53286 2738 53338
rect 2790 53286 2802 53338
rect 2854 53286 2866 53338
rect 2918 53286 7610 53338
rect 7662 53286 7674 53338
rect 7726 53286 7738 53338
rect 7790 53286 7802 53338
rect 7854 53286 7866 53338
rect 7918 53286 12610 53338
rect 12662 53286 12674 53338
rect 12726 53286 12738 53338
rect 12790 53286 12802 53338
rect 12854 53286 12866 53338
rect 12918 53286 17610 53338
rect 17662 53286 17674 53338
rect 17726 53286 17738 53338
rect 17790 53286 17802 53338
rect 17854 53286 17866 53338
rect 17918 53286 22610 53338
rect 22662 53286 22674 53338
rect 22726 53286 22738 53338
rect 22790 53286 22802 53338
rect 22854 53286 22866 53338
rect 22918 53286 27610 53338
rect 27662 53286 27674 53338
rect 27726 53286 27738 53338
rect 27790 53286 27802 53338
rect 27854 53286 27866 53338
rect 27918 53286 32610 53338
rect 32662 53286 32674 53338
rect 32726 53286 32738 53338
rect 32790 53286 32802 53338
rect 32854 53286 32866 53338
rect 32918 53286 37610 53338
rect 37662 53286 37674 53338
rect 37726 53286 37738 53338
rect 37790 53286 37802 53338
rect 37854 53286 37866 53338
rect 37918 53286 40848 53338
rect 1104 53264 40848 53286
rect 22370 53184 22376 53236
rect 22428 53224 22434 53236
rect 31570 53224 31576 53236
rect 22428 53196 31576 53224
rect 22428 53184 22434 53196
rect 31570 53184 31576 53196
rect 31628 53184 31634 53236
rect 6362 53116 6368 53168
rect 6420 53156 6426 53168
rect 6420 53128 23506 53156
rect 6420 53116 6426 53128
rect 22925 53023 22983 53029
rect 22925 52989 22937 53023
rect 22971 53020 22983 53023
rect 23290 53020 23296 53032
rect 22971 52992 23296 53020
rect 22971 52989 22983 52992
rect 22925 52983 22983 52989
rect 23290 52980 23296 52992
rect 23348 52980 23354 53032
rect 24670 52980 24676 53032
rect 24728 52980 24734 53032
rect 24949 53023 25007 53029
rect 24949 52989 24961 53023
rect 24995 53020 25007 53023
rect 28902 53020 28908 53032
rect 24995 52992 28908 53020
rect 24995 52989 25007 52992
rect 24949 52983 25007 52989
rect 28902 52980 28908 52992
rect 28960 52980 28966 53032
rect 5258 52844 5264 52896
rect 5316 52884 5322 52896
rect 25038 52884 25044 52896
rect 5316 52856 25044 52884
rect 5316 52844 5322 52856
rect 25038 52844 25044 52856
rect 25096 52844 25102 52896
rect 1104 52794 40848 52816
rect 1104 52742 1950 52794
rect 2002 52742 2014 52794
rect 2066 52742 2078 52794
rect 2130 52742 2142 52794
rect 2194 52742 2206 52794
rect 2258 52742 6950 52794
rect 7002 52742 7014 52794
rect 7066 52742 7078 52794
rect 7130 52742 7142 52794
rect 7194 52742 7206 52794
rect 7258 52742 11950 52794
rect 12002 52742 12014 52794
rect 12066 52742 12078 52794
rect 12130 52742 12142 52794
rect 12194 52742 12206 52794
rect 12258 52742 16950 52794
rect 17002 52742 17014 52794
rect 17066 52742 17078 52794
rect 17130 52742 17142 52794
rect 17194 52742 17206 52794
rect 17258 52742 21950 52794
rect 22002 52742 22014 52794
rect 22066 52742 22078 52794
rect 22130 52742 22142 52794
rect 22194 52742 22206 52794
rect 22258 52742 26950 52794
rect 27002 52742 27014 52794
rect 27066 52742 27078 52794
rect 27130 52742 27142 52794
rect 27194 52742 27206 52794
rect 27258 52742 31950 52794
rect 32002 52742 32014 52794
rect 32066 52742 32078 52794
rect 32130 52742 32142 52794
rect 32194 52742 32206 52794
rect 32258 52742 36950 52794
rect 37002 52742 37014 52794
rect 37066 52742 37078 52794
rect 37130 52742 37142 52794
rect 37194 52742 37206 52794
rect 37258 52742 40848 52794
rect 1104 52720 40848 52742
rect 4062 52640 4068 52692
rect 4120 52680 4126 52692
rect 36449 52683 36507 52689
rect 36449 52680 36461 52683
rect 4120 52652 36461 52680
rect 4120 52640 4126 52652
rect 36449 52649 36461 52652
rect 36495 52680 36507 52683
rect 37093 52683 37151 52689
rect 37093 52680 37105 52683
rect 36495 52652 37105 52680
rect 36495 52649 36507 52652
rect 36449 52643 36507 52649
rect 37093 52649 37105 52652
rect 37139 52649 37151 52683
rect 37093 52643 37151 52649
rect 24121 52615 24179 52621
rect 24121 52581 24133 52615
rect 24167 52612 24179 52615
rect 33134 52612 33140 52624
rect 24167 52584 33140 52612
rect 24167 52581 24179 52584
rect 24121 52575 24179 52581
rect 33134 52572 33140 52584
rect 33192 52572 33198 52624
rect 25314 52544 25320 52556
rect 5368 52516 25320 52544
rect 5074 52436 5080 52488
rect 5132 52436 5138 52488
rect 5258 52436 5264 52488
rect 5316 52436 5322 52488
rect 5368 52485 5396 52516
rect 25314 52504 25320 52516
rect 25372 52504 25378 52556
rect 5353 52479 5411 52485
rect 5353 52445 5365 52479
rect 5399 52445 5411 52479
rect 5353 52439 5411 52445
rect 5626 52436 5632 52488
rect 5684 52436 5690 52488
rect 15930 52436 15936 52488
rect 15988 52476 15994 52488
rect 23937 52479 23995 52485
rect 23937 52476 23949 52479
rect 15988 52448 23949 52476
rect 15988 52436 15994 52448
rect 23937 52445 23949 52448
rect 23983 52445 23995 52479
rect 23937 52439 23995 52445
rect 24118 52436 24124 52488
rect 24176 52436 24182 52488
rect 25038 52436 25044 52488
rect 25096 52476 25102 52488
rect 26050 52476 26056 52488
rect 25096 52448 26056 52476
rect 25096 52436 25102 52448
rect 26050 52436 26056 52448
rect 26108 52436 26114 52488
rect 30852 52448 31248 52476
rect 4338 52368 4344 52420
rect 4396 52408 4402 52420
rect 4709 52411 4767 52417
rect 4709 52408 4721 52411
rect 4396 52380 4721 52408
rect 4396 52368 4402 52380
rect 4709 52377 4721 52380
rect 4755 52408 4767 52411
rect 5276 52408 5304 52436
rect 4755 52380 5304 52408
rect 4755 52377 4767 52380
rect 4709 52371 4767 52377
rect 18690 52368 18696 52420
rect 18748 52408 18754 52420
rect 28534 52408 28540 52420
rect 18748 52380 28540 52408
rect 18748 52368 18754 52380
rect 28534 52368 28540 52380
rect 28592 52408 28598 52420
rect 28810 52408 28816 52420
rect 28592 52380 28816 52408
rect 28592 52368 28598 52380
rect 28810 52368 28816 52380
rect 28868 52368 28874 52420
rect 5445 52343 5503 52349
rect 5445 52309 5457 52343
rect 5491 52340 5503 52343
rect 6178 52340 6184 52352
rect 5491 52312 6184 52340
rect 5491 52309 5503 52312
rect 5445 52303 5503 52309
rect 6178 52300 6184 52312
rect 6236 52300 6242 52352
rect 25498 52300 25504 52352
rect 25556 52340 25562 52352
rect 30852 52340 30880 52448
rect 31220 52408 31248 52448
rect 36354 52436 36360 52488
rect 36412 52476 36418 52488
rect 36817 52479 36875 52485
rect 36817 52476 36829 52479
rect 36412 52448 36829 52476
rect 36412 52436 36418 52448
rect 36817 52445 36829 52448
rect 36863 52445 36875 52479
rect 36817 52439 36875 52445
rect 37093 52411 37151 52417
rect 37093 52408 37105 52411
rect 31220 52380 37105 52408
rect 37093 52377 37105 52380
rect 37139 52377 37151 52411
rect 37093 52371 37151 52377
rect 37277 52411 37335 52417
rect 37277 52377 37289 52411
rect 37323 52408 37335 52411
rect 38194 52408 38200 52420
rect 37323 52380 38200 52408
rect 37323 52377 37335 52380
rect 37277 52371 37335 52377
rect 25556 52312 30880 52340
rect 25556 52300 25562 52312
rect 34146 52300 34152 52352
rect 34204 52340 34210 52352
rect 37292 52340 37320 52371
rect 38194 52368 38200 52380
rect 38252 52368 38258 52420
rect 34204 52312 37320 52340
rect 34204 52300 34210 52312
rect 1104 52250 40848 52272
rect 1104 52198 2610 52250
rect 2662 52198 2674 52250
rect 2726 52198 2738 52250
rect 2790 52198 2802 52250
rect 2854 52198 2866 52250
rect 2918 52198 7610 52250
rect 7662 52198 7674 52250
rect 7726 52198 7738 52250
rect 7790 52198 7802 52250
rect 7854 52198 7866 52250
rect 7918 52198 12610 52250
rect 12662 52198 12674 52250
rect 12726 52198 12738 52250
rect 12790 52198 12802 52250
rect 12854 52198 12866 52250
rect 12918 52198 17610 52250
rect 17662 52198 17674 52250
rect 17726 52198 17738 52250
rect 17790 52198 17802 52250
rect 17854 52198 17866 52250
rect 17918 52198 22610 52250
rect 22662 52198 22674 52250
rect 22726 52198 22738 52250
rect 22790 52198 22802 52250
rect 22854 52198 22866 52250
rect 22918 52198 27610 52250
rect 27662 52198 27674 52250
rect 27726 52198 27738 52250
rect 27790 52198 27802 52250
rect 27854 52198 27866 52250
rect 27918 52198 32610 52250
rect 32662 52198 32674 52250
rect 32726 52198 32738 52250
rect 32790 52198 32802 52250
rect 32854 52198 32866 52250
rect 32918 52198 37610 52250
rect 37662 52198 37674 52250
rect 37726 52198 37738 52250
rect 37790 52198 37802 52250
rect 37854 52198 37866 52250
rect 37918 52198 40848 52250
rect 1104 52176 40848 52198
rect 4338 52096 4344 52148
rect 4396 52096 4402 52148
rect 11054 52096 11060 52148
rect 11112 52136 11118 52148
rect 12342 52136 12348 52148
rect 11112 52108 12348 52136
rect 11112 52096 11118 52108
rect 12342 52096 12348 52108
rect 12400 52136 12406 52148
rect 12400 52108 31616 52136
rect 12400 52096 12406 52108
rect 6886 52040 10732 52068
rect 4062 51960 4068 52012
rect 4120 52000 4126 52012
rect 6886 52000 6914 52040
rect 4120 51972 6914 52000
rect 4120 51960 4126 51972
rect 10410 51960 10416 52012
rect 10468 51960 10474 52012
rect 10704 52009 10732 52040
rect 10689 52003 10747 52009
rect 10689 51969 10701 52003
rect 10735 52000 10747 52003
rect 13814 52000 13820 52012
rect 10735 51972 13820 52000
rect 10735 51969 10747 51972
rect 10689 51963 10747 51969
rect 13814 51960 13820 51972
rect 13872 51960 13878 52012
rect 31588 52009 31616 52108
rect 31481 52003 31539 52009
rect 31481 52000 31493 52003
rect 26206 51972 31493 52000
rect 10226 51892 10232 51944
rect 10284 51892 10290 51944
rect 17494 51892 17500 51944
rect 17552 51932 17558 51944
rect 26206 51932 26234 51972
rect 31481 51969 31493 51972
rect 31527 51969 31539 52003
rect 31481 51963 31539 51969
rect 31573 52003 31631 52009
rect 31573 51969 31585 52003
rect 31619 51969 31631 52003
rect 31573 51963 31631 51969
rect 31757 52003 31815 52009
rect 31757 51969 31769 52003
rect 31803 52000 31815 52003
rect 32306 52000 32312 52012
rect 31803 51972 32312 52000
rect 31803 51969 31815 51972
rect 31757 51963 31815 51969
rect 32306 51960 32312 51972
rect 32364 51960 32370 52012
rect 33045 52003 33103 52009
rect 33045 51969 33057 52003
rect 33091 51969 33103 52003
rect 33045 51963 33103 51969
rect 17552 51904 26234 51932
rect 17552 51892 17558 51904
rect 27522 51892 27528 51944
rect 27580 51932 27586 51944
rect 33060 51932 33088 51963
rect 27580 51904 33088 51932
rect 27580 51892 27586 51904
rect 10597 51867 10655 51873
rect 10597 51833 10609 51867
rect 10643 51864 10655 51867
rect 21358 51864 21364 51876
rect 10643 51836 21364 51864
rect 10643 51833 10655 51836
rect 10597 51827 10655 51833
rect 21358 51824 21364 51836
rect 21416 51824 21422 51876
rect 31665 51867 31723 51873
rect 31665 51833 31677 51867
rect 31711 51864 31723 51867
rect 33042 51864 33048 51876
rect 31711 51836 33048 51864
rect 31711 51833 31723 51836
rect 31665 51827 31723 51833
rect 33042 51824 33048 51836
rect 33100 51824 33106 51876
rect 31294 51756 31300 51808
rect 31352 51756 31358 51808
rect 33134 51756 33140 51808
rect 33192 51796 33198 51808
rect 33229 51799 33287 51805
rect 33229 51796 33241 51799
rect 33192 51768 33241 51796
rect 33192 51756 33198 51768
rect 33229 51765 33241 51768
rect 33275 51765 33287 51799
rect 33229 51759 33287 51765
rect 1104 51706 40848 51728
rect 1104 51654 1950 51706
rect 2002 51654 2014 51706
rect 2066 51654 2078 51706
rect 2130 51654 2142 51706
rect 2194 51654 2206 51706
rect 2258 51654 6950 51706
rect 7002 51654 7014 51706
rect 7066 51654 7078 51706
rect 7130 51654 7142 51706
rect 7194 51654 7206 51706
rect 7258 51654 11950 51706
rect 12002 51654 12014 51706
rect 12066 51654 12078 51706
rect 12130 51654 12142 51706
rect 12194 51654 12206 51706
rect 12258 51654 16950 51706
rect 17002 51654 17014 51706
rect 17066 51654 17078 51706
rect 17130 51654 17142 51706
rect 17194 51654 17206 51706
rect 17258 51654 21950 51706
rect 22002 51654 22014 51706
rect 22066 51654 22078 51706
rect 22130 51654 22142 51706
rect 22194 51654 22206 51706
rect 22258 51654 26950 51706
rect 27002 51654 27014 51706
rect 27066 51654 27078 51706
rect 27130 51654 27142 51706
rect 27194 51654 27206 51706
rect 27258 51654 31950 51706
rect 32002 51654 32014 51706
rect 32066 51654 32078 51706
rect 32130 51654 32142 51706
rect 32194 51654 32206 51706
rect 32258 51654 36950 51706
rect 37002 51654 37014 51706
rect 37066 51654 37078 51706
rect 37130 51654 37142 51706
rect 37194 51654 37206 51706
rect 37258 51654 40848 51706
rect 1104 51632 40848 51654
rect 28810 51552 28816 51604
rect 28868 51592 28874 51604
rect 34146 51592 34152 51604
rect 28868 51564 34152 51592
rect 28868 51552 28874 51564
rect 34146 51552 34152 51564
rect 34204 51552 34210 51604
rect 11698 51456 11704 51468
rect 11440 51428 11704 51456
rect 11238 51348 11244 51400
rect 11296 51388 11302 51400
rect 11440 51388 11468 51428
rect 11698 51416 11704 51428
rect 11756 51416 11762 51468
rect 18690 51456 18696 51468
rect 16776 51428 18696 51456
rect 11296 51360 11468 51388
rect 11517 51391 11575 51397
rect 11296 51348 11302 51360
rect 11517 51357 11529 51391
rect 11563 51357 11575 51391
rect 11517 51351 11575 51357
rect 10778 51280 10784 51332
rect 10836 51280 10842 51332
rect 11330 51280 11336 51332
rect 11388 51280 11394 51332
rect 11532 51320 11560 51351
rect 16574 51348 16580 51400
rect 16632 51348 16638 51400
rect 16776 51397 16804 51428
rect 18690 51416 18696 51428
rect 18748 51416 18754 51468
rect 16761 51391 16819 51397
rect 16761 51357 16773 51391
rect 16807 51357 16819 51391
rect 16761 51351 16819 51357
rect 16850 51348 16856 51400
rect 16908 51348 16914 51400
rect 16945 51391 17003 51397
rect 16945 51357 16957 51391
rect 16991 51388 17003 51391
rect 17310 51388 17316 51400
rect 16991 51360 17316 51388
rect 16991 51357 17003 51360
rect 16945 51351 17003 51357
rect 17310 51348 17316 51360
rect 17368 51348 17374 51400
rect 17494 51348 17500 51400
rect 17552 51388 17558 51400
rect 17954 51388 17960 51400
rect 17552 51360 17960 51388
rect 17552 51348 17558 51360
rect 17954 51348 17960 51360
rect 18012 51348 18018 51400
rect 19610 51320 19616 51332
rect 11532 51292 19616 51320
rect 19610 51280 19616 51292
rect 19668 51320 19674 51332
rect 19978 51320 19984 51332
rect 19668 51292 19984 51320
rect 19668 51280 19674 51292
rect 19978 51280 19984 51292
rect 20036 51280 20042 51332
rect 34514 51320 34520 51332
rect 26206 51292 34520 51320
rect 11348 51252 11376 51280
rect 11606 51252 11612 51264
rect 11348 51224 11612 51252
rect 11606 51212 11612 51224
rect 11664 51212 11670 51264
rect 17221 51255 17279 51261
rect 17221 51221 17233 51255
rect 17267 51252 17279 51255
rect 26206 51252 26234 51292
rect 34514 51280 34520 51292
rect 34572 51280 34578 51332
rect 17267 51224 26234 51252
rect 17267 51221 17279 51224
rect 17221 51215 17279 51221
rect 33134 51212 33140 51264
rect 33192 51212 33198 51264
rect 1104 51162 40848 51184
rect 1104 51110 2610 51162
rect 2662 51110 2674 51162
rect 2726 51110 2738 51162
rect 2790 51110 2802 51162
rect 2854 51110 2866 51162
rect 2918 51110 7610 51162
rect 7662 51110 7674 51162
rect 7726 51110 7738 51162
rect 7790 51110 7802 51162
rect 7854 51110 7866 51162
rect 7918 51110 12610 51162
rect 12662 51110 12674 51162
rect 12726 51110 12738 51162
rect 12790 51110 12802 51162
rect 12854 51110 12866 51162
rect 12918 51110 17610 51162
rect 17662 51110 17674 51162
rect 17726 51110 17738 51162
rect 17790 51110 17802 51162
rect 17854 51110 17866 51162
rect 17918 51110 22610 51162
rect 22662 51110 22674 51162
rect 22726 51110 22738 51162
rect 22790 51110 22802 51162
rect 22854 51110 22866 51162
rect 22918 51110 27610 51162
rect 27662 51110 27674 51162
rect 27726 51110 27738 51162
rect 27790 51110 27802 51162
rect 27854 51110 27866 51162
rect 27918 51110 32610 51162
rect 32662 51110 32674 51162
rect 32726 51110 32738 51162
rect 32790 51110 32802 51162
rect 32854 51110 32866 51162
rect 32918 51110 37610 51162
rect 37662 51110 37674 51162
rect 37726 51110 37738 51162
rect 37790 51110 37802 51162
rect 37854 51110 37866 51162
rect 37918 51110 40848 51162
rect 1104 51088 40848 51110
rect 13078 50872 13084 50924
rect 13136 50872 13142 50924
rect 12434 50804 12440 50856
rect 12492 50844 12498 50856
rect 12805 50847 12863 50853
rect 12805 50844 12817 50847
rect 12492 50816 12817 50844
rect 12492 50804 12498 50816
rect 12805 50813 12817 50816
rect 12851 50844 12863 50847
rect 29086 50844 29092 50856
rect 12851 50816 29092 50844
rect 12851 50813 12863 50816
rect 12805 50807 12863 50813
rect 29086 50804 29092 50816
rect 29144 50804 29150 50856
rect 8294 50736 8300 50788
rect 8352 50776 8358 50788
rect 8478 50776 8484 50788
rect 8352 50748 8484 50776
rect 8352 50736 8358 50748
rect 8478 50736 8484 50748
rect 8536 50736 8542 50788
rect 12986 50736 12992 50788
rect 13044 50736 13050 50788
rect 13081 50711 13139 50717
rect 13081 50677 13093 50711
rect 13127 50708 13139 50711
rect 22370 50708 22376 50720
rect 13127 50680 22376 50708
rect 13127 50677 13139 50680
rect 13081 50671 13139 50677
rect 22370 50668 22376 50680
rect 22428 50668 22434 50720
rect 1104 50618 40848 50640
rect 1104 50566 1950 50618
rect 2002 50566 2014 50618
rect 2066 50566 2078 50618
rect 2130 50566 2142 50618
rect 2194 50566 2206 50618
rect 2258 50566 6950 50618
rect 7002 50566 7014 50618
rect 7066 50566 7078 50618
rect 7130 50566 7142 50618
rect 7194 50566 7206 50618
rect 7258 50566 11950 50618
rect 12002 50566 12014 50618
rect 12066 50566 12078 50618
rect 12130 50566 12142 50618
rect 12194 50566 12206 50618
rect 12258 50566 16950 50618
rect 17002 50566 17014 50618
rect 17066 50566 17078 50618
rect 17130 50566 17142 50618
rect 17194 50566 17206 50618
rect 17258 50566 21950 50618
rect 22002 50566 22014 50618
rect 22066 50566 22078 50618
rect 22130 50566 22142 50618
rect 22194 50566 22206 50618
rect 22258 50566 26950 50618
rect 27002 50566 27014 50618
rect 27066 50566 27078 50618
rect 27130 50566 27142 50618
rect 27194 50566 27206 50618
rect 27258 50566 31950 50618
rect 32002 50566 32014 50618
rect 32066 50566 32078 50618
rect 32130 50566 32142 50618
rect 32194 50566 32206 50618
rect 32258 50566 36950 50618
rect 37002 50566 37014 50618
rect 37066 50566 37078 50618
rect 37130 50566 37142 50618
rect 37194 50566 37206 50618
rect 37258 50566 40848 50618
rect 1104 50544 40848 50566
rect 29546 50464 29552 50516
rect 29604 50504 29610 50516
rect 33965 50507 34023 50513
rect 33965 50504 33977 50507
rect 29604 50476 33977 50504
rect 29604 50464 29610 50476
rect 33965 50473 33977 50476
rect 34011 50473 34023 50507
rect 33965 50467 34023 50473
rect 25317 50371 25375 50377
rect 25317 50337 25329 50371
rect 25363 50337 25375 50371
rect 25317 50331 25375 50337
rect 24946 50260 24952 50312
rect 25004 50260 25010 50312
rect 14366 50192 14372 50244
rect 14424 50232 14430 50244
rect 14826 50232 14832 50244
rect 14424 50204 14832 50232
rect 14424 50192 14430 50204
rect 14826 50192 14832 50204
rect 14884 50232 14890 50244
rect 24854 50232 24860 50244
rect 14884 50204 24860 50232
rect 14884 50192 14890 50204
rect 24854 50192 24860 50204
rect 24912 50232 24918 50244
rect 25332 50232 25360 50331
rect 37458 50328 37464 50380
rect 37516 50368 37522 50380
rect 37645 50371 37703 50377
rect 37645 50368 37657 50371
rect 37516 50340 37657 50368
rect 37516 50328 37522 50340
rect 37645 50337 37657 50340
rect 37691 50337 37703 50371
rect 37645 50331 37703 50337
rect 37921 50371 37979 50377
rect 37921 50337 37933 50371
rect 37967 50368 37979 50371
rect 38378 50368 38384 50380
rect 37967 50340 38384 50368
rect 37967 50337 37979 50340
rect 37921 50331 37979 50337
rect 38378 50328 38384 50340
rect 38436 50328 38442 50380
rect 24912 50204 25360 50232
rect 24912 50192 24918 50204
rect 34146 50192 34152 50244
rect 34204 50192 34210 50244
rect 38654 50192 38660 50244
rect 38712 50192 38718 50244
rect 39669 50235 39727 50241
rect 39669 50201 39681 50235
rect 39715 50201 39727 50235
rect 39669 50195 39727 50201
rect 33778 50124 33784 50176
rect 33836 50124 33842 50176
rect 33962 50124 33968 50176
rect 34020 50124 34026 50176
rect 36538 50124 36544 50176
rect 36596 50164 36602 50176
rect 39684 50164 39712 50195
rect 36596 50136 39712 50164
rect 36596 50124 36602 50136
rect 1104 50074 40848 50096
rect 1104 50022 2610 50074
rect 2662 50022 2674 50074
rect 2726 50022 2738 50074
rect 2790 50022 2802 50074
rect 2854 50022 2866 50074
rect 2918 50022 7610 50074
rect 7662 50022 7674 50074
rect 7726 50022 7738 50074
rect 7790 50022 7802 50074
rect 7854 50022 7866 50074
rect 7918 50022 12610 50074
rect 12662 50022 12674 50074
rect 12726 50022 12738 50074
rect 12790 50022 12802 50074
rect 12854 50022 12866 50074
rect 12918 50022 17610 50074
rect 17662 50022 17674 50074
rect 17726 50022 17738 50074
rect 17790 50022 17802 50074
rect 17854 50022 17866 50074
rect 17918 50022 22610 50074
rect 22662 50022 22674 50074
rect 22726 50022 22738 50074
rect 22790 50022 22802 50074
rect 22854 50022 22866 50074
rect 22918 50022 27610 50074
rect 27662 50022 27674 50074
rect 27726 50022 27738 50074
rect 27790 50022 27802 50074
rect 27854 50022 27866 50074
rect 27918 50022 32610 50074
rect 32662 50022 32674 50074
rect 32726 50022 32738 50074
rect 32790 50022 32802 50074
rect 32854 50022 32866 50074
rect 32918 50022 37610 50074
rect 37662 50022 37674 50074
rect 37726 50022 37738 50074
rect 37790 50022 37802 50074
rect 37854 50022 37866 50074
rect 37918 50022 40848 50074
rect 1104 50000 40848 50022
rect 29273 49963 29331 49969
rect 29273 49929 29285 49963
rect 29319 49960 29331 49963
rect 29362 49960 29368 49972
rect 29319 49932 29368 49960
rect 29319 49929 29331 49932
rect 29273 49923 29331 49929
rect 29362 49920 29368 49932
rect 29420 49920 29426 49972
rect 22066 49864 29316 49892
rect 10962 49784 10968 49836
rect 11020 49824 11026 49836
rect 15102 49824 15108 49836
rect 11020 49796 15108 49824
rect 11020 49784 11026 49796
rect 15102 49784 15108 49796
rect 15160 49824 15166 49836
rect 22066 49824 22094 49864
rect 15160 49796 22094 49824
rect 15160 49784 15166 49796
rect 29086 49784 29092 49836
rect 29144 49784 29150 49836
rect 29288 49833 29316 49864
rect 29273 49827 29331 49833
rect 29273 49793 29285 49827
rect 29319 49793 29331 49827
rect 29273 49787 29331 49793
rect 36538 49716 36544 49768
rect 36596 49756 36602 49768
rect 36722 49756 36728 49768
rect 36596 49728 36728 49756
rect 36596 49716 36602 49728
rect 36722 49716 36728 49728
rect 36780 49716 36786 49768
rect 1104 49530 40848 49552
rect 1104 49478 1950 49530
rect 2002 49478 2014 49530
rect 2066 49478 2078 49530
rect 2130 49478 2142 49530
rect 2194 49478 2206 49530
rect 2258 49478 6950 49530
rect 7002 49478 7014 49530
rect 7066 49478 7078 49530
rect 7130 49478 7142 49530
rect 7194 49478 7206 49530
rect 7258 49478 11950 49530
rect 12002 49478 12014 49530
rect 12066 49478 12078 49530
rect 12130 49478 12142 49530
rect 12194 49478 12206 49530
rect 12258 49478 16950 49530
rect 17002 49478 17014 49530
rect 17066 49478 17078 49530
rect 17130 49478 17142 49530
rect 17194 49478 17206 49530
rect 17258 49478 21950 49530
rect 22002 49478 22014 49530
rect 22066 49478 22078 49530
rect 22130 49478 22142 49530
rect 22194 49478 22206 49530
rect 22258 49478 26950 49530
rect 27002 49478 27014 49530
rect 27066 49478 27078 49530
rect 27130 49478 27142 49530
rect 27194 49478 27206 49530
rect 27258 49478 31950 49530
rect 32002 49478 32014 49530
rect 32066 49478 32078 49530
rect 32130 49478 32142 49530
rect 32194 49478 32206 49530
rect 32258 49478 36950 49530
rect 37002 49478 37014 49530
rect 37066 49478 37078 49530
rect 37130 49478 37142 49530
rect 37194 49478 37206 49530
rect 37258 49478 40848 49530
rect 1104 49456 40848 49478
rect 24581 49419 24639 49425
rect 24581 49385 24593 49419
rect 24627 49416 24639 49419
rect 24762 49416 24768 49428
rect 24627 49388 24768 49416
rect 24627 49385 24639 49388
rect 24581 49379 24639 49385
rect 24762 49376 24768 49388
rect 24820 49376 24826 49428
rect 33137 49419 33195 49425
rect 33137 49385 33149 49419
rect 33183 49416 33195 49419
rect 33410 49416 33416 49428
rect 33183 49388 33416 49416
rect 33183 49385 33195 49388
rect 33137 49379 33195 49385
rect 33410 49376 33416 49388
rect 33468 49416 33474 49428
rect 33594 49416 33600 49428
rect 33468 49388 33600 49416
rect 33468 49376 33474 49388
rect 33594 49376 33600 49388
rect 33652 49376 33658 49428
rect 22066 49184 24808 49212
rect 14458 49104 14464 49156
rect 14516 49144 14522 49156
rect 15010 49144 15016 49156
rect 14516 49116 15016 49144
rect 14516 49104 14522 49116
rect 15010 49104 15016 49116
rect 15068 49144 15074 49156
rect 22066 49144 22094 49184
rect 24780 49153 24808 49184
rect 24549 49147 24607 49153
rect 24549 49144 24561 49147
rect 15068 49116 22094 49144
rect 24044 49116 24561 49144
rect 15068 49104 15074 49116
rect 9030 49036 9036 49088
rect 9088 49076 9094 49088
rect 24044 49076 24072 49116
rect 24549 49113 24561 49116
rect 24595 49144 24607 49147
rect 24765 49147 24823 49153
rect 24595 49113 24624 49144
rect 24549 49107 24624 49113
rect 24765 49113 24777 49147
rect 24811 49144 24823 49147
rect 26510 49144 26516 49156
rect 24811 49116 26516 49144
rect 24811 49113 24823 49116
rect 24765 49107 24823 49113
rect 9088 49048 24072 49076
rect 9088 49036 9094 49048
rect 24394 49036 24400 49088
rect 24452 49036 24458 49088
rect 24596 49076 24624 49107
rect 26510 49104 26516 49116
rect 26568 49104 26574 49156
rect 33318 49104 33324 49156
rect 33376 49104 33382 49156
rect 25041 49079 25099 49085
rect 25041 49076 25053 49079
rect 24596 49048 25053 49076
rect 25041 49045 25053 49048
rect 25087 49045 25099 49079
rect 25041 49039 25099 49045
rect 31754 49036 31760 49088
rect 31812 49076 31818 49088
rect 33134 49085 33140 49088
rect 32953 49079 33011 49085
rect 32953 49076 32965 49079
rect 31812 49048 32965 49076
rect 31812 49036 31818 49048
rect 32953 49045 32965 49048
rect 32999 49045 33011 49079
rect 32953 49039 33011 49045
rect 33121 49079 33140 49085
rect 33121 49045 33133 49079
rect 33121 49039 33140 49045
rect 33134 49036 33140 49039
rect 33192 49036 33198 49088
rect 1104 48986 40848 49008
rect 1104 48934 2610 48986
rect 2662 48934 2674 48986
rect 2726 48934 2738 48986
rect 2790 48934 2802 48986
rect 2854 48934 2866 48986
rect 2918 48934 7610 48986
rect 7662 48934 7674 48986
rect 7726 48934 7738 48986
rect 7790 48934 7802 48986
rect 7854 48934 7866 48986
rect 7918 48934 12610 48986
rect 12662 48934 12674 48986
rect 12726 48934 12738 48986
rect 12790 48934 12802 48986
rect 12854 48934 12866 48986
rect 12918 48934 17610 48986
rect 17662 48934 17674 48986
rect 17726 48934 17738 48986
rect 17790 48934 17802 48986
rect 17854 48934 17866 48986
rect 17918 48934 22610 48986
rect 22662 48934 22674 48986
rect 22726 48934 22738 48986
rect 22790 48934 22802 48986
rect 22854 48934 22866 48986
rect 22918 48934 27610 48986
rect 27662 48934 27674 48986
rect 27726 48934 27738 48986
rect 27790 48934 27802 48986
rect 27854 48934 27866 48986
rect 27918 48934 32610 48986
rect 32662 48934 32674 48986
rect 32726 48934 32738 48986
rect 32790 48934 32802 48986
rect 32854 48934 32866 48986
rect 32918 48934 37610 48986
rect 37662 48934 37674 48986
rect 37726 48934 37738 48986
rect 37790 48934 37802 48986
rect 37854 48934 37866 48986
rect 37918 48934 40848 48986
rect 1104 48912 40848 48934
rect 9398 48696 9404 48748
rect 9456 48736 9462 48748
rect 11149 48739 11207 48745
rect 11149 48736 11161 48739
rect 9456 48708 11161 48736
rect 9456 48696 9462 48708
rect 11149 48705 11161 48708
rect 11195 48705 11207 48739
rect 11149 48699 11207 48705
rect 11333 48739 11391 48745
rect 11333 48705 11345 48739
rect 11379 48736 11391 48739
rect 12434 48736 12440 48748
rect 11379 48708 12440 48736
rect 11379 48705 11391 48708
rect 11333 48699 11391 48705
rect 12434 48696 12440 48708
rect 12492 48696 12498 48748
rect 21634 48696 21640 48748
rect 21692 48696 21698 48748
rect 4982 48492 4988 48544
rect 5040 48532 5046 48544
rect 11149 48535 11207 48541
rect 11149 48532 11161 48535
rect 5040 48504 11161 48532
rect 5040 48492 5046 48504
rect 11149 48501 11161 48504
rect 11195 48501 11207 48535
rect 11149 48495 11207 48501
rect 20990 48492 20996 48544
rect 21048 48532 21054 48544
rect 21453 48535 21511 48541
rect 21453 48532 21465 48535
rect 21048 48504 21465 48532
rect 21048 48492 21054 48504
rect 21453 48501 21465 48504
rect 21499 48501 21511 48535
rect 21453 48495 21511 48501
rect 1104 48442 40848 48464
rect 1104 48390 1950 48442
rect 2002 48390 2014 48442
rect 2066 48390 2078 48442
rect 2130 48390 2142 48442
rect 2194 48390 2206 48442
rect 2258 48390 6950 48442
rect 7002 48390 7014 48442
rect 7066 48390 7078 48442
rect 7130 48390 7142 48442
rect 7194 48390 7206 48442
rect 7258 48390 11950 48442
rect 12002 48390 12014 48442
rect 12066 48390 12078 48442
rect 12130 48390 12142 48442
rect 12194 48390 12206 48442
rect 12258 48390 16950 48442
rect 17002 48390 17014 48442
rect 17066 48390 17078 48442
rect 17130 48390 17142 48442
rect 17194 48390 17206 48442
rect 17258 48390 21950 48442
rect 22002 48390 22014 48442
rect 22066 48390 22078 48442
rect 22130 48390 22142 48442
rect 22194 48390 22206 48442
rect 22258 48390 26950 48442
rect 27002 48390 27014 48442
rect 27066 48390 27078 48442
rect 27130 48390 27142 48442
rect 27194 48390 27206 48442
rect 27258 48390 31950 48442
rect 32002 48390 32014 48442
rect 32066 48390 32078 48442
rect 32130 48390 32142 48442
rect 32194 48390 32206 48442
rect 32258 48390 36950 48442
rect 37002 48390 37014 48442
rect 37066 48390 37078 48442
rect 37130 48390 37142 48442
rect 37194 48390 37206 48442
rect 37258 48390 40848 48442
rect 1104 48368 40848 48390
rect 26510 48288 26516 48340
rect 26568 48328 26574 48340
rect 33410 48328 33416 48340
rect 26568 48300 33416 48328
rect 26568 48288 26574 48300
rect 33410 48288 33416 48300
rect 33468 48288 33474 48340
rect 25774 48260 25780 48272
rect 6886 48232 25780 48260
rect 3418 48192 3424 48204
rect 2424 48164 3424 48192
rect 2424 48133 2452 48164
rect 3418 48152 3424 48164
rect 3476 48192 3482 48204
rect 4062 48192 4068 48204
rect 3476 48164 4068 48192
rect 3476 48152 3482 48164
rect 4062 48152 4068 48164
rect 4120 48152 4126 48204
rect 2409 48127 2467 48133
rect 2409 48093 2421 48127
rect 2455 48093 2467 48127
rect 2409 48087 2467 48093
rect 2685 48127 2743 48133
rect 2685 48093 2697 48127
rect 2731 48124 2743 48127
rect 6886 48124 6914 48232
rect 25774 48220 25780 48232
rect 25832 48220 25838 48272
rect 33594 48152 33600 48204
rect 33652 48192 33658 48204
rect 34425 48195 34483 48201
rect 34425 48192 34437 48195
rect 33652 48164 34437 48192
rect 33652 48152 33658 48164
rect 34425 48161 34437 48164
rect 34471 48161 34483 48195
rect 34425 48155 34483 48161
rect 2731 48096 6914 48124
rect 2731 48093 2743 48096
rect 2685 48087 2743 48093
rect 30374 48084 30380 48136
rect 30432 48084 30438 48136
rect 33870 48084 33876 48136
rect 33928 48084 33934 48136
rect 33965 48127 34023 48133
rect 33965 48093 33977 48127
rect 34011 48093 34023 48127
rect 33965 48087 34023 48093
rect 2869 48059 2927 48065
rect 2869 48025 2881 48059
rect 2915 48056 2927 48059
rect 15930 48056 15936 48068
rect 2915 48028 15936 48056
rect 2915 48025 2927 48028
rect 2869 48019 2927 48025
rect 15930 48016 15936 48028
rect 15988 48016 15994 48068
rect 29730 48016 29736 48068
rect 29788 48016 29794 48068
rect 33980 48056 34008 48087
rect 33520 48028 34008 48056
rect 6086 47948 6092 48000
rect 6144 47988 6150 48000
rect 6822 47988 6828 48000
rect 6144 47960 6828 47988
rect 6144 47948 6150 47960
rect 6822 47948 6828 47960
rect 6880 47988 6886 48000
rect 33520 47997 33548 48028
rect 33505 47991 33563 47997
rect 33505 47988 33517 47991
rect 6880 47960 33517 47988
rect 6880 47948 6886 47960
rect 33505 47957 33517 47960
rect 33551 47957 33563 47991
rect 33505 47951 33563 47957
rect 1104 47898 40848 47920
rect 1104 47846 2610 47898
rect 2662 47846 2674 47898
rect 2726 47846 2738 47898
rect 2790 47846 2802 47898
rect 2854 47846 2866 47898
rect 2918 47846 7610 47898
rect 7662 47846 7674 47898
rect 7726 47846 7738 47898
rect 7790 47846 7802 47898
rect 7854 47846 7866 47898
rect 7918 47846 12610 47898
rect 12662 47846 12674 47898
rect 12726 47846 12738 47898
rect 12790 47846 12802 47898
rect 12854 47846 12866 47898
rect 12918 47846 17610 47898
rect 17662 47846 17674 47898
rect 17726 47846 17738 47898
rect 17790 47846 17802 47898
rect 17854 47846 17866 47898
rect 17918 47846 22610 47898
rect 22662 47846 22674 47898
rect 22726 47846 22738 47898
rect 22790 47846 22802 47898
rect 22854 47846 22866 47898
rect 22918 47846 27610 47898
rect 27662 47846 27674 47898
rect 27726 47846 27738 47898
rect 27790 47846 27802 47898
rect 27854 47846 27866 47898
rect 27918 47846 32610 47898
rect 32662 47846 32674 47898
rect 32726 47846 32738 47898
rect 32790 47846 32802 47898
rect 32854 47846 32866 47898
rect 32918 47846 37610 47898
rect 37662 47846 37674 47898
rect 37726 47846 37738 47898
rect 37790 47846 37802 47898
rect 37854 47846 37866 47898
rect 37918 47846 40848 47898
rect 1104 47824 40848 47846
rect 30374 47608 30380 47660
rect 30432 47648 30438 47660
rect 35253 47651 35311 47657
rect 35253 47648 35265 47651
rect 30432 47620 35265 47648
rect 30432 47608 30438 47620
rect 35253 47617 35265 47620
rect 35299 47648 35311 47651
rect 40218 47648 40224 47660
rect 35299 47620 40224 47648
rect 35299 47617 35311 47620
rect 35253 47611 35311 47617
rect 40218 47608 40224 47620
rect 40276 47608 40282 47660
rect 13814 47540 13820 47592
rect 13872 47580 13878 47592
rect 21450 47580 21456 47592
rect 13872 47552 21456 47580
rect 13872 47540 13878 47552
rect 21450 47540 21456 47552
rect 21508 47540 21514 47592
rect 35158 47404 35164 47456
rect 35216 47404 35222 47456
rect 1104 47354 40848 47376
rect 1104 47302 1950 47354
rect 2002 47302 2014 47354
rect 2066 47302 2078 47354
rect 2130 47302 2142 47354
rect 2194 47302 2206 47354
rect 2258 47302 6950 47354
rect 7002 47302 7014 47354
rect 7066 47302 7078 47354
rect 7130 47302 7142 47354
rect 7194 47302 7206 47354
rect 7258 47302 11950 47354
rect 12002 47302 12014 47354
rect 12066 47302 12078 47354
rect 12130 47302 12142 47354
rect 12194 47302 12206 47354
rect 12258 47302 16950 47354
rect 17002 47302 17014 47354
rect 17066 47302 17078 47354
rect 17130 47302 17142 47354
rect 17194 47302 17206 47354
rect 17258 47302 21950 47354
rect 22002 47302 22014 47354
rect 22066 47302 22078 47354
rect 22130 47302 22142 47354
rect 22194 47302 22206 47354
rect 22258 47302 26950 47354
rect 27002 47302 27014 47354
rect 27066 47302 27078 47354
rect 27130 47302 27142 47354
rect 27194 47302 27206 47354
rect 27258 47302 31950 47354
rect 32002 47302 32014 47354
rect 32066 47302 32078 47354
rect 32130 47302 32142 47354
rect 32194 47302 32206 47354
rect 32258 47302 36950 47354
rect 37002 47302 37014 47354
rect 37066 47302 37078 47354
rect 37130 47302 37142 47354
rect 37194 47302 37206 47354
rect 37258 47302 40848 47354
rect 1104 47280 40848 47302
rect 36725 47243 36783 47249
rect 36725 47209 36737 47243
rect 36771 47240 36783 47243
rect 37461 47243 37519 47249
rect 37461 47240 37473 47243
rect 36771 47212 37473 47240
rect 36771 47209 36783 47212
rect 36725 47203 36783 47209
rect 37461 47209 37473 47212
rect 37507 47240 37519 47243
rect 38102 47240 38108 47252
rect 37507 47212 38108 47240
rect 37507 47209 37519 47212
rect 37461 47203 37519 47209
rect 38102 47200 38108 47212
rect 38160 47200 38166 47252
rect 33042 47132 33048 47184
rect 33100 47172 33106 47184
rect 37001 47175 37059 47181
rect 37001 47172 37013 47175
rect 33100 47144 37013 47172
rect 33100 47132 33106 47144
rect 37001 47141 37013 47144
rect 37047 47141 37059 47175
rect 37001 47135 37059 47141
rect 10597 47107 10655 47113
rect 10597 47073 10609 47107
rect 10643 47104 10655 47107
rect 13814 47104 13820 47116
rect 10643 47076 13820 47104
rect 10643 47073 10655 47076
rect 10597 47067 10655 47073
rect 13814 47064 13820 47076
rect 13872 47064 13878 47116
rect 25406 47064 25412 47116
rect 25464 47104 25470 47116
rect 25774 47104 25780 47116
rect 25464 47076 25780 47104
rect 25464 47064 25470 47076
rect 25774 47064 25780 47076
rect 25832 47064 25838 47116
rect 37737 47107 37795 47113
rect 37737 47104 37749 47107
rect 37200 47076 37749 47104
rect 1670 46996 1676 47048
rect 1728 46996 1734 47048
rect 10318 46996 10324 47048
rect 10376 47036 10382 47048
rect 10965 47039 11023 47045
rect 10965 47036 10977 47039
rect 10376 47008 10977 47036
rect 10376 46996 10382 47008
rect 10965 47005 10977 47008
rect 11011 47036 11023 47039
rect 30374 47036 30380 47048
rect 11011 47008 30380 47036
rect 11011 47005 11023 47008
rect 10965 46999 11023 47005
rect 30374 46996 30380 47008
rect 30432 46996 30438 47048
rect 30466 46996 30472 47048
rect 30524 47036 30530 47048
rect 37200 47045 37228 47076
rect 37737 47073 37749 47076
rect 37783 47073 37795 47107
rect 37737 47067 37795 47073
rect 37185 47039 37243 47045
rect 37185 47036 37197 47039
rect 30524 47008 37197 47036
rect 30524 46996 30530 47008
rect 37185 47005 37197 47008
rect 37231 47005 37243 47039
rect 37185 46999 37243 47005
rect 37277 47039 37335 47045
rect 37277 47005 37289 47039
rect 37323 47036 37335 47039
rect 38194 47036 38200 47048
rect 37323 47008 38200 47036
rect 37323 47005 37335 47008
rect 37277 46999 37335 47005
rect 38194 46996 38200 47008
rect 38252 46996 38258 47048
rect 19886 46928 19892 46980
rect 19944 46968 19950 46980
rect 36265 46971 36323 46977
rect 36265 46968 36277 46971
rect 19944 46940 36277 46968
rect 19944 46928 19950 46940
rect 36265 46937 36277 46940
rect 36311 46968 36323 46971
rect 37461 46971 37519 46977
rect 37461 46968 37473 46971
rect 36311 46940 37473 46968
rect 36311 46937 36323 46940
rect 36265 46931 36323 46937
rect 37461 46937 37473 46940
rect 37507 46937 37519 46971
rect 37461 46931 37519 46937
rect 1854 46860 1860 46912
rect 1912 46860 1918 46912
rect 1104 46810 40848 46832
rect 1104 46758 2610 46810
rect 2662 46758 2674 46810
rect 2726 46758 2738 46810
rect 2790 46758 2802 46810
rect 2854 46758 2866 46810
rect 2918 46758 7610 46810
rect 7662 46758 7674 46810
rect 7726 46758 7738 46810
rect 7790 46758 7802 46810
rect 7854 46758 7866 46810
rect 7918 46758 12610 46810
rect 12662 46758 12674 46810
rect 12726 46758 12738 46810
rect 12790 46758 12802 46810
rect 12854 46758 12866 46810
rect 12918 46758 17610 46810
rect 17662 46758 17674 46810
rect 17726 46758 17738 46810
rect 17790 46758 17802 46810
rect 17854 46758 17866 46810
rect 17918 46758 22610 46810
rect 22662 46758 22674 46810
rect 22726 46758 22738 46810
rect 22790 46758 22802 46810
rect 22854 46758 22866 46810
rect 22918 46758 27610 46810
rect 27662 46758 27674 46810
rect 27726 46758 27738 46810
rect 27790 46758 27802 46810
rect 27854 46758 27866 46810
rect 27918 46758 32610 46810
rect 32662 46758 32674 46810
rect 32726 46758 32738 46810
rect 32790 46758 32802 46810
rect 32854 46758 32866 46810
rect 32918 46758 37610 46810
rect 37662 46758 37674 46810
rect 37726 46758 37738 46810
rect 37790 46758 37802 46810
rect 37854 46758 37866 46810
rect 37918 46758 40848 46810
rect 1104 46736 40848 46758
rect 28810 46520 28816 46572
rect 28868 46520 28874 46572
rect 28902 46316 28908 46368
rect 28960 46356 28966 46368
rect 30101 46359 30159 46365
rect 30101 46356 30113 46359
rect 28960 46328 30113 46356
rect 28960 46316 28966 46328
rect 30101 46325 30113 46328
rect 30147 46325 30159 46359
rect 30101 46319 30159 46325
rect 1104 46266 40848 46288
rect 1104 46214 1950 46266
rect 2002 46214 2014 46266
rect 2066 46214 2078 46266
rect 2130 46214 2142 46266
rect 2194 46214 2206 46266
rect 2258 46214 6950 46266
rect 7002 46214 7014 46266
rect 7066 46214 7078 46266
rect 7130 46214 7142 46266
rect 7194 46214 7206 46266
rect 7258 46214 11950 46266
rect 12002 46214 12014 46266
rect 12066 46214 12078 46266
rect 12130 46214 12142 46266
rect 12194 46214 12206 46266
rect 12258 46214 16950 46266
rect 17002 46214 17014 46266
rect 17066 46214 17078 46266
rect 17130 46214 17142 46266
rect 17194 46214 17206 46266
rect 17258 46214 21950 46266
rect 22002 46214 22014 46266
rect 22066 46214 22078 46266
rect 22130 46214 22142 46266
rect 22194 46214 22206 46266
rect 22258 46214 26950 46266
rect 27002 46214 27014 46266
rect 27066 46214 27078 46266
rect 27130 46214 27142 46266
rect 27194 46214 27206 46266
rect 27258 46214 31950 46266
rect 32002 46214 32014 46266
rect 32066 46214 32078 46266
rect 32130 46214 32142 46266
rect 32194 46214 32206 46266
rect 32258 46214 36950 46266
rect 37002 46214 37014 46266
rect 37066 46214 37078 46266
rect 37130 46214 37142 46266
rect 37194 46214 37206 46266
rect 37258 46214 40848 46266
rect 1104 46192 40848 46214
rect 26329 46155 26387 46161
rect 26329 46121 26341 46155
rect 26375 46152 26387 46155
rect 34606 46152 34612 46164
rect 26375 46124 34612 46152
rect 26375 46121 26387 46124
rect 26329 46115 26387 46121
rect 34606 46112 34612 46124
rect 34664 46112 34670 46164
rect 9582 45908 9588 45960
rect 9640 45948 9646 45960
rect 14185 45951 14243 45957
rect 14185 45948 14197 45951
rect 9640 45920 14197 45948
rect 9640 45908 9646 45920
rect 14185 45917 14197 45920
rect 14231 45948 14243 45951
rect 16117 45951 16175 45957
rect 16117 45948 16129 45951
rect 14231 45920 16129 45948
rect 14231 45917 14243 45920
rect 14185 45911 14243 45917
rect 16117 45917 16129 45920
rect 16163 45917 16175 45951
rect 18601 45951 18659 45957
rect 18601 45948 18613 45951
rect 16117 45911 16175 45917
rect 16546 45920 18613 45948
rect 14550 45840 14556 45892
rect 14608 45840 14614 45892
rect 15378 45840 15384 45892
rect 15436 45880 15442 45892
rect 16546 45880 16574 45920
rect 18601 45917 18613 45920
rect 18647 45948 18659 45951
rect 29730 45948 29736 45960
rect 18647 45920 29736 45948
rect 18647 45917 18659 45920
rect 18601 45911 18659 45917
rect 29730 45908 29736 45920
rect 29788 45908 29794 45960
rect 15436 45852 16574 45880
rect 15436 45840 15442 45852
rect 23014 45840 23020 45892
rect 23072 45880 23078 45892
rect 26329 45883 26387 45889
rect 26329 45880 26341 45883
rect 23072 45852 26341 45880
rect 23072 45840 23078 45852
rect 26329 45849 26341 45852
rect 26375 45849 26387 45883
rect 26329 45843 26387 45849
rect 26510 45840 26516 45892
rect 26568 45840 26574 45892
rect 28902 45840 28908 45892
rect 28960 45840 28966 45892
rect 18690 45772 18696 45824
rect 18748 45772 18754 45824
rect 25958 45772 25964 45824
rect 26016 45812 26022 45824
rect 26145 45815 26203 45821
rect 26145 45812 26157 45815
rect 26016 45784 26157 45812
rect 26016 45772 26022 45784
rect 26145 45781 26157 45784
rect 26191 45781 26203 45815
rect 26145 45775 26203 45781
rect 1104 45722 40848 45744
rect 1104 45670 2610 45722
rect 2662 45670 2674 45722
rect 2726 45670 2738 45722
rect 2790 45670 2802 45722
rect 2854 45670 2866 45722
rect 2918 45670 7610 45722
rect 7662 45670 7674 45722
rect 7726 45670 7738 45722
rect 7790 45670 7802 45722
rect 7854 45670 7866 45722
rect 7918 45670 12610 45722
rect 12662 45670 12674 45722
rect 12726 45670 12738 45722
rect 12790 45670 12802 45722
rect 12854 45670 12866 45722
rect 12918 45670 17610 45722
rect 17662 45670 17674 45722
rect 17726 45670 17738 45722
rect 17790 45670 17802 45722
rect 17854 45670 17866 45722
rect 17918 45670 22610 45722
rect 22662 45670 22674 45722
rect 22726 45670 22738 45722
rect 22790 45670 22802 45722
rect 22854 45670 22866 45722
rect 22918 45670 27610 45722
rect 27662 45670 27674 45722
rect 27726 45670 27738 45722
rect 27790 45670 27802 45722
rect 27854 45670 27866 45722
rect 27918 45670 32610 45722
rect 32662 45670 32674 45722
rect 32726 45670 32738 45722
rect 32790 45670 32802 45722
rect 32854 45670 32866 45722
rect 32918 45670 37610 45722
rect 37662 45670 37674 45722
rect 37726 45670 37738 45722
rect 37790 45670 37802 45722
rect 37854 45670 37866 45722
rect 37918 45670 40848 45722
rect 1104 45648 40848 45670
rect 8294 45568 8300 45620
rect 8352 45608 8358 45620
rect 9582 45608 9588 45620
rect 8352 45580 9588 45608
rect 8352 45568 8358 45580
rect 9582 45568 9588 45580
rect 9640 45568 9646 45620
rect 3050 45500 3056 45552
rect 3108 45540 3114 45552
rect 14826 45540 14832 45552
rect 3108 45512 14832 45540
rect 3108 45500 3114 45512
rect 14826 45500 14832 45512
rect 14884 45500 14890 45552
rect 3421 45475 3479 45481
rect 1394 45364 1400 45416
rect 1452 45364 1458 45416
rect 2056 45268 2084 45458
rect 3421 45441 3433 45475
rect 3467 45472 3479 45475
rect 8294 45472 8300 45484
rect 3467 45444 8300 45472
rect 3467 45441 3479 45444
rect 3421 45435 3479 45441
rect 8294 45432 8300 45444
rect 8352 45432 8358 45484
rect 16850 45432 16856 45484
rect 16908 45472 16914 45484
rect 25041 45475 25099 45481
rect 25041 45472 25053 45475
rect 16908 45444 25053 45472
rect 16908 45432 16914 45444
rect 25041 45441 25053 45444
rect 25087 45441 25099 45475
rect 25041 45435 25099 45441
rect 3142 45364 3148 45416
rect 3200 45364 3206 45416
rect 14274 45364 14280 45416
rect 14332 45404 14338 45416
rect 24949 45407 25007 45413
rect 24949 45404 24961 45407
rect 14332 45376 24961 45404
rect 14332 45364 14338 45376
rect 24949 45373 24961 45376
rect 24995 45373 25007 45407
rect 24949 45367 25007 45373
rect 35158 45336 35164 45348
rect 21376 45308 35164 45336
rect 3789 45271 3847 45277
rect 3789 45268 3801 45271
rect 2056 45240 3801 45268
rect 3789 45237 3801 45240
rect 3835 45268 3847 45271
rect 21376 45268 21404 45308
rect 35158 45296 35164 45308
rect 35216 45296 35222 45348
rect 3835 45240 21404 45268
rect 3835 45237 3847 45240
rect 3789 45231 3847 45237
rect 1104 45178 40848 45200
rect 1104 45126 1950 45178
rect 2002 45126 2014 45178
rect 2066 45126 2078 45178
rect 2130 45126 2142 45178
rect 2194 45126 2206 45178
rect 2258 45126 6950 45178
rect 7002 45126 7014 45178
rect 7066 45126 7078 45178
rect 7130 45126 7142 45178
rect 7194 45126 7206 45178
rect 7258 45126 11950 45178
rect 12002 45126 12014 45178
rect 12066 45126 12078 45178
rect 12130 45126 12142 45178
rect 12194 45126 12206 45178
rect 12258 45126 16950 45178
rect 17002 45126 17014 45178
rect 17066 45126 17078 45178
rect 17130 45126 17142 45178
rect 17194 45126 17206 45178
rect 17258 45126 21950 45178
rect 22002 45126 22014 45178
rect 22066 45126 22078 45178
rect 22130 45126 22142 45178
rect 22194 45126 22206 45178
rect 22258 45126 26950 45178
rect 27002 45126 27014 45178
rect 27066 45126 27078 45178
rect 27130 45126 27142 45178
rect 27194 45126 27206 45178
rect 27258 45126 31950 45178
rect 32002 45126 32014 45178
rect 32066 45126 32078 45178
rect 32130 45126 32142 45178
rect 32194 45126 32206 45178
rect 32258 45126 36950 45178
rect 37002 45126 37014 45178
rect 37066 45126 37078 45178
rect 37130 45126 37142 45178
rect 37194 45126 37206 45178
rect 37258 45126 40848 45178
rect 1104 45104 40848 45126
rect 1394 45024 1400 45076
rect 1452 45064 1458 45076
rect 10410 45064 10416 45076
rect 1452 45036 10416 45064
rect 1452 45024 1458 45036
rect 10410 45024 10416 45036
rect 10468 45024 10474 45076
rect 5350 44996 5356 45008
rect 2884 44968 5356 44996
rect 2884 44869 2912 44968
rect 5350 44956 5356 44968
rect 5408 44996 5414 45008
rect 19426 44996 19432 45008
rect 5408 44968 19432 44996
rect 5408 44956 5414 44968
rect 19426 44956 19432 44968
rect 19484 44956 19490 45008
rect 2961 44931 3019 44937
rect 2961 44897 2973 44931
rect 3007 44928 3019 44931
rect 3050 44928 3056 44940
rect 3007 44900 3056 44928
rect 3007 44897 3019 44900
rect 2961 44891 3019 44897
rect 3050 44888 3056 44900
rect 3108 44888 3114 44940
rect 3145 44931 3203 44937
rect 3145 44897 3157 44931
rect 3191 44897 3203 44931
rect 3145 44891 3203 44897
rect 3329 44931 3387 44937
rect 3329 44897 3341 44931
rect 3375 44928 3387 44931
rect 5534 44928 5540 44940
rect 3375 44900 5540 44928
rect 3375 44897 3387 44900
rect 3329 44891 3387 44897
rect 2869 44863 2927 44869
rect 2869 44829 2881 44863
rect 2915 44829 2927 44863
rect 2869 44823 2927 44829
rect 2498 44752 2504 44804
rect 2556 44792 2562 44804
rect 2685 44795 2743 44801
rect 2685 44792 2697 44795
rect 2556 44764 2697 44792
rect 2556 44752 2562 44764
rect 2685 44761 2697 44764
rect 2731 44761 2743 44795
rect 3160 44792 3188 44891
rect 5534 44888 5540 44900
rect 5592 44888 5598 44940
rect 10410 44888 10416 44940
rect 10468 44928 10474 44940
rect 20898 44928 20904 44940
rect 10468 44900 20904 44928
rect 10468 44888 10474 44900
rect 20898 44888 20904 44900
rect 20956 44888 20962 44940
rect 35986 44928 35992 44940
rect 22572 44900 35992 44928
rect 3237 44863 3295 44869
rect 5258 44864 5264 44872
rect 3237 44829 3249 44863
rect 3283 44860 3295 44863
rect 5092 44860 5264 44864
rect 3283 44836 5264 44860
rect 3283 44832 5120 44836
rect 3283 44829 3295 44832
rect 3237 44823 3295 44829
rect 5258 44820 5264 44836
rect 5316 44820 5322 44872
rect 5718 44860 5724 44872
rect 5368 44832 5724 44860
rect 3160 44764 3372 44792
rect 2685 44755 2743 44761
rect 3344 44724 3372 44764
rect 5368 44724 5396 44832
rect 5718 44820 5724 44832
rect 5776 44820 5782 44872
rect 19426 44820 19432 44872
rect 19484 44860 19490 44872
rect 22572 44869 22600 44900
rect 35986 44888 35992 44900
rect 36044 44888 36050 44940
rect 22557 44863 22615 44869
rect 22557 44860 22569 44863
rect 19484 44832 22569 44860
rect 19484 44820 19490 44832
rect 22557 44829 22569 44832
rect 22603 44829 22615 44863
rect 22557 44823 22615 44829
rect 22833 44863 22891 44869
rect 22833 44829 22845 44863
rect 22879 44860 22891 44863
rect 30558 44860 30564 44872
rect 22879 44832 30564 44860
rect 22879 44829 22891 44832
rect 22833 44823 22891 44829
rect 30558 44820 30564 44832
rect 30616 44820 30622 44872
rect 5442 44752 5448 44804
rect 5500 44792 5506 44804
rect 8478 44792 8484 44804
rect 5500 44764 8484 44792
rect 5500 44752 5506 44764
rect 8478 44752 8484 44764
rect 8536 44752 8542 44804
rect 22278 44792 22284 44804
rect 16546 44764 22284 44792
rect 3344 44696 5396 44724
rect 5534 44684 5540 44736
rect 5592 44724 5598 44736
rect 16546 44724 16574 44764
rect 22278 44752 22284 44764
rect 22336 44792 22342 44804
rect 22462 44792 22468 44804
rect 22336 44764 22468 44792
rect 22336 44752 22342 44764
rect 22462 44752 22468 44764
rect 22520 44792 22526 44804
rect 22741 44795 22799 44801
rect 22741 44792 22753 44795
rect 22520 44764 22753 44792
rect 22520 44752 22526 44764
rect 22741 44761 22753 44764
rect 22787 44761 22799 44795
rect 22741 44755 22799 44761
rect 5592 44696 16574 44724
rect 5592 44684 5598 44696
rect 22370 44684 22376 44736
rect 22428 44684 22434 44736
rect 1104 44634 40848 44656
rect 1104 44582 2610 44634
rect 2662 44582 2674 44634
rect 2726 44582 2738 44634
rect 2790 44582 2802 44634
rect 2854 44582 2866 44634
rect 2918 44582 7610 44634
rect 7662 44582 7674 44634
rect 7726 44582 7738 44634
rect 7790 44582 7802 44634
rect 7854 44582 7866 44634
rect 7918 44582 12610 44634
rect 12662 44582 12674 44634
rect 12726 44582 12738 44634
rect 12790 44582 12802 44634
rect 12854 44582 12866 44634
rect 12918 44582 17610 44634
rect 17662 44582 17674 44634
rect 17726 44582 17738 44634
rect 17790 44582 17802 44634
rect 17854 44582 17866 44634
rect 17918 44582 22610 44634
rect 22662 44582 22674 44634
rect 22726 44582 22738 44634
rect 22790 44582 22802 44634
rect 22854 44582 22866 44634
rect 22918 44582 27610 44634
rect 27662 44582 27674 44634
rect 27726 44582 27738 44634
rect 27790 44582 27802 44634
rect 27854 44582 27866 44634
rect 27918 44582 32610 44634
rect 32662 44582 32674 44634
rect 32726 44582 32738 44634
rect 32790 44582 32802 44634
rect 32854 44582 32866 44634
rect 32918 44582 37610 44634
rect 37662 44582 37674 44634
rect 37726 44582 37738 44634
rect 37790 44582 37802 44634
rect 37854 44582 37866 44634
rect 37918 44582 40848 44634
rect 1104 44560 40848 44582
rect 14274 44140 14280 44192
rect 14332 44180 14338 44192
rect 14642 44180 14648 44192
rect 14332 44152 14648 44180
rect 14332 44140 14338 44152
rect 14642 44140 14648 44152
rect 14700 44140 14706 44192
rect 16850 44140 16856 44192
rect 16908 44180 16914 44192
rect 17310 44180 17316 44192
rect 16908 44152 17316 44180
rect 16908 44140 16914 44152
rect 17310 44140 17316 44152
rect 17368 44140 17374 44192
rect 1104 44090 40848 44112
rect 1104 44038 1950 44090
rect 2002 44038 2014 44090
rect 2066 44038 2078 44090
rect 2130 44038 2142 44090
rect 2194 44038 2206 44090
rect 2258 44038 6950 44090
rect 7002 44038 7014 44090
rect 7066 44038 7078 44090
rect 7130 44038 7142 44090
rect 7194 44038 7206 44090
rect 7258 44038 11950 44090
rect 12002 44038 12014 44090
rect 12066 44038 12078 44090
rect 12130 44038 12142 44090
rect 12194 44038 12206 44090
rect 12258 44038 16950 44090
rect 17002 44038 17014 44090
rect 17066 44038 17078 44090
rect 17130 44038 17142 44090
rect 17194 44038 17206 44090
rect 17258 44038 21950 44090
rect 22002 44038 22014 44090
rect 22066 44038 22078 44090
rect 22130 44038 22142 44090
rect 22194 44038 22206 44090
rect 22258 44038 26950 44090
rect 27002 44038 27014 44090
rect 27066 44038 27078 44090
rect 27130 44038 27142 44090
rect 27194 44038 27206 44090
rect 27258 44038 31950 44090
rect 32002 44038 32014 44090
rect 32066 44038 32078 44090
rect 32130 44038 32142 44090
rect 32194 44038 32206 44090
rect 32258 44038 36950 44090
rect 37002 44038 37014 44090
rect 37066 44038 37078 44090
rect 37130 44038 37142 44090
rect 37194 44038 37206 44090
rect 37258 44038 40848 44090
rect 1104 44016 40848 44038
rect 24854 43800 24860 43852
rect 24912 43800 24918 43852
rect 25498 43800 25504 43852
rect 25556 43800 25562 43852
rect 24673 43775 24731 43781
rect 24673 43741 24685 43775
rect 24719 43741 24731 43775
rect 24673 43735 24731 43741
rect 25225 43775 25283 43781
rect 25225 43741 25237 43775
rect 25271 43772 25283 43775
rect 28258 43772 28264 43784
rect 25271 43744 28264 43772
rect 25271 43741 25283 43744
rect 25225 43735 25283 43741
rect 24688 43704 24716 43735
rect 28258 43732 28264 43744
rect 28316 43732 28322 43784
rect 29086 43704 29092 43716
rect 24688 43676 29092 43704
rect 29086 43664 29092 43676
rect 29144 43704 29150 43716
rect 29270 43704 29276 43716
rect 29144 43676 29276 43704
rect 29144 43664 29150 43676
rect 29270 43664 29276 43676
rect 29328 43664 29334 43716
rect 4798 43596 4804 43648
rect 4856 43636 4862 43648
rect 24765 43639 24823 43645
rect 24765 43636 24777 43639
rect 4856 43608 24777 43636
rect 4856 43596 4862 43608
rect 24765 43605 24777 43608
rect 24811 43605 24823 43639
rect 24765 43599 24823 43605
rect 1104 43546 40848 43568
rect 1104 43494 2610 43546
rect 2662 43494 2674 43546
rect 2726 43494 2738 43546
rect 2790 43494 2802 43546
rect 2854 43494 2866 43546
rect 2918 43494 7610 43546
rect 7662 43494 7674 43546
rect 7726 43494 7738 43546
rect 7790 43494 7802 43546
rect 7854 43494 7866 43546
rect 7918 43494 12610 43546
rect 12662 43494 12674 43546
rect 12726 43494 12738 43546
rect 12790 43494 12802 43546
rect 12854 43494 12866 43546
rect 12918 43494 17610 43546
rect 17662 43494 17674 43546
rect 17726 43494 17738 43546
rect 17790 43494 17802 43546
rect 17854 43494 17866 43546
rect 17918 43494 22610 43546
rect 22662 43494 22674 43546
rect 22726 43494 22738 43546
rect 22790 43494 22802 43546
rect 22854 43494 22866 43546
rect 22918 43494 27610 43546
rect 27662 43494 27674 43546
rect 27726 43494 27738 43546
rect 27790 43494 27802 43546
rect 27854 43494 27866 43546
rect 27918 43494 32610 43546
rect 32662 43494 32674 43546
rect 32726 43494 32738 43546
rect 32790 43494 32802 43546
rect 32854 43494 32866 43546
rect 32918 43494 37610 43546
rect 37662 43494 37674 43546
rect 37726 43494 37738 43546
rect 37790 43494 37802 43546
rect 37854 43494 37866 43546
rect 37918 43494 40848 43546
rect 1104 43472 40848 43494
rect 1104 43002 40848 43024
rect 1104 42950 1950 43002
rect 2002 42950 2014 43002
rect 2066 42950 2078 43002
rect 2130 42950 2142 43002
rect 2194 42950 2206 43002
rect 2258 42950 6950 43002
rect 7002 42950 7014 43002
rect 7066 42950 7078 43002
rect 7130 42950 7142 43002
rect 7194 42950 7206 43002
rect 7258 42950 11950 43002
rect 12002 42950 12014 43002
rect 12066 42950 12078 43002
rect 12130 42950 12142 43002
rect 12194 42950 12206 43002
rect 12258 42950 16950 43002
rect 17002 42950 17014 43002
rect 17066 42950 17078 43002
rect 17130 42950 17142 43002
rect 17194 42950 17206 43002
rect 17258 42950 21950 43002
rect 22002 42950 22014 43002
rect 22066 42950 22078 43002
rect 22130 42950 22142 43002
rect 22194 42950 22206 43002
rect 22258 42950 26950 43002
rect 27002 42950 27014 43002
rect 27066 42950 27078 43002
rect 27130 42950 27142 43002
rect 27194 42950 27206 43002
rect 27258 42950 31950 43002
rect 32002 42950 32014 43002
rect 32066 42950 32078 43002
rect 32130 42950 32142 43002
rect 32194 42950 32206 43002
rect 32258 42950 36950 43002
rect 37002 42950 37014 43002
rect 37066 42950 37078 43002
rect 37130 42950 37142 43002
rect 37194 42950 37206 43002
rect 37258 42950 40848 43002
rect 1104 42928 40848 42950
rect 1104 42458 40848 42480
rect 1104 42406 2610 42458
rect 2662 42406 2674 42458
rect 2726 42406 2738 42458
rect 2790 42406 2802 42458
rect 2854 42406 2866 42458
rect 2918 42406 7610 42458
rect 7662 42406 7674 42458
rect 7726 42406 7738 42458
rect 7790 42406 7802 42458
rect 7854 42406 7866 42458
rect 7918 42406 12610 42458
rect 12662 42406 12674 42458
rect 12726 42406 12738 42458
rect 12790 42406 12802 42458
rect 12854 42406 12866 42458
rect 12918 42406 17610 42458
rect 17662 42406 17674 42458
rect 17726 42406 17738 42458
rect 17790 42406 17802 42458
rect 17854 42406 17866 42458
rect 17918 42406 22610 42458
rect 22662 42406 22674 42458
rect 22726 42406 22738 42458
rect 22790 42406 22802 42458
rect 22854 42406 22866 42458
rect 22918 42406 27610 42458
rect 27662 42406 27674 42458
rect 27726 42406 27738 42458
rect 27790 42406 27802 42458
rect 27854 42406 27866 42458
rect 27918 42406 32610 42458
rect 32662 42406 32674 42458
rect 32726 42406 32738 42458
rect 32790 42406 32802 42458
rect 32854 42406 32866 42458
rect 32918 42406 37610 42458
rect 37662 42406 37674 42458
rect 37726 42406 37738 42458
rect 37790 42406 37802 42458
rect 37854 42406 37866 42458
rect 37918 42406 40848 42458
rect 1104 42384 40848 42406
rect 1104 41914 40848 41936
rect 1104 41862 1950 41914
rect 2002 41862 2014 41914
rect 2066 41862 2078 41914
rect 2130 41862 2142 41914
rect 2194 41862 2206 41914
rect 2258 41862 6950 41914
rect 7002 41862 7014 41914
rect 7066 41862 7078 41914
rect 7130 41862 7142 41914
rect 7194 41862 7206 41914
rect 7258 41862 11950 41914
rect 12002 41862 12014 41914
rect 12066 41862 12078 41914
rect 12130 41862 12142 41914
rect 12194 41862 12206 41914
rect 12258 41862 16950 41914
rect 17002 41862 17014 41914
rect 17066 41862 17078 41914
rect 17130 41862 17142 41914
rect 17194 41862 17206 41914
rect 17258 41862 21950 41914
rect 22002 41862 22014 41914
rect 22066 41862 22078 41914
rect 22130 41862 22142 41914
rect 22194 41862 22206 41914
rect 22258 41862 26950 41914
rect 27002 41862 27014 41914
rect 27066 41862 27078 41914
rect 27130 41862 27142 41914
rect 27194 41862 27206 41914
rect 27258 41862 31950 41914
rect 32002 41862 32014 41914
rect 32066 41862 32078 41914
rect 32130 41862 32142 41914
rect 32194 41862 32206 41914
rect 32258 41862 36950 41914
rect 37002 41862 37014 41914
rect 37066 41862 37078 41914
rect 37130 41862 37142 41914
rect 37194 41862 37206 41914
rect 37258 41862 40848 41914
rect 1104 41840 40848 41862
rect 13538 41760 13544 41812
rect 13596 41800 13602 41812
rect 36541 41803 36599 41809
rect 36541 41800 36553 41803
rect 13596 41772 36553 41800
rect 13596 41760 13602 41772
rect 36541 41769 36553 41772
rect 36587 41769 36599 41803
rect 36541 41763 36599 41769
rect 26050 41692 26056 41744
rect 26108 41732 26114 41744
rect 30742 41732 30748 41744
rect 26108 41704 30748 41732
rect 26108 41692 26114 41704
rect 30742 41692 30748 41704
rect 30800 41692 30806 41744
rect 24765 41667 24823 41673
rect 24765 41633 24777 41667
rect 24811 41664 24823 41667
rect 28902 41664 28908 41676
rect 24811 41636 28908 41664
rect 24811 41633 24823 41636
rect 24765 41627 24823 41633
rect 28902 41624 28908 41636
rect 28960 41624 28966 41676
rect 30466 41664 30472 41676
rect 29012 41636 30472 41664
rect 13814 41556 13820 41608
rect 13872 41596 13878 41608
rect 14274 41596 14280 41608
rect 13872 41568 14280 41596
rect 13872 41556 13878 41568
rect 14274 41556 14280 41568
rect 14332 41596 14338 41608
rect 14369 41599 14427 41605
rect 14369 41596 14381 41599
rect 14332 41568 14381 41596
rect 14332 41556 14338 41568
rect 14369 41565 14381 41568
rect 14415 41565 14427 41599
rect 14369 41559 14427 41565
rect 14918 41556 14924 41608
rect 14976 41596 14982 41608
rect 15378 41596 15384 41608
rect 14976 41568 15384 41596
rect 14976 41556 14982 41568
rect 15378 41556 15384 41568
rect 15436 41556 15442 41608
rect 26789 41599 26847 41605
rect 26789 41596 26801 41599
rect 26436 41568 26801 41596
rect 25038 41488 25044 41540
rect 25096 41488 25102 41540
rect 26326 41528 26332 41540
rect 26266 41500 26332 41528
rect 26326 41488 26332 41500
rect 26384 41488 26390 41540
rect 5258 41420 5264 41472
rect 5316 41460 5322 41472
rect 14277 41463 14335 41469
rect 14277 41460 14289 41463
rect 5316 41432 14289 41460
rect 5316 41420 5322 41432
rect 14277 41429 14289 41432
rect 14323 41429 14335 41463
rect 14277 41423 14335 41429
rect 15473 41463 15531 41469
rect 15473 41429 15485 41463
rect 15519 41460 15531 41463
rect 15562 41460 15568 41472
rect 15519 41432 15568 41460
rect 15519 41429 15531 41432
rect 15473 41423 15531 41429
rect 15562 41420 15568 41432
rect 15620 41420 15626 41472
rect 19978 41420 19984 41472
rect 20036 41460 20042 41472
rect 26436 41460 26464 41568
rect 26789 41565 26801 41568
rect 26835 41596 26847 41599
rect 29012 41596 29040 41636
rect 30466 41624 30472 41636
rect 30524 41624 30530 41676
rect 36556 41664 36584 41763
rect 37185 41667 37243 41673
rect 37185 41664 37197 41667
rect 36556 41636 37197 41664
rect 37185 41633 37197 41636
rect 37231 41633 37243 41667
rect 37185 41627 37243 41633
rect 36814 41596 36820 41608
rect 26835 41568 29040 41596
rect 31726 41568 36820 41596
rect 26835 41565 26847 41568
rect 26789 41559 26847 41565
rect 26694 41488 26700 41540
rect 26752 41528 26758 41540
rect 27982 41528 27988 41540
rect 26752 41500 27988 41528
rect 26752 41488 26758 41500
rect 27982 41488 27988 41500
rect 28040 41488 28046 41540
rect 28902 41488 28908 41540
rect 28960 41528 28966 41540
rect 31726 41528 31754 41568
rect 36814 41556 36820 41568
rect 36872 41596 36878 41608
rect 36909 41599 36967 41605
rect 36909 41596 36921 41599
rect 36872 41568 36921 41596
rect 36872 41556 36878 41568
rect 36909 41565 36921 41568
rect 36955 41565 36967 41599
rect 36909 41559 36967 41565
rect 28960 41500 31754 41528
rect 28960 41488 28966 41500
rect 37274 41488 37280 41540
rect 37332 41528 37338 41540
rect 38933 41531 38991 41537
rect 37332 41500 37674 41528
rect 37332 41488 37338 41500
rect 38933 41497 38945 41531
rect 38979 41497 38991 41531
rect 38933 41491 38991 41497
rect 20036 41432 26464 41460
rect 20036 41420 20042 41432
rect 30742 41420 30748 41472
rect 30800 41460 30806 41472
rect 38948 41460 38976 41491
rect 30800 41432 38976 41460
rect 30800 41420 30806 41432
rect 1104 41370 40848 41392
rect 1104 41318 2610 41370
rect 2662 41318 2674 41370
rect 2726 41318 2738 41370
rect 2790 41318 2802 41370
rect 2854 41318 2866 41370
rect 2918 41318 7610 41370
rect 7662 41318 7674 41370
rect 7726 41318 7738 41370
rect 7790 41318 7802 41370
rect 7854 41318 7866 41370
rect 7918 41318 12610 41370
rect 12662 41318 12674 41370
rect 12726 41318 12738 41370
rect 12790 41318 12802 41370
rect 12854 41318 12866 41370
rect 12918 41318 17610 41370
rect 17662 41318 17674 41370
rect 17726 41318 17738 41370
rect 17790 41318 17802 41370
rect 17854 41318 17866 41370
rect 17918 41318 22610 41370
rect 22662 41318 22674 41370
rect 22726 41318 22738 41370
rect 22790 41318 22802 41370
rect 22854 41318 22866 41370
rect 22918 41318 27610 41370
rect 27662 41318 27674 41370
rect 27726 41318 27738 41370
rect 27790 41318 27802 41370
rect 27854 41318 27866 41370
rect 27918 41318 32610 41370
rect 32662 41318 32674 41370
rect 32726 41318 32738 41370
rect 32790 41318 32802 41370
rect 32854 41318 32866 41370
rect 32918 41318 37610 41370
rect 37662 41318 37674 41370
rect 37726 41318 37738 41370
rect 37790 41318 37802 41370
rect 37854 41318 37866 41370
rect 37918 41318 40848 41370
rect 1104 41296 40848 41318
rect 16114 41216 16120 41268
rect 16172 41256 16178 41268
rect 16666 41256 16672 41268
rect 16172 41228 16672 41256
rect 16172 41216 16178 41228
rect 16666 41216 16672 41228
rect 16724 41216 16730 41268
rect 22370 41188 22376 41200
rect 7300 41160 22376 41188
rect 7300 41129 7328 41160
rect 22370 41148 22376 41160
rect 22428 41148 22434 41200
rect 7193 41123 7251 41129
rect 7193 41089 7205 41123
rect 7239 41089 7251 41123
rect 7193 41083 7251 41089
rect 7285 41123 7343 41129
rect 7285 41089 7297 41123
rect 7331 41089 7343 41123
rect 7285 41083 7343 41089
rect 7469 41123 7527 41129
rect 7469 41089 7481 41123
rect 7515 41120 7527 41123
rect 7558 41120 7564 41132
rect 7515 41092 7564 41120
rect 7515 41089 7527 41092
rect 7469 41083 7527 41089
rect 7208 41052 7236 41083
rect 7558 41080 7564 41092
rect 7616 41120 7622 41132
rect 7837 41123 7895 41129
rect 7616 41092 7788 41120
rect 7616 41080 7622 41092
rect 7374 41052 7380 41064
rect 7208 41024 7380 41052
rect 7374 41012 7380 41024
rect 7432 41012 7438 41064
rect 7760 41052 7788 41092
rect 7837 41089 7849 41123
rect 7883 41120 7895 41123
rect 8294 41120 8300 41132
rect 7883 41092 8300 41120
rect 7883 41089 7895 41092
rect 7837 41083 7895 41089
rect 8294 41080 8300 41092
rect 8352 41080 8358 41132
rect 25590 41080 25596 41132
rect 25648 41080 25654 41132
rect 8113 41055 8171 41061
rect 7760 41024 8064 41052
rect 8036 40984 8064 41024
rect 8113 41021 8125 41055
rect 8159 41052 8171 41055
rect 8202 41052 8208 41064
rect 8159 41024 8208 41052
rect 8159 41021 8171 41024
rect 8113 41015 8171 41021
rect 8202 41012 8208 41024
rect 8260 41052 8266 41064
rect 14182 41052 14188 41064
rect 8260 41024 14188 41052
rect 8260 41012 8266 41024
rect 14182 41012 14188 41024
rect 14240 41012 14246 41064
rect 33870 41052 33876 41064
rect 16546 41024 33876 41052
rect 16546 40984 16574 41024
rect 33870 41012 33876 41024
rect 33928 41012 33934 41064
rect 8036 40956 16574 40984
rect 7466 40876 7472 40928
rect 7524 40916 7530 40928
rect 25501 40919 25559 40925
rect 25501 40916 25513 40919
rect 7524 40888 25513 40916
rect 7524 40876 7530 40888
rect 25501 40885 25513 40888
rect 25547 40885 25559 40919
rect 25501 40879 25559 40885
rect 1104 40826 40848 40848
rect 1104 40774 1950 40826
rect 2002 40774 2014 40826
rect 2066 40774 2078 40826
rect 2130 40774 2142 40826
rect 2194 40774 2206 40826
rect 2258 40774 6950 40826
rect 7002 40774 7014 40826
rect 7066 40774 7078 40826
rect 7130 40774 7142 40826
rect 7194 40774 7206 40826
rect 7258 40774 11950 40826
rect 12002 40774 12014 40826
rect 12066 40774 12078 40826
rect 12130 40774 12142 40826
rect 12194 40774 12206 40826
rect 12258 40774 16950 40826
rect 17002 40774 17014 40826
rect 17066 40774 17078 40826
rect 17130 40774 17142 40826
rect 17194 40774 17206 40826
rect 17258 40774 21950 40826
rect 22002 40774 22014 40826
rect 22066 40774 22078 40826
rect 22130 40774 22142 40826
rect 22194 40774 22206 40826
rect 22258 40774 26950 40826
rect 27002 40774 27014 40826
rect 27066 40774 27078 40826
rect 27130 40774 27142 40826
rect 27194 40774 27206 40826
rect 27258 40774 31950 40826
rect 32002 40774 32014 40826
rect 32066 40774 32078 40826
rect 32130 40774 32142 40826
rect 32194 40774 32206 40826
rect 32258 40774 36950 40826
rect 37002 40774 37014 40826
rect 37066 40774 37078 40826
rect 37130 40774 37142 40826
rect 37194 40774 37206 40826
rect 37258 40774 40848 40826
rect 1104 40752 40848 40774
rect 10594 40712 10600 40724
rect 6886 40684 10600 40712
rect 6886 40644 6914 40684
rect 10594 40672 10600 40684
rect 10652 40712 10658 40724
rect 10778 40712 10784 40724
rect 10652 40684 10784 40712
rect 10652 40672 10658 40684
rect 10778 40672 10784 40684
rect 10836 40672 10842 40724
rect 2976 40616 6914 40644
rect 2685 40511 2743 40517
rect 2685 40477 2697 40511
rect 2731 40508 2743 40511
rect 2976 40508 3004 40616
rect 7374 40604 7380 40656
rect 7432 40644 7438 40656
rect 31294 40644 31300 40656
rect 7432 40616 31300 40644
rect 7432 40604 7438 40616
rect 31294 40604 31300 40616
rect 31352 40604 31358 40656
rect 3602 40536 3608 40588
rect 3660 40536 3666 40588
rect 2731 40480 3004 40508
rect 3053 40511 3111 40517
rect 2731 40477 2743 40480
rect 2685 40471 2743 40477
rect 3053 40477 3065 40511
rect 3099 40477 3111 40511
rect 3053 40471 3111 40477
rect 3421 40511 3479 40517
rect 3421 40477 3433 40511
rect 3467 40508 3479 40511
rect 16758 40508 16764 40520
rect 3467 40480 16764 40508
rect 3467 40477 3479 40480
rect 3421 40471 3479 40477
rect 3068 40440 3096 40471
rect 16758 40468 16764 40480
rect 16816 40508 16822 40520
rect 17494 40508 17500 40520
rect 16816 40480 17500 40508
rect 16816 40468 16822 40480
rect 17494 40468 17500 40480
rect 17552 40468 17558 40520
rect 15838 40440 15844 40452
rect 3068 40412 15844 40440
rect 15838 40400 15844 40412
rect 15896 40440 15902 40452
rect 16114 40440 16120 40452
rect 15896 40412 16120 40440
rect 15896 40400 15902 40412
rect 16114 40400 16120 40412
rect 16172 40400 16178 40452
rect 1104 40282 40848 40304
rect 1104 40230 2610 40282
rect 2662 40230 2674 40282
rect 2726 40230 2738 40282
rect 2790 40230 2802 40282
rect 2854 40230 2866 40282
rect 2918 40230 7610 40282
rect 7662 40230 7674 40282
rect 7726 40230 7738 40282
rect 7790 40230 7802 40282
rect 7854 40230 7866 40282
rect 7918 40230 12610 40282
rect 12662 40230 12674 40282
rect 12726 40230 12738 40282
rect 12790 40230 12802 40282
rect 12854 40230 12866 40282
rect 12918 40230 17610 40282
rect 17662 40230 17674 40282
rect 17726 40230 17738 40282
rect 17790 40230 17802 40282
rect 17854 40230 17866 40282
rect 17918 40230 22610 40282
rect 22662 40230 22674 40282
rect 22726 40230 22738 40282
rect 22790 40230 22802 40282
rect 22854 40230 22866 40282
rect 22918 40230 27610 40282
rect 27662 40230 27674 40282
rect 27726 40230 27738 40282
rect 27790 40230 27802 40282
rect 27854 40230 27866 40282
rect 27918 40230 32610 40282
rect 32662 40230 32674 40282
rect 32726 40230 32738 40282
rect 32790 40230 32802 40282
rect 32854 40230 32866 40282
rect 32918 40230 37610 40282
rect 37662 40230 37674 40282
rect 37726 40230 37738 40282
rect 37790 40230 37802 40282
rect 37854 40230 37866 40282
rect 37918 40230 40848 40282
rect 1104 40208 40848 40230
rect 1104 39738 40848 39760
rect 1104 39686 1950 39738
rect 2002 39686 2014 39738
rect 2066 39686 2078 39738
rect 2130 39686 2142 39738
rect 2194 39686 2206 39738
rect 2258 39686 6950 39738
rect 7002 39686 7014 39738
rect 7066 39686 7078 39738
rect 7130 39686 7142 39738
rect 7194 39686 7206 39738
rect 7258 39686 11950 39738
rect 12002 39686 12014 39738
rect 12066 39686 12078 39738
rect 12130 39686 12142 39738
rect 12194 39686 12206 39738
rect 12258 39686 16950 39738
rect 17002 39686 17014 39738
rect 17066 39686 17078 39738
rect 17130 39686 17142 39738
rect 17194 39686 17206 39738
rect 17258 39686 21950 39738
rect 22002 39686 22014 39738
rect 22066 39686 22078 39738
rect 22130 39686 22142 39738
rect 22194 39686 22206 39738
rect 22258 39686 26950 39738
rect 27002 39686 27014 39738
rect 27066 39686 27078 39738
rect 27130 39686 27142 39738
rect 27194 39686 27206 39738
rect 27258 39686 31950 39738
rect 32002 39686 32014 39738
rect 32066 39686 32078 39738
rect 32130 39686 32142 39738
rect 32194 39686 32206 39738
rect 32258 39686 36950 39738
rect 37002 39686 37014 39738
rect 37066 39686 37078 39738
rect 37130 39686 37142 39738
rect 37194 39686 37206 39738
rect 37258 39686 40848 39738
rect 1104 39664 40848 39686
rect 22002 39448 22008 39500
rect 22060 39488 22066 39500
rect 25222 39488 25228 39500
rect 22060 39460 25228 39488
rect 22060 39448 22066 39460
rect 25222 39448 25228 39460
rect 25280 39448 25286 39500
rect 14182 39380 14188 39432
rect 14240 39420 14246 39432
rect 23750 39420 23756 39432
rect 14240 39392 23756 39420
rect 14240 39380 14246 39392
rect 23750 39380 23756 39392
rect 23808 39420 23814 39432
rect 26050 39420 26056 39432
rect 23808 39392 26056 39420
rect 23808 39380 23814 39392
rect 26050 39380 26056 39392
rect 26108 39380 26114 39432
rect 29730 39380 29736 39432
rect 29788 39420 29794 39432
rect 30929 39423 30987 39429
rect 30929 39420 30941 39423
rect 29788 39392 30941 39420
rect 29788 39380 29794 39392
rect 30929 39389 30941 39392
rect 30975 39389 30987 39423
rect 30929 39383 30987 39389
rect 8110 39312 8116 39364
rect 8168 39352 8174 39364
rect 22186 39352 22192 39364
rect 8168 39324 22192 39352
rect 8168 39312 8174 39324
rect 22186 39312 22192 39324
rect 22244 39312 22250 39364
rect 30834 39244 30840 39296
rect 30892 39244 30898 39296
rect 1104 39194 40848 39216
rect 1104 39142 2610 39194
rect 2662 39142 2674 39194
rect 2726 39142 2738 39194
rect 2790 39142 2802 39194
rect 2854 39142 2866 39194
rect 2918 39142 7610 39194
rect 7662 39142 7674 39194
rect 7726 39142 7738 39194
rect 7790 39142 7802 39194
rect 7854 39142 7866 39194
rect 7918 39142 12610 39194
rect 12662 39142 12674 39194
rect 12726 39142 12738 39194
rect 12790 39142 12802 39194
rect 12854 39142 12866 39194
rect 12918 39142 17610 39194
rect 17662 39142 17674 39194
rect 17726 39142 17738 39194
rect 17790 39142 17802 39194
rect 17854 39142 17866 39194
rect 17918 39142 22610 39194
rect 22662 39142 22674 39194
rect 22726 39142 22738 39194
rect 22790 39142 22802 39194
rect 22854 39142 22866 39194
rect 22918 39142 27610 39194
rect 27662 39142 27674 39194
rect 27726 39142 27738 39194
rect 27790 39142 27802 39194
rect 27854 39142 27866 39194
rect 27918 39142 32610 39194
rect 32662 39142 32674 39194
rect 32726 39142 32738 39194
rect 32790 39142 32802 39194
rect 32854 39142 32866 39194
rect 32918 39142 37610 39194
rect 37662 39142 37674 39194
rect 37726 39142 37738 39194
rect 37790 39142 37802 39194
rect 37854 39142 37866 39194
rect 37918 39142 40848 39194
rect 1104 39120 40848 39142
rect 14182 39040 14188 39092
rect 14240 39040 14246 39092
rect 22186 39040 22192 39092
rect 22244 39080 22250 39092
rect 24121 39083 24179 39089
rect 24121 39080 24133 39083
rect 22244 39052 24133 39080
rect 22244 39040 22250 39052
rect 24121 39049 24133 39052
rect 24167 39049 24179 39083
rect 24121 39043 24179 39049
rect 14001 39015 14059 39021
rect 14001 38981 14013 39015
rect 14047 39012 14059 39015
rect 22002 39012 22008 39024
rect 14047 38984 22008 39012
rect 14047 38981 14059 38984
rect 14001 38975 14059 38981
rect 22002 38972 22008 38984
rect 22060 38972 22066 39024
rect 22097 39015 22155 39021
rect 22097 38981 22109 39015
rect 22143 39012 22155 39015
rect 22204 39012 22232 39040
rect 22143 38984 22232 39012
rect 22143 38981 22155 38984
rect 22097 38975 22155 38981
rect 14277 38947 14335 38953
rect 14277 38913 14289 38947
rect 14323 38944 14335 38947
rect 18874 38944 18880 38956
rect 14323 38916 18880 38944
rect 14323 38913 14335 38916
rect 14277 38907 14335 38913
rect 18874 38904 18880 38916
rect 18932 38904 18938 38956
rect 20898 38904 20904 38956
rect 20956 38904 20962 38956
rect 21358 38904 21364 38956
rect 21416 38904 21422 38956
rect 21821 38947 21879 38953
rect 21821 38944 21833 38947
rect 21468 38916 21833 38944
rect 8386 38836 8392 38888
rect 8444 38876 8450 38888
rect 9582 38876 9588 38888
rect 8444 38848 9588 38876
rect 8444 38836 8450 38848
rect 9582 38836 9588 38848
rect 9640 38876 9646 38888
rect 21468 38876 21496 38916
rect 21821 38913 21833 38916
rect 21867 38913 21879 38947
rect 21821 38907 21879 38913
rect 23198 38904 23204 38956
rect 23256 38904 23262 38956
rect 24118 38944 24124 38956
rect 23400 38916 24124 38944
rect 9640 38848 21496 38876
rect 21637 38879 21695 38885
rect 9640 38836 9646 38848
rect 21637 38845 21649 38879
rect 21683 38876 21695 38879
rect 23400 38876 23428 38916
rect 24118 38904 24124 38916
rect 24176 38904 24182 38956
rect 21683 38848 23428 38876
rect 23845 38879 23903 38885
rect 21683 38845 21695 38848
rect 21637 38839 21695 38845
rect 23845 38845 23857 38879
rect 23891 38845 23903 38879
rect 23845 38839 23903 38845
rect 12986 38768 12992 38820
rect 13044 38808 13050 38820
rect 14001 38811 14059 38817
rect 14001 38808 14013 38811
rect 13044 38780 14013 38808
rect 13044 38768 13050 38780
rect 14001 38777 14013 38780
rect 14047 38777 14059 38811
rect 14001 38771 14059 38777
rect 21726 38700 21732 38752
rect 21784 38740 21790 38752
rect 23860 38740 23888 38839
rect 21784 38712 23888 38740
rect 21784 38700 21790 38712
rect 25222 38700 25228 38752
rect 25280 38740 25286 38752
rect 26050 38740 26056 38752
rect 25280 38712 26056 38740
rect 25280 38700 25286 38712
rect 26050 38700 26056 38712
rect 26108 38700 26114 38752
rect 1104 38650 40848 38672
rect 1104 38598 1950 38650
rect 2002 38598 2014 38650
rect 2066 38598 2078 38650
rect 2130 38598 2142 38650
rect 2194 38598 2206 38650
rect 2258 38598 6950 38650
rect 7002 38598 7014 38650
rect 7066 38598 7078 38650
rect 7130 38598 7142 38650
rect 7194 38598 7206 38650
rect 7258 38598 11950 38650
rect 12002 38598 12014 38650
rect 12066 38598 12078 38650
rect 12130 38598 12142 38650
rect 12194 38598 12206 38650
rect 12258 38598 16950 38650
rect 17002 38598 17014 38650
rect 17066 38598 17078 38650
rect 17130 38598 17142 38650
rect 17194 38598 17206 38650
rect 17258 38598 21950 38650
rect 22002 38598 22014 38650
rect 22066 38598 22078 38650
rect 22130 38598 22142 38650
rect 22194 38598 22206 38650
rect 22258 38598 26950 38650
rect 27002 38598 27014 38650
rect 27066 38598 27078 38650
rect 27130 38598 27142 38650
rect 27194 38598 27206 38650
rect 27258 38598 31950 38650
rect 32002 38598 32014 38650
rect 32066 38598 32078 38650
rect 32130 38598 32142 38650
rect 32194 38598 32206 38650
rect 32258 38598 36950 38650
rect 37002 38598 37014 38650
rect 37066 38598 37078 38650
rect 37130 38598 37142 38650
rect 37194 38598 37206 38650
rect 37258 38598 40848 38650
rect 1104 38576 40848 38598
rect 25590 38496 25596 38548
rect 25648 38536 25654 38548
rect 26786 38536 26792 38548
rect 25648 38508 26792 38536
rect 25648 38496 25654 38508
rect 26786 38496 26792 38508
rect 26844 38496 26850 38548
rect 6089 38403 6147 38409
rect 6089 38369 6101 38403
rect 6135 38400 6147 38403
rect 9214 38400 9220 38412
rect 6135 38372 9220 38400
rect 6135 38369 6147 38372
rect 6089 38363 6147 38369
rect 9214 38360 9220 38372
rect 9272 38360 9278 38412
rect 6362 38292 6368 38344
rect 6420 38292 6426 38344
rect 1104 38106 40848 38128
rect 1104 38054 2610 38106
rect 2662 38054 2674 38106
rect 2726 38054 2738 38106
rect 2790 38054 2802 38106
rect 2854 38054 2866 38106
rect 2918 38054 7610 38106
rect 7662 38054 7674 38106
rect 7726 38054 7738 38106
rect 7790 38054 7802 38106
rect 7854 38054 7866 38106
rect 7918 38054 12610 38106
rect 12662 38054 12674 38106
rect 12726 38054 12738 38106
rect 12790 38054 12802 38106
rect 12854 38054 12866 38106
rect 12918 38054 17610 38106
rect 17662 38054 17674 38106
rect 17726 38054 17738 38106
rect 17790 38054 17802 38106
rect 17854 38054 17866 38106
rect 17918 38054 22610 38106
rect 22662 38054 22674 38106
rect 22726 38054 22738 38106
rect 22790 38054 22802 38106
rect 22854 38054 22866 38106
rect 22918 38054 27610 38106
rect 27662 38054 27674 38106
rect 27726 38054 27738 38106
rect 27790 38054 27802 38106
rect 27854 38054 27866 38106
rect 27918 38054 32610 38106
rect 32662 38054 32674 38106
rect 32726 38054 32738 38106
rect 32790 38054 32802 38106
rect 32854 38054 32866 38106
rect 32918 38054 37610 38106
rect 37662 38054 37674 38106
rect 37726 38054 37738 38106
rect 37790 38054 37802 38106
rect 37854 38054 37866 38106
rect 37918 38054 40848 38106
rect 1104 38032 40848 38054
rect 5718 37952 5724 38004
rect 5776 37992 5782 38004
rect 5776 37964 29224 37992
rect 5776 37952 5782 37964
rect 25590 37924 25596 37936
rect 16546 37896 25596 37924
rect 7009 37859 7067 37865
rect 7009 37825 7021 37859
rect 7055 37856 7067 37859
rect 16546 37856 16574 37896
rect 25590 37884 25596 37896
rect 25648 37884 25654 37936
rect 7055 37828 16574 37856
rect 7055 37825 7067 37828
rect 7009 37819 7067 37825
rect 24946 37816 24952 37868
rect 25004 37856 25010 37868
rect 29196 37865 29224 37964
rect 31570 37884 31576 37936
rect 31628 37924 31634 37936
rect 31846 37924 31852 37936
rect 31628 37896 31852 37924
rect 31628 37884 31634 37896
rect 31846 37884 31852 37896
rect 31904 37884 31910 37936
rect 28629 37859 28687 37865
rect 28629 37856 28641 37859
rect 25004 37828 28641 37856
rect 25004 37816 25010 37828
rect 28629 37825 28641 37828
rect 28675 37856 28687 37859
rect 29181 37859 29239 37865
rect 28675 37828 29132 37856
rect 28675 37825 28687 37828
rect 28629 37819 28687 37825
rect 28994 37788 29000 37800
rect 22066 37760 29000 37788
rect 18966 37680 18972 37732
rect 19024 37720 19030 37732
rect 22066 37720 22094 37760
rect 28994 37748 29000 37760
rect 29052 37748 29058 37800
rect 29104 37788 29132 37828
rect 29181 37825 29193 37859
rect 29227 37856 29239 37859
rect 32398 37856 32404 37868
rect 29227 37828 32404 37856
rect 29227 37825 29239 37828
rect 29181 37819 29239 37825
rect 32398 37816 32404 37828
rect 32456 37816 32462 37868
rect 31846 37788 31852 37800
rect 29104 37760 31852 37788
rect 31846 37748 31852 37760
rect 31904 37748 31910 37800
rect 19024 37692 22094 37720
rect 24688 37692 35894 37720
rect 19024 37680 19030 37692
rect 7101 37655 7159 37661
rect 7101 37621 7113 37655
rect 7147 37652 7159 37655
rect 24688 37652 24716 37692
rect 7147 37624 24716 37652
rect 35866 37652 35894 37692
rect 37274 37652 37280 37664
rect 35866 37624 37280 37652
rect 7147 37621 7159 37624
rect 7101 37615 7159 37621
rect 37274 37612 37280 37624
rect 37332 37612 37338 37664
rect 1104 37562 40848 37584
rect 1104 37510 1950 37562
rect 2002 37510 2014 37562
rect 2066 37510 2078 37562
rect 2130 37510 2142 37562
rect 2194 37510 2206 37562
rect 2258 37510 6950 37562
rect 7002 37510 7014 37562
rect 7066 37510 7078 37562
rect 7130 37510 7142 37562
rect 7194 37510 7206 37562
rect 7258 37510 11950 37562
rect 12002 37510 12014 37562
rect 12066 37510 12078 37562
rect 12130 37510 12142 37562
rect 12194 37510 12206 37562
rect 12258 37510 16950 37562
rect 17002 37510 17014 37562
rect 17066 37510 17078 37562
rect 17130 37510 17142 37562
rect 17194 37510 17206 37562
rect 17258 37510 21950 37562
rect 22002 37510 22014 37562
rect 22066 37510 22078 37562
rect 22130 37510 22142 37562
rect 22194 37510 22206 37562
rect 22258 37510 26950 37562
rect 27002 37510 27014 37562
rect 27066 37510 27078 37562
rect 27130 37510 27142 37562
rect 27194 37510 27206 37562
rect 27258 37510 31950 37562
rect 32002 37510 32014 37562
rect 32066 37510 32078 37562
rect 32130 37510 32142 37562
rect 32194 37510 32206 37562
rect 32258 37510 36950 37562
rect 37002 37510 37014 37562
rect 37066 37510 37078 37562
rect 37130 37510 37142 37562
rect 37194 37510 37206 37562
rect 37258 37510 40848 37562
rect 1104 37488 40848 37510
rect 28994 37408 29000 37460
rect 29052 37448 29058 37460
rect 40034 37448 40040 37460
rect 29052 37420 40040 37448
rect 29052 37408 29058 37420
rect 40034 37408 40040 37420
rect 40092 37408 40098 37460
rect 14274 37204 14280 37256
rect 14332 37244 14338 37256
rect 27801 37247 27859 37253
rect 27801 37244 27813 37247
rect 14332 37216 27813 37244
rect 14332 37204 14338 37216
rect 27801 37213 27813 37216
rect 27847 37213 27859 37247
rect 27801 37207 27859 37213
rect 27709 37179 27767 37185
rect 27709 37145 27721 37179
rect 27755 37176 27767 37179
rect 27982 37176 27988 37188
rect 27755 37148 27988 37176
rect 27755 37145 27767 37148
rect 27709 37139 27767 37145
rect 27982 37136 27988 37148
rect 28040 37136 28046 37188
rect 1104 37018 40848 37040
rect 1104 36966 2610 37018
rect 2662 36966 2674 37018
rect 2726 36966 2738 37018
rect 2790 36966 2802 37018
rect 2854 36966 2866 37018
rect 2918 36966 7610 37018
rect 7662 36966 7674 37018
rect 7726 36966 7738 37018
rect 7790 36966 7802 37018
rect 7854 36966 7866 37018
rect 7918 36966 12610 37018
rect 12662 36966 12674 37018
rect 12726 36966 12738 37018
rect 12790 36966 12802 37018
rect 12854 36966 12866 37018
rect 12918 36966 17610 37018
rect 17662 36966 17674 37018
rect 17726 36966 17738 37018
rect 17790 36966 17802 37018
rect 17854 36966 17866 37018
rect 17918 36966 22610 37018
rect 22662 36966 22674 37018
rect 22726 36966 22738 37018
rect 22790 36966 22802 37018
rect 22854 36966 22866 37018
rect 22918 36966 27610 37018
rect 27662 36966 27674 37018
rect 27726 36966 27738 37018
rect 27790 36966 27802 37018
rect 27854 36966 27866 37018
rect 27918 36966 32610 37018
rect 32662 36966 32674 37018
rect 32726 36966 32738 37018
rect 32790 36966 32802 37018
rect 32854 36966 32866 37018
rect 32918 36966 37610 37018
rect 37662 36966 37674 37018
rect 37726 36966 37738 37018
rect 37790 36966 37802 37018
rect 37854 36966 37866 37018
rect 37918 36966 40848 37018
rect 1104 36944 40848 36966
rect 8294 36864 8300 36916
rect 8352 36904 8358 36916
rect 27065 36907 27123 36913
rect 8352 36876 9904 36904
rect 8352 36864 8358 36876
rect 8386 36836 8392 36848
rect 7852 36808 8392 36836
rect 7852 36777 7880 36808
rect 8386 36796 8392 36808
rect 8444 36796 8450 36848
rect 7837 36771 7895 36777
rect 7837 36737 7849 36771
rect 7883 36737 7895 36771
rect 7837 36731 7895 36737
rect 9214 36728 9220 36780
rect 9272 36728 9278 36780
rect 9876 36709 9904 36876
rect 27065 36873 27077 36907
rect 27111 36904 27123 36907
rect 27430 36904 27436 36916
rect 27111 36876 27436 36904
rect 27111 36873 27123 36876
rect 27065 36867 27123 36873
rect 27430 36864 27436 36876
rect 27488 36864 27494 36916
rect 26786 36728 26792 36780
rect 26844 36768 26850 36780
rect 26973 36771 27031 36777
rect 26973 36768 26985 36771
rect 26844 36740 26985 36768
rect 26844 36728 26850 36740
rect 26973 36737 26985 36740
rect 27019 36737 27031 36771
rect 26973 36731 27031 36737
rect 7561 36703 7619 36709
rect 7561 36669 7573 36703
rect 7607 36700 7619 36703
rect 8113 36703 8171 36709
rect 8113 36700 8125 36703
rect 7607 36672 8125 36700
rect 7607 36669 7619 36672
rect 7561 36663 7619 36669
rect 8113 36669 8125 36672
rect 8159 36700 8171 36703
rect 9861 36703 9919 36709
rect 8159 36672 9812 36700
rect 8159 36669 8171 36672
rect 8113 36663 8171 36669
rect 9784 36632 9812 36672
rect 9861 36669 9873 36703
rect 9907 36700 9919 36703
rect 31478 36700 31484 36712
rect 9907 36672 31484 36700
rect 9907 36669 9919 36672
rect 9861 36663 9919 36669
rect 31478 36660 31484 36672
rect 31536 36660 31542 36712
rect 31570 36632 31576 36644
rect 9784 36604 31576 36632
rect 31570 36592 31576 36604
rect 31628 36592 31634 36644
rect 1104 36474 40848 36496
rect 1104 36422 1950 36474
rect 2002 36422 2014 36474
rect 2066 36422 2078 36474
rect 2130 36422 2142 36474
rect 2194 36422 2206 36474
rect 2258 36422 6950 36474
rect 7002 36422 7014 36474
rect 7066 36422 7078 36474
rect 7130 36422 7142 36474
rect 7194 36422 7206 36474
rect 7258 36422 11950 36474
rect 12002 36422 12014 36474
rect 12066 36422 12078 36474
rect 12130 36422 12142 36474
rect 12194 36422 12206 36474
rect 12258 36422 16950 36474
rect 17002 36422 17014 36474
rect 17066 36422 17078 36474
rect 17130 36422 17142 36474
rect 17194 36422 17206 36474
rect 17258 36422 21950 36474
rect 22002 36422 22014 36474
rect 22066 36422 22078 36474
rect 22130 36422 22142 36474
rect 22194 36422 22206 36474
rect 22258 36422 26950 36474
rect 27002 36422 27014 36474
rect 27066 36422 27078 36474
rect 27130 36422 27142 36474
rect 27194 36422 27206 36474
rect 27258 36422 31950 36474
rect 32002 36422 32014 36474
rect 32066 36422 32078 36474
rect 32130 36422 32142 36474
rect 32194 36422 32206 36474
rect 32258 36422 36950 36474
rect 37002 36422 37014 36474
rect 37066 36422 37078 36474
rect 37130 36422 37142 36474
rect 37194 36422 37206 36474
rect 37258 36422 40848 36474
rect 1104 36400 40848 36422
rect 9398 36320 9404 36372
rect 9456 36360 9462 36372
rect 9493 36363 9551 36369
rect 9493 36360 9505 36363
rect 9456 36332 9505 36360
rect 9456 36320 9462 36332
rect 9493 36329 9505 36332
rect 9539 36329 9551 36363
rect 9493 36323 9551 36329
rect 30650 36252 30656 36304
rect 30708 36292 30714 36304
rect 32214 36292 32220 36304
rect 30708 36264 32220 36292
rect 30708 36252 30714 36264
rect 32214 36252 32220 36264
rect 32272 36252 32278 36304
rect 9217 36227 9275 36233
rect 9217 36193 9229 36227
rect 9263 36193 9275 36227
rect 18966 36224 18972 36236
rect 9217 36187 9275 36193
rect 16546 36196 18972 36224
rect 8478 36116 8484 36168
rect 8536 36156 8542 36168
rect 9125 36159 9183 36165
rect 9125 36156 9137 36159
rect 8536 36128 9137 36156
rect 8536 36116 8542 36128
rect 9125 36125 9137 36128
rect 9171 36125 9183 36159
rect 9232 36156 9260 36187
rect 16546 36156 16574 36196
rect 18966 36184 18972 36196
rect 19024 36184 19030 36236
rect 32398 36224 32404 36236
rect 32140 36196 32404 36224
rect 9232 36128 16574 36156
rect 9125 36119 9183 36125
rect 31846 36116 31852 36168
rect 31904 36156 31910 36168
rect 32030 36156 32036 36168
rect 31904 36128 32036 36156
rect 31904 36116 31910 36128
rect 32030 36116 32036 36128
rect 32088 36116 32094 36168
rect 18598 35980 18604 36032
rect 18656 36020 18662 36032
rect 32140 36029 32168 36196
rect 32398 36184 32404 36196
rect 32456 36224 32462 36236
rect 33042 36224 33048 36236
rect 32456 36196 33048 36224
rect 32456 36184 32462 36196
rect 33042 36184 33048 36196
rect 33100 36184 33106 36236
rect 40218 36184 40224 36236
rect 40276 36184 40282 36236
rect 40494 36116 40500 36168
rect 40552 36116 40558 36168
rect 32398 36048 32404 36100
rect 32456 36048 32462 36100
rect 31941 36023 31999 36029
rect 31941 36020 31953 36023
rect 18656 35992 31953 36020
rect 18656 35980 18662 35992
rect 31941 35989 31953 35992
rect 31987 35989 31999 36023
rect 31941 35983 31999 35989
rect 32125 36023 32183 36029
rect 32125 35989 32137 36023
rect 32171 35989 32183 36023
rect 32125 35983 32183 35989
rect 32214 35980 32220 36032
rect 32272 36020 32278 36032
rect 32950 36020 32956 36032
rect 32272 35992 32956 36020
rect 32272 35980 32278 35992
rect 32950 35980 32956 35992
rect 33008 35980 33014 36032
rect 1104 35930 40848 35952
rect 1104 35878 2610 35930
rect 2662 35878 2674 35930
rect 2726 35878 2738 35930
rect 2790 35878 2802 35930
rect 2854 35878 2866 35930
rect 2918 35878 7610 35930
rect 7662 35878 7674 35930
rect 7726 35878 7738 35930
rect 7790 35878 7802 35930
rect 7854 35878 7866 35930
rect 7918 35878 12610 35930
rect 12662 35878 12674 35930
rect 12726 35878 12738 35930
rect 12790 35878 12802 35930
rect 12854 35878 12866 35930
rect 12918 35878 17610 35930
rect 17662 35878 17674 35930
rect 17726 35878 17738 35930
rect 17790 35878 17802 35930
rect 17854 35878 17866 35930
rect 17918 35878 22610 35930
rect 22662 35878 22674 35930
rect 22726 35878 22738 35930
rect 22790 35878 22802 35930
rect 22854 35878 22866 35930
rect 22918 35878 27610 35930
rect 27662 35878 27674 35930
rect 27726 35878 27738 35930
rect 27790 35878 27802 35930
rect 27854 35878 27866 35930
rect 27918 35878 32610 35930
rect 32662 35878 32674 35930
rect 32726 35878 32738 35930
rect 32790 35878 32802 35930
rect 32854 35878 32866 35930
rect 32918 35878 37610 35930
rect 37662 35878 37674 35930
rect 37726 35878 37738 35930
rect 37790 35878 37802 35930
rect 37854 35878 37866 35930
rect 37918 35878 40848 35930
rect 1104 35856 40848 35878
rect 34977 35819 35035 35825
rect 34977 35785 34989 35819
rect 35023 35816 35035 35819
rect 35023 35788 35112 35816
rect 35023 35785 35035 35788
rect 34977 35779 35035 35785
rect 34974 35680 34980 35692
rect 34935 35652 34980 35680
rect 34974 35640 34980 35652
rect 35032 35640 35038 35692
rect 20346 35504 20352 35556
rect 20404 35544 20410 35556
rect 34793 35547 34851 35553
rect 34793 35544 34805 35547
rect 20404 35516 34805 35544
rect 20404 35504 20410 35516
rect 34793 35513 34805 35516
rect 34839 35513 34851 35547
rect 34793 35507 34851 35513
rect 15930 35436 15936 35488
rect 15988 35476 15994 35488
rect 34333 35479 34391 35485
rect 34333 35476 34345 35479
rect 15988 35448 34345 35476
rect 15988 35436 15994 35448
rect 34333 35445 34345 35448
rect 34379 35476 34391 35479
rect 35084 35476 35112 35788
rect 35434 35572 35440 35624
rect 35492 35572 35498 35624
rect 34379 35448 35112 35476
rect 34379 35445 34391 35448
rect 34333 35439 34391 35445
rect 35342 35436 35348 35488
rect 35400 35476 35406 35488
rect 39022 35476 39028 35488
rect 35400 35448 39028 35476
rect 35400 35436 35406 35448
rect 39022 35436 39028 35448
rect 39080 35436 39086 35488
rect 1104 35386 40848 35408
rect 1104 35334 1950 35386
rect 2002 35334 2014 35386
rect 2066 35334 2078 35386
rect 2130 35334 2142 35386
rect 2194 35334 2206 35386
rect 2258 35334 6950 35386
rect 7002 35334 7014 35386
rect 7066 35334 7078 35386
rect 7130 35334 7142 35386
rect 7194 35334 7206 35386
rect 7258 35334 11950 35386
rect 12002 35334 12014 35386
rect 12066 35334 12078 35386
rect 12130 35334 12142 35386
rect 12194 35334 12206 35386
rect 12258 35334 16950 35386
rect 17002 35334 17014 35386
rect 17066 35334 17078 35386
rect 17130 35334 17142 35386
rect 17194 35334 17206 35386
rect 17258 35334 21950 35386
rect 22002 35334 22014 35386
rect 22066 35334 22078 35386
rect 22130 35334 22142 35386
rect 22194 35334 22206 35386
rect 22258 35334 26950 35386
rect 27002 35334 27014 35386
rect 27066 35334 27078 35386
rect 27130 35334 27142 35386
rect 27194 35334 27206 35386
rect 27258 35334 31950 35386
rect 32002 35334 32014 35386
rect 32066 35334 32078 35386
rect 32130 35334 32142 35386
rect 32194 35334 32206 35386
rect 32258 35334 36950 35386
rect 37002 35334 37014 35386
rect 37066 35334 37078 35386
rect 37130 35334 37142 35386
rect 37194 35334 37206 35386
rect 37258 35334 40848 35386
rect 1104 35312 40848 35334
rect 29822 35164 29828 35216
rect 29880 35204 29886 35216
rect 36722 35204 36728 35216
rect 29880 35176 36728 35204
rect 29880 35164 29886 35176
rect 36722 35164 36728 35176
rect 36780 35164 36786 35216
rect 1104 34842 40848 34864
rect 1104 34790 2610 34842
rect 2662 34790 2674 34842
rect 2726 34790 2738 34842
rect 2790 34790 2802 34842
rect 2854 34790 2866 34842
rect 2918 34790 7610 34842
rect 7662 34790 7674 34842
rect 7726 34790 7738 34842
rect 7790 34790 7802 34842
rect 7854 34790 7866 34842
rect 7918 34790 12610 34842
rect 12662 34790 12674 34842
rect 12726 34790 12738 34842
rect 12790 34790 12802 34842
rect 12854 34790 12866 34842
rect 12918 34790 17610 34842
rect 17662 34790 17674 34842
rect 17726 34790 17738 34842
rect 17790 34790 17802 34842
rect 17854 34790 17866 34842
rect 17918 34790 22610 34842
rect 22662 34790 22674 34842
rect 22726 34790 22738 34842
rect 22790 34790 22802 34842
rect 22854 34790 22866 34842
rect 22918 34790 27610 34842
rect 27662 34790 27674 34842
rect 27726 34790 27738 34842
rect 27790 34790 27802 34842
rect 27854 34790 27866 34842
rect 27918 34790 32610 34842
rect 32662 34790 32674 34842
rect 32726 34790 32738 34842
rect 32790 34790 32802 34842
rect 32854 34790 32866 34842
rect 32918 34790 37610 34842
rect 37662 34790 37674 34842
rect 37726 34790 37738 34842
rect 37790 34790 37802 34842
rect 37854 34790 37866 34842
rect 37918 34790 40848 34842
rect 1104 34768 40848 34790
rect 17402 34620 17408 34672
rect 17460 34660 17466 34672
rect 17460 34632 22094 34660
rect 17460 34620 17466 34632
rect 15470 34552 15476 34604
rect 15528 34592 15534 34604
rect 15930 34592 15936 34604
rect 15528 34564 15936 34592
rect 15528 34552 15534 34564
rect 15930 34552 15936 34564
rect 15988 34552 15994 34604
rect 22066 34592 22094 34632
rect 32677 34595 32735 34601
rect 32677 34592 32689 34595
rect 22066 34564 32689 34592
rect 32677 34561 32689 34564
rect 32723 34561 32735 34595
rect 32677 34555 32735 34561
rect 32953 34595 33011 34601
rect 32953 34561 32965 34595
rect 32999 34592 33011 34595
rect 35434 34592 35440 34604
rect 32999 34564 35440 34592
rect 32999 34561 33011 34564
rect 32953 34555 33011 34561
rect 35434 34552 35440 34564
rect 35492 34552 35498 34604
rect 8662 34484 8668 34536
rect 8720 34524 8726 34536
rect 32585 34527 32643 34533
rect 32585 34524 32597 34527
rect 8720 34496 32597 34524
rect 8720 34484 8726 34496
rect 32585 34493 32597 34496
rect 32631 34493 32643 34527
rect 32585 34487 32643 34493
rect 1104 34298 40848 34320
rect 1104 34246 1950 34298
rect 2002 34246 2014 34298
rect 2066 34246 2078 34298
rect 2130 34246 2142 34298
rect 2194 34246 2206 34298
rect 2258 34246 6950 34298
rect 7002 34246 7014 34298
rect 7066 34246 7078 34298
rect 7130 34246 7142 34298
rect 7194 34246 7206 34298
rect 7258 34246 11950 34298
rect 12002 34246 12014 34298
rect 12066 34246 12078 34298
rect 12130 34246 12142 34298
rect 12194 34246 12206 34298
rect 12258 34246 16950 34298
rect 17002 34246 17014 34298
rect 17066 34246 17078 34298
rect 17130 34246 17142 34298
rect 17194 34246 17206 34298
rect 17258 34246 21950 34298
rect 22002 34246 22014 34298
rect 22066 34246 22078 34298
rect 22130 34246 22142 34298
rect 22194 34246 22206 34298
rect 22258 34246 26950 34298
rect 27002 34246 27014 34298
rect 27066 34246 27078 34298
rect 27130 34246 27142 34298
rect 27194 34246 27206 34298
rect 27258 34246 31950 34298
rect 32002 34246 32014 34298
rect 32066 34246 32078 34298
rect 32130 34246 32142 34298
rect 32194 34246 32206 34298
rect 32258 34246 36950 34298
rect 37002 34246 37014 34298
rect 37066 34246 37078 34298
rect 37130 34246 37142 34298
rect 37194 34246 37206 34298
rect 37258 34246 40848 34298
rect 1104 34224 40848 34246
rect 18874 34144 18880 34196
rect 18932 34184 18938 34196
rect 25130 34184 25136 34196
rect 18932 34156 25136 34184
rect 18932 34144 18938 34156
rect 25130 34144 25136 34156
rect 25188 34144 25194 34196
rect 10686 34076 10692 34128
rect 10744 34116 10750 34128
rect 10744 34088 20576 34116
rect 10744 34076 10750 34088
rect 19610 33940 19616 33992
rect 19668 33940 19674 33992
rect 20548 33980 20576 34088
rect 23290 34008 23296 34060
rect 23348 34048 23354 34060
rect 23348 34020 24716 34048
rect 23348 34008 23354 34020
rect 24688 33989 24716 34020
rect 25130 34008 25136 34060
rect 25188 34008 25194 34060
rect 24397 33983 24455 33989
rect 24397 33980 24409 33983
rect 20548 33952 24409 33980
rect 24397 33949 24409 33952
rect 24443 33949 24455 33983
rect 24397 33943 24455 33949
rect 24673 33983 24731 33989
rect 24673 33949 24685 33983
rect 24719 33949 24731 33983
rect 24673 33943 24731 33949
rect 14826 33872 14832 33924
rect 14884 33912 14890 33924
rect 15102 33912 15108 33924
rect 14884 33884 15108 33912
rect 14884 33872 14890 33884
rect 15102 33872 15108 33884
rect 15160 33912 15166 33924
rect 24765 33915 24823 33921
rect 24765 33912 24777 33915
rect 15160 33884 22094 33912
rect 15160 33872 15166 33884
rect 21082 33804 21088 33856
rect 21140 33804 21146 33856
rect 22066 33844 22094 33884
rect 24504 33884 24777 33912
rect 24504 33844 24532 33884
rect 24765 33881 24777 33884
rect 24811 33881 24823 33915
rect 24765 33875 24823 33881
rect 22066 33816 24532 33844
rect 24578 33804 24584 33856
rect 24636 33804 24642 33856
rect 1104 33754 40848 33776
rect 1104 33702 2610 33754
rect 2662 33702 2674 33754
rect 2726 33702 2738 33754
rect 2790 33702 2802 33754
rect 2854 33702 2866 33754
rect 2918 33702 7610 33754
rect 7662 33702 7674 33754
rect 7726 33702 7738 33754
rect 7790 33702 7802 33754
rect 7854 33702 7866 33754
rect 7918 33702 12610 33754
rect 12662 33702 12674 33754
rect 12726 33702 12738 33754
rect 12790 33702 12802 33754
rect 12854 33702 12866 33754
rect 12918 33702 17610 33754
rect 17662 33702 17674 33754
rect 17726 33702 17738 33754
rect 17790 33702 17802 33754
rect 17854 33702 17866 33754
rect 17918 33702 22610 33754
rect 22662 33702 22674 33754
rect 22726 33702 22738 33754
rect 22790 33702 22802 33754
rect 22854 33702 22866 33754
rect 22918 33702 27610 33754
rect 27662 33702 27674 33754
rect 27726 33702 27738 33754
rect 27790 33702 27802 33754
rect 27854 33702 27866 33754
rect 27918 33702 32610 33754
rect 32662 33702 32674 33754
rect 32726 33702 32738 33754
rect 32790 33702 32802 33754
rect 32854 33702 32866 33754
rect 32918 33702 37610 33754
rect 37662 33702 37674 33754
rect 37726 33702 37738 33754
rect 37790 33702 37802 33754
rect 37854 33702 37866 33754
rect 37918 33702 40848 33754
rect 1104 33680 40848 33702
rect 9214 33600 9220 33652
rect 9272 33640 9278 33652
rect 10413 33643 10471 33649
rect 10413 33640 10425 33643
rect 9272 33612 10425 33640
rect 9272 33600 9278 33612
rect 10413 33609 10425 33612
rect 10459 33609 10471 33643
rect 10413 33603 10471 33609
rect 10502 33600 10508 33652
rect 10560 33640 10566 33652
rect 14366 33640 14372 33652
rect 10560 33612 14372 33640
rect 10560 33600 10566 33612
rect 14366 33600 14372 33612
rect 14424 33640 14430 33652
rect 24578 33640 24584 33652
rect 14424 33612 24584 33640
rect 14424 33600 14430 33612
rect 24578 33600 24584 33612
rect 24636 33600 24642 33652
rect 10505 33507 10563 33513
rect 10505 33473 10517 33507
rect 10551 33504 10563 33507
rect 14918 33504 14924 33516
rect 10551 33476 14924 33504
rect 10551 33473 10563 33476
rect 10505 33467 10563 33473
rect 14918 33464 14924 33476
rect 14976 33464 14982 33516
rect 31754 33464 31760 33516
rect 31812 33504 31818 33516
rect 33045 33507 33103 33513
rect 33045 33504 33057 33507
rect 31812 33476 33057 33504
rect 31812 33464 31818 33476
rect 33045 33473 33057 33476
rect 33091 33473 33103 33507
rect 33045 33467 33103 33473
rect 10410 33260 10416 33312
rect 10468 33300 10474 33312
rect 10686 33300 10692 33312
rect 10468 33272 10692 33300
rect 10468 33260 10474 33272
rect 10686 33260 10692 33272
rect 10744 33260 10750 33312
rect 18598 33260 18604 33312
rect 18656 33300 18662 33312
rect 18874 33300 18880 33312
rect 18656 33272 18880 33300
rect 18656 33260 18662 33272
rect 18874 33260 18880 33272
rect 18932 33260 18938 33312
rect 24670 33260 24676 33312
rect 24728 33300 24734 33312
rect 32861 33303 32919 33309
rect 32861 33300 32873 33303
rect 24728 33272 32873 33300
rect 24728 33260 24734 33272
rect 32861 33269 32873 33272
rect 32907 33269 32919 33303
rect 32861 33263 32919 33269
rect 1104 33210 40848 33232
rect 1104 33158 1950 33210
rect 2002 33158 2014 33210
rect 2066 33158 2078 33210
rect 2130 33158 2142 33210
rect 2194 33158 2206 33210
rect 2258 33158 6950 33210
rect 7002 33158 7014 33210
rect 7066 33158 7078 33210
rect 7130 33158 7142 33210
rect 7194 33158 7206 33210
rect 7258 33158 11950 33210
rect 12002 33158 12014 33210
rect 12066 33158 12078 33210
rect 12130 33158 12142 33210
rect 12194 33158 12206 33210
rect 12258 33158 16950 33210
rect 17002 33158 17014 33210
rect 17066 33158 17078 33210
rect 17130 33158 17142 33210
rect 17194 33158 17206 33210
rect 17258 33158 21950 33210
rect 22002 33158 22014 33210
rect 22066 33158 22078 33210
rect 22130 33158 22142 33210
rect 22194 33158 22206 33210
rect 22258 33158 26950 33210
rect 27002 33158 27014 33210
rect 27066 33158 27078 33210
rect 27130 33158 27142 33210
rect 27194 33158 27206 33210
rect 27258 33158 31950 33210
rect 32002 33158 32014 33210
rect 32066 33158 32078 33210
rect 32130 33158 32142 33210
rect 32194 33158 32206 33210
rect 32258 33158 36950 33210
rect 37002 33158 37014 33210
rect 37066 33158 37078 33210
rect 37130 33158 37142 33210
rect 37194 33158 37206 33210
rect 37258 33158 40848 33210
rect 1104 33136 40848 33158
rect 15378 32716 15384 32768
rect 15436 32756 15442 32768
rect 16482 32756 16488 32768
rect 15436 32728 16488 32756
rect 15436 32716 15442 32728
rect 16482 32716 16488 32728
rect 16540 32756 16546 32768
rect 31478 32756 31484 32768
rect 16540 32728 31484 32756
rect 16540 32716 16546 32728
rect 31478 32716 31484 32728
rect 31536 32716 31542 32768
rect 38102 32716 38108 32768
rect 38160 32756 38166 32768
rect 38562 32756 38568 32768
rect 38160 32728 38568 32756
rect 38160 32716 38166 32728
rect 38562 32716 38568 32728
rect 38620 32716 38626 32768
rect 1104 32666 40848 32688
rect 1104 32614 2610 32666
rect 2662 32614 2674 32666
rect 2726 32614 2738 32666
rect 2790 32614 2802 32666
rect 2854 32614 2866 32666
rect 2918 32614 7610 32666
rect 7662 32614 7674 32666
rect 7726 32614 7738 32666
rect 7790 32614 7802 32666
rect 7854 32614 7866 32666
rect 7918 32614 12610 32666
rect 12662 32614 12674 32666
rect 12726 32614 12738 32666
rect 12790 32614 12802 32666
rect 12854 32614 12866 32666
rect 12918 32614 17610 32666
rect 17662 32614 17674 32666
rect 17726 32614 17738 32666
rect 17790 32614 17802 32666
rect 17854 32614 17866 32666
rect 17918 32614 22610 32666
rect 22662 32614 22674 32666
rect 22726 32614 22738 32666
rect 22790 32614 22802 32666
rect 22854 32614 22866 32666
rect 22918 32614 27610 32666
rect 27662 32614 27674 32666
rect 27726 32614 27738 32666
rect 27790 32614 27802 32666
rect 27854 32614 27866 32666
rect 27918 32614 32610 32666
rect 32662 32614 32674 32666
rect 32726 32614 32738 32666
rect 32790 32614 32802 32666
rect 32854 32614 32866 32666
rect 32918 32614 37610 32666
rect 37662 32614 37674 32666
rect 37726 32614 37738 32666
rect 37790 32614 37802 32666
rect 37854 32614 37866 32666
rect 37918 32614 40848 32666
rect 1104 32592 40848 32614
rect 6362 32512 6368 32564
rect 6420 32552 6426 32564
rect 40126 32552 40132 32564
rect 6420 32524 40132 32552
rect 6420 32512 6426 32524
rect 40126 32512 40132 32524
rect 40184 32512 40190 32564
rect 13078 32444 13084 32496
rect 13136 32484 13142 32496
rect 13136 32456 22094 32484
rect 13136 32444 13142 32456
rect 6822 32376 6828 32428
rect 6880 32416 6886 32428
rect 18509 32419 18567 32425
rect 18509 32416 18521 32419
rect 6880 32388 18521 32416
rect 6880 32376 6886 32388
rect 18509 32385 18521 32388
rect 18555 32385 18567 32419
rect 22066 32416 22094 32456
rect 28258 32444 28264 32496
rect 28316 32484 28322 32496
rect 31389 32487 31447 32493
rect 31389 32484 31401 32487
rect 28316 32456 31401 32484
rect 28316 32444 28322 32456
rect 31389 32453 31401 32456
rect 31435 32453 31447 32487
rect 31389 32447 31447 32453
rect 28902 32416 28908 32428
rect 22066 32388 28908 32416
rect 18509 32379 18567 32385
rect 28902 32376 28908 32388
rect 28960 32376 28966 32428
rect 31478 32376 31484 32428
rect 31536 32376 31542 32428
rect 36814 32376 36820 32428
rect 36872 32416 36878 32428
rect 37277 32419 37335 32425
rect 37277 32416 37289 32419
rect 36872 32388 37289 32416
rect 36872 32376 36878 32388
rect 37277 32385 37289 32388
rect 37323 32385 37335 32419
rect 37277 32379 37335 32385
rect 38654 32376 38660 32428
rect 38712 32376 38718 32428
rect 18046 32308 18052 32360
rect 18104 32308 18110 32360
rect 18601 32351 18659 32357
rect 18601 32317 18613 32351
rect 18647 32348 18659 32351
rect 19150 32348 19156 32360
rect 18647 32320 19156 32348
rect 18647 32317 18659 32320
rect 18601 32311 18659 32317
rect 19150 32308 19156 32320
rect 19208 32308 19214 32360
rect 28920 32348 28948 32376
rect 35434 32348 35440 32360
rect 28920 32320 35440 32348
rect 35434 32308 35440 32320
rect 35492 32308 35498 32360
rect 37553 32351 37611 32357
rect 37553 32317 37565 32351
rect 37599 32348 37611 32351
rect 38286 32348 38292 32360
rect 37599 32320 38292 32348
rect 37599 32317 37611 32320
rect 37553 32311 37611 32317
rect 38286 32308 38292 32320
rect 38344 32308 38350 32360
rect 38562 32308 38568 32360
rect 38620 32348 38626 32360
rect 39301 32351 39359 32357
rect 39301 32348 39313 32351
rect 38620 32320 39313 32348
rect 38620 32308 38626 32320
rect 39301 32317 39313 32320
rect 39347 32317 39359 32351
rect 39301 32311 39359 32317
rect 25222 32240 25228 32292
rect 25280 32280 25286 32292
rect 25280 32252 31754 32280
rect 25280 32240 25286 32252
rect 31726 32212 31754 32252
rect 35342 32212 35348 32224
rect 31726 32184 35348 32212
rect 35342 32172 35348 32184
rect 35400 32172 35406 32224
rect 1104 32122 40848 32144
rect 1104 32070 1950 32122
rect 2002 32070 2014 32122
rect 2066 32070 2078 32122
rect 2130 32070 2142 32122
rect 2194 32070 2206 32122
rect 2258 32070 6950 32122
rect 7002 32070 7014 32122
rect 7066 32070 7078 32122
rect 7130 32070 7142 32122
rect 7194 32070 7206 32122
rect 7258 32070 11950 32122
rect 12002 32070 12014 32122
rect 12066 32070 12078 32122
rect 12130 32070 12142 32122
rect 12194 32070 12206 32122
rect 12258 32070 16950 32122
rect 17002 32070 17014 32122
rect 17066 32070 17078 32122
rect 17130 32070 17142 32122
rect 17194 32070 17206 32122
rect 17258 32070 21950 32122
rect 22002 32070 22014 32122
rect 22066 32070 22078 32122
rect 22130 32070 22142 32122
rect 22194 32070 22206 32122
rect 22258 32070 26950 32122
rect 27002 32070 27014 32122
rect 27066 32070 27078 32122
rect 27130 32070 27142 32122
rect 27194 32070 27206 32122
rect 27258 32070 31950 32122
rect 32002 32070 32014 32122
rect 32066 32070 32078 32122
rect 32130 32070 32142 32122
rect 32194 32070 32206 32122
rect 32258 32070 36950 32122
rect 37002 32070 37014 32122
rect 37066 32070 37078 32122
rect 37130 32070 37142 32122
rect 37194 32070 37206 32122
rect 37258 32070 40848 32122
rect 1104 32048 40848 32070
rect 24210 31968 24216 32020
rect 24268 32008 24274 32020
rect 29641 32011 29699 32017
rect 29641 32008 29653 32011
rect 24268 31980 29653 32008
rect 24268 31968 24274 31980
rect 29641 31977 29653 31980
rect 29687 31977 29699 32011
rect 29641 31971 29699 31977
rect 39482 31968 39488 32020
rect 39540 32008 39546 32020
rect 39666 32008 39672 32020
rect 39540 31980 39672 32008
rect 39540 31968 39546 31980
rect 39666 31968 39672 31980
rect 39724 32008 39730 32020
rect 39853 32011 39911 32017
rect 39853 32008 39865 32011
rect 39724 31980 39865 32008
rect 39724 31968 39730 31980
rect 39853 31977 39865 31980
rect 39899 31977 39911 32011
rect 39853 31971 39911 31977
rect 40126 31968 40132 32020
rect 40184 32008 40190 32020
rect 40221 32011 40279 32017
rect 40221 32008 40233 32011
rect 40184 31980 40233 32008
rect 40184 31968 40190 31980
rect 40221 31977 40233 31980
rect 40267 31977 40279 32011
rect 40221 31971 40279 31977
rect 6178 31900 6184 31952
rect 6236 31940 6242 31952
rect 28718 31940 28724 31952
rect 6236 31912 28724 31940
rect 6236 31900 6242 31912
rect 28718 31900 28724 31912
rect 28776 31940 28782 31952
rect 28776 31912 36216 31940
rect 28776 31900 28782 31912
rect 25406 31832 25412 31884
rect 25464 31832 25470 31884
rect 35434 31832 35440 31884
rect 35492 31872 35498 31884
rect 35492 31844 36124 31872
rect 35492 31832 35498 31844
rect 20898 31764 20904 31816
rect 20956 31804 20962 31816
rect 21358 31804 21364 31816
rect 20956 31776 21364 31804
rect 20956 31764 20962 31776
rect 21358 31764 21364 31776
rect 21416 31804 21422 31816
rect 25222 31804 25228 31816
rect 21416 31776 25228 31804
rect 21416 31764 21422 31776
rect 25222 31764 25228 31776
rect 25280 31764 25286 31816
rect 25777 31807 25835 31813
rect 25777 31773 25789 31807
rect 25823 31804 25835 31807
rect 29733 31807 29791 31813
rect 25823 31776 29592 31804
rect 25823 31773 25835 31776
rect 25777 31767 25835 31773
rect 29564 31754 29592 31776
rect 29733 31773 29745 31807
rect 29779 31804 29791 31807
rect 29822 31804 29828 31816
rect 29779 31776 29828 31804
rect 29779 31773 29791 31776
rect 29733 31767 29791 31773
rect 29822 31764 29828 31776
rect 29880 31764 29886 31816
rect 34882 31804 34888 31816
rect 29932 31776 34888 31804
rect 7374 31696 7380 31748
rect 7432 31736 7438 31748
rect 29454 31736 29460 31748
rect 7432 31708 29460 31736
rect 7432 31696 7438 31708
rect 29454 31696 29460 31708
rect 29512 31696 29518 31748
rect 29564 31726 29684 31754
rect 29656 31668 29684 31726
rect 29932 31668 29960 31776
rect 34882 31764 34888 31776
rect 34940 31764 34946 31816
rect 36096 31736 36124 31844
rect 36188 31813 36216 31912
rect 36446 31832 36452 31884
rect 36504 31872 36510 31884
rect 39393 31875 39451 31881
rect 39393 31872 39405 31875
rect 36504 31844 39405 31872
rect 36504 31832 36510 31844
rect 39393 31841 39405 31844
rect 39439 31872 39451 31875
rect 39945 31875 40003 31881
rect 39945 31872 39957 31875
rect 39439 31844 39957 31872
rect 39439 31841 39451 31844
rect 39393 31835 39451 31841
rect 39945 31841 39957 31844
rect 39991 31841 40003 31875
rect 39945 31835 40003 31841
rect 36173 31807 36231 31813
rect 36173 31773 36185 31807
rect 36219 31773 36231 31807
rect 36173 31767 36231 31773
rect 36538 31764 36544 31816
rect 36596 31764 36602 31816
rect 36633 31807 36691 31813
rect 36633 31773 36645 31807
rect 36679 31773 36691 31807
rect 36633 31767 36691 31773
rect 36648 31736 36676 31767
rect 39758 31764 39764 31816
rect 39816 31804 39822 31816
rect 39853 31807 39911 31813
rect 39853 31804 39865 31807
rect 39816 31776 39865 31804
rect 39816 31764 39822 31776
rect 39853 31773 39865 31776
rect 39899 31773 39911 31807
rect 39853 31767 39911 31773
rect 36096 31708 36676 31736
rect 29656 31640 29960 31668
rect 1104 31578 40848 31600
rect 1104 31526 2610 31578
rect 2662 31526 2674 31578
rect 2726 31526 2738 31578
rect 2790 31526 2802 31578
rect 2854 31526 2866 31578
rect 2918 31526 7610 31578
rect 7662 31526 7674 31578
rect 7726 31526 7738 31578
rect 7790 31526 7802 31578
rect 7854 31526 7866 31578
rect 7918 31526 12610 31578
rect 12662 31526 12674 31578
rect 12726 31526 12738 31578
rect 12790 31526 12802 31578
rect 12854 31526 12866 31578
rect 12918 31526 17610 31578
rect 17662 31526 17674 31578
rect 17726 31526 17738 31578
rect 17790 31526 17802 31578
rect 17854 31526 17866 31578
rect 17918 31526 22610 31578
rect 22662 31526 22674 31578
rect 22726 31526 22738 31578
rect 22790 31526 22802 31578
rect 22854 31526 22866 31578
rect 22918 31526 27610 31578
rect 27662 31526 27674 31578
rect 27726 31526 27738 31578
rect 27790 31526 27802 31578
rect 27854 31526 27866 31578
rect 27918 31526 32610 31578
rect 32662 31526 32674 31578
rect 32726 31526 32738 31578
rect 32790 31526 32802 31578
rect 32854 31526 32866 31578
rect 32918 31526 37610 31578
rect 37662 31526 37674 31578
rect 37726 31526 37738 31578
rect 37790 31526 37802 31578
rect 37854 31526 37866 31578
rect 37918 31526 40848 31578
rect 1104 31504 40848 31526
rect 7561 31467 7619 31473
rect 7561 31433 7573 31467
rect 7607 31464 7619 31467
rect 14642 31464 14648 31476
rect 7607 31436 14648 31464
rect 7607 31433 7619 31436
rect 7561 31427 7619 31433
rect 14642 31424 14648 31436
rect 14700 31424 14706 31476
rect 17402 31424 17408 31476
rect 17460 31464 17466 31476
rect 17460 31436 26234 31464
rect 17460 31424 17466 31436
rect 19610 31356 19616 31408
rect 19668 31356 19674 31408
rect 7374 31288 7380 31340
rect 7432 31288 7438 31340
rect 7653 31331 7711 31337
rect 7653 31297 7665 31331
rect 7699 31328 7711 31331
rect 8202 31328 8208 31340
rect 7699 31300 8208 31328
rect 7699 31297 7711 31300
rect 7653 31291 7711 31297
rect 8202 31288 8208 31300
rect 8260 31288 8266 31340
rect 18138 31220 18144 31272
rect 18196 31260 18202 31272
rect 18877 31263 18935 31269
rect 18877 31260 18889 31263
rect 18196 31232 18889 31260
rect 18196 31220 18202 31232
rect 18877 31229 18889 31232
rect 18923 31229 18935 31263
rect 19153 31263 19211 31269
rect 19153 31260 19165 31263
rect 18877 31223 18935 31229
rect 18984 31232 19165 31260
rect 2406 31152 2412 31204
rect 2464 31192 2470 31204
rect 18509 31195 18567 31201
rect 18509 31192 18521 31195
rect 2464 31164 18521 31192
rect 2464 31152 2470 31164
rect 18509 31161 18521 31164
rect 18555 31192 18567 31195
rect 18984 31192 19012 31232
rect 19153 31229 19165 31232
rect 19199 31229 19211 31263
rect 19153 31223 19211 31229
rect 20898 31220 20904 31272
rect 20956 31220 20962 31272
rect 18555 31164 19012 31192
rect 26206 31192 26234 31436
rect 31570 31424 31576 31476
rect 31628 31464 31634 31476
rect 33137 31467 33195 31473
rect 33137 31464 33149 31467
rect 31628 31436 33149 31464
rect 31628 31424 31634 31436
rect 33137 31433 33149 31436
rect 33183 31433 33195 31467
rect 33137 31427 33195 31433
rect 33152 31328 33180 31427
rect 33594 31356 33600 31408
rect 33652 31396 33658 31408
rect 33652 31368 33824 31396
rect 33652 31356 33658 31368
rect 33796 31337 33824 31368
rect 33505 31331 33563 31337
rect 33505 31328 33517 31331
rect 33152 31300 33517 31328
rect 33505 31297 33517 31300
rect 33551 31297 33563 31331
rect 33505 31291 33563 31297
rect 33689 31331 33747 31337
rect 33689 31297 33701 31331
rect 33735 31297 33747 31331
rect 33689 31291 33747 31297
rect 33781 31331 33839 31337
rect 33781 31297 33793 31331
rect 33827 31297 33839 31331
rect 33781 31291 33839 31297
rect 31846 31220 31852 31272
rect 31904 31260 31910 31272
rect 33704 31260 33732 31291
rect 31904 31232 33732 31260
rect 31904 31220 31910 31232
rect 33226 31192 33232 31204
rect 26206 31164 33232 31192
rect 18555 31161 18567 31164
rect 18509 31155 18567 31161
rect 33226 31152 33232 31164
rect 33284 31152 33290 31204
rect 7193 31127 7251 31133
rect 7193 31093 7205 31127
rect 7239 31124 7251 31127
rect 16574 31124 16580 31136
rect 7239 31096 16580 31124
rect 7239 31093 7251 31096
rect 7193 31087 7251 31093
rect 16574 31084 16580 31096
rect 16632 31084 16638 31136
rect 29454 31084 29460 31136
rect 29512 31124 29518 31136
rect 33502 31124 33508 31136
rect 29512 31096 33508 31124
rect 29512 31084 29518 31096
rect 33502 31084 33508 31096
rect 33560 31124 33566 31136
rect 33965 31127 34023 31133
rect 33965 31124 33977 31127
rect 33560 31096 33977 31124
rect 33560 31084 33566 31096
rect 33965 31093 33977 31096
rect 34011 31093 34023 31127
rect 33965 31087 34023 31093
rect 1104 31034 40848 31056
rect 1104 30982 1950 31034
rect 2002 30982 2014 31034
rect 2066 30982 2078 31034
rect 2130 30982 2142 31034
rect 2194 30982 2206 31034
rect 2258 30982 6950 31034
rect 7002 30982 7014 31034
rect 7066 30982 7078 31034
rect 7130 30982 7142 31034
rect 7194 30982 7206 31034
rect 7258 30982 11950 31034
rect 12002 30982 12014 31034
rect 12066 30982 12078 31034
rect 12130 30982 12142 31034
rect 12194 30982 12206 31034
rect 12258 30982 16950 31034
rect 17002 30982 17014 31034
rect 17066 30982 17078 31034
rect 17130 30982 17142 31034
rect 17194 30982 17206 31034
rect 17258 30982 21950 31034
rect 22002 30982 22014 31034
rect 22066 30982 22078 31034
rect 22130 30982 22142 31034
rect 22194 30982 22206 31034
rect 22258 30982 26950 31034
rect 27002 30982 27014 31034
rect 27066 30982 27078 31034
rect 27130 30982 27142 31034
rect 27194 30982 27206 31034
rect 27258 30982 31950 31034
rect 32002 30982 32014 31034
rect 32066 30982 32078 31034
rect 32130 30982 32142 31034
rect 32194 30982 32206 31034
rect 32258 30982 36950 31034
rect 37002 30982 37014 31034
rect 37066 30982 37078 31034
rect 37130 30982 37142 31034
rect 37194 30982 37206 31034
rect 37258 30982 40848 31034
rect 1104 30960 40848 30982
rect 9232 30892 12434 30920
rect 9030 30812 9036 30864
rect 9088 30812 9094 30864
rect 9232 30725 9260 30892
rect 12406 30852 12434 30892
rect 14090 30880 14096 30932
rect 14148 30920 14154 30932
rect 39025 30923 39083 30929
rect 39025 30920 39037 30923
rect 14148 30892 39037 30920
rect 14148 30880 14154 30892
rect 39025 30889 39037 30892
rect 39071 30920 39083 30923
rect 40037 30923 40095 30929
rect 40037 30920 40049 30923
rect 39071 30892 40049 30920
rect 39071 30889 39083 30892
rect 39025 30883 39083 30889
rect 40037 30889 40049 30892
rect 40083 30889 40095 30923
rect 40037 30883 40095 30889
rect 14550 30852 14556 30864
rect 12406 30824 14556 30852
rect 14550 30812 14556 30824
rect 14608 30852 14614 30864
rect 21174 30852 21180 30864
rect 14608 30824 21180 30852
rect 14608 30812 14614 30824
rect 21174 30812 21180 30824
rect 21232 30812 21238 30864
rect 9490 30744 9496 30796
rect 9548 30784 9554 30796
rect 9548 30756 10548 30784
rect 9548 30744 9554 30756
rect 9217 30719 9275 30725
rect 9217 30685 9229 30719
rect 9263 30685 9275 30719
rect 9217 30679 9275 30685
rect 9324 30688 10088 30716
rect 10520 30702 10548 30756
rect 11606 30744 11612 30796
rect 11664 30784 11670 30796
rect 11885 30787 11943 30793
rect 11885 30784 11897 30787
rect 11664 30756 11897 30784
rect 11664 30744 11670 30756
rect 11885 30753 11897 30756
rect 11931 30753 11943 30787
rect 11885 30747 11943 30753
rect 6454 30608 6460 30660
rect 6512 30648 6518 30660
rect 9324 30648 9352 30688
rect 9861 30651 9919 30657
rect 9861 30648 9873 30651
rect 6512 30620 9352 30648
rect 9416 30620 9873 30648
rect 6512 30608 6518 30620
rect 5626 30540 5632 30592
rect 5684 30580 5690 30592
rect 6270 30580 6276 30592
rect 5684 30552 6276 30580
rect 5684 30540 5690 30552
rect 6270 30540 6276 30552
rect 6328 30580 6334 30592
rect 9416 30580 9444 30620
rect 9861 30617 9873 30620
rect 9907 30617 9919 30651
rect 9861 30611 9919 30617
rect 6328 30552 9444 30580
rect 10060 30580 10088 30688
rect 33226 30676 33232 30728
rect 33284 30716 33290 30728
rect 34146 30716 34152 30728
rect 33284 30688 34152 30716
rect 33284 30676 33290 30688
rect 34146 30676 34152 30688
rect 34204 30716 34210 30728
rect 39393 30719 39451 30725
rect 39393 30716 39405 30719
rect 34204 30688 39405 30716
rect 34204 30676 34210 30688
rect 39393 30685 39405 30688
rect 39439 30716 39451 30719
rect 39439 30688 39896 30716
rect 39439 30685 39451 30688
rect 39393 30679 39451 30685
rect 11330 30608 11336 30660
rect 11388 30648 11394 30660
rect 39868 30657 39896 30688
rect 11609 30651 11667 30657
rect 11609 30648 11621 30651
rect 11388 30620 11621 30648
rect 11388 30608 11394 30620
rect 11609 30617 11621 30620
rect 11655 30617 11667 30651
rect 39853 30651 39911 30657
rect 11609 30611 11667 30617
rect 38028 30620 39528 30648
rect 38028 30580 38056 30620
rect 10060 30552 38056 30580
rect 39500 30580 39528 30620
rect 39853 30617 39865 30651
rect 39899 30617 39911 30651
rect 39853 30611 39911 30617
rect 40034 30608 40040 30660
rect 40092 30608 40098 30660
rect 40221 30583 40279 30589
rect 40221 30580 40233 30583
rect 39500 30552 40233 30580
rect 6328 30540 6334 30552
rect 40221 30549 40233 30552
rect 40267 30549 40279 30583
rect 40221 30543 40279 30549
rect 1104 30490 40848 30512
rect 1104 30438 2610 30490
rect 2662 30438 2674 30490
rect 2726 30438 2738 30490
rect 2790 30438 2802 30490
rect 2854 30438 2866 30490
rect 2918 30438 7610 30490
rect 7662 30438 7674 30490
rect 7726 30438 7738 30490
rect 7790 30438 7802 30490
rect 7854 30438 7866 30490
rect 7918 30438 12610 30490
rect 12662 30438 12674 30490
rect 12726 30438 12738 30490
rect 12790 30438 12802 30490
rect 12854 30438 12866 30490
rect 12918 30438 17610 30490
rect 17662 30438 17674 30490
rect 17726 30438 17738 30490
rect 17790 30438 17802 30490
rect 17854 30438 17866 30490
rect 17918 30438 22610 30490
rect 22662 30438 22674 30490
rect 22726 30438 22738 30490
rect 22790 30438 22802 30490
rect 22854 30438 22866 30490
rect 22918 30438 27610 30490
rect 27662 30438 27674 30490
rect 27726 30438 27738 30490
rect 27790 30438 27802 30490
rect 27854 30438 27866 30490
rect 27918 30438 32610 30490
rect 32662 30438 32674 30490
rect 32726 30438 32738 30490
rect 32790 30438 32802 30490
rect 32854 30438 32866 30490
rect 32918 30438 37610 30490
rect 37662 30438 37674 30490
rect 37726 30438 37738 30490
rect 37790 30438 37802 30490
rect 37854 30438 37866 30490
rect 37918 30438 40848 30490
rect 1104 30416 40848 30438
rect 3050 30336 3056 30388
rect 3108 30376 3114 30388
rect 11330 30376 11336 30388
rect 3108 30348 11336 30376
rect 3108 30336 3114 30348
rect 11330 30336 11336 30348
rect 11388 30336 11394 30388
rect 11514 30268 11520 30320
rect 11572 30308 11578 30320
rect 11885 30311 11943 30317
rect 11885 30308 11897 30311
rect 11572 30280 11897 30308
rect 11572 30268 11578 30280
rect 11885 30277 11897 30280
rect 11931 30277 11943 30311
rect 11885 30271 11943 30277
rect 22462 30268 22468 30320
rect 22520 30308 22526 30320
rect 23014 30308 23020 30320
rect 22520 30280 23020 30308
rect 22520 30268 22526 30280
rect 23014 30268 23020 30280
rect 23072 30308 23078 30320
rect 32398 30308 32404 30320
rect 23072 30280 32404 30308
rect 23072 30268 23078 30280
rect 32398 30268 32404 30280
rect 32456 30268 32462 30320
rect 11698 30200 11704 30252
rect 11756 30200 11762 30252
rect 18233 30243 18291 30249
rect 18233 30240 18245 30243
rect 12406 30212 18245 30240
rect 5074 30132 5080 30184
rect 5132 30172 5138 30184
rect 12406 30172 12434 30212
rect 18233 30209 18245 30212
rect 18279 30240 18291 30243
rect 18874 30240 18880 30252
rect 18279 30212 18880 30240
rect 18279 30209 18291 30212
rect 18233 30203 18291 30209
rect 18874 30200 18880 30212
rect 18932 30200 18938 30252
rect 5132 30144 12434 30172
rect 18141 30175 18199 30181
rect 5132 30132 5138 30144
rect 18141 30141 18153 30175
rect 18187 30172 18199 30175
rect 18598 30172 18604 30184
rect 18187 30144 18604 30172
rect 18187 30141 18199 30144
rect 18141 30135 18199 30141
rect 18598 30132 18604 30144
rect 18656 30172 18662 30184
rect 18782 30172 18788 30184
rect 18656 30144 18788 30172
rect 18656 30132 18662 30144
rect 18782 30132 18788 30144
rect 18840 30132 18846 30184
rect 12069 30107 12127 30113
rect 12069 30073 12081 30107
rect 12115 30104 12127 30107
rect 28626 30104 28632 30116
rect 12115 30076 28632 30104
rect 12115 30073 12127 30076
rect 12069 30067 12127 30073
rect 28626 30064 28632 30076
rect 28684 30064 28690 30116
rect 16850 29996 16856 30048
rect 16908 30036 16914 30048
rect 18414 30036 18420 30048
rect 16908 30008 18420 30036
rect 16908 29996 16914 30008
rect 18414 29996 18420 30008
rect 18472 29996 18478 30048
rect 28994 29996 29000 30048
rect 29052 30036 29058 30048
rect 29270 30036 29276 30048
rect 29052 30008 29276 30036
rect 29052 29996 29058 30008
rect 29270 29996 29276 30008
rect 29328 29996 29334 30048
rect 1104 29946 40848 29968
rect 1104 29894 1950 29946
rect 2002 29894 2014 29946
rect 2066 29894 2078 29946
rect 2130 29894 2142 29946
rect 2194 29894 2206 29946
rect 2258 29894 6950 29946
rect 7002 29894 7014 29946
rect 7066 29894 7078 29946
rect 7130 29894 7142 29946
rect 7194 29894 7206 29946
rect 7258 29894 11950 29946
rect 12002 29894 12014 29946
rect 12066 29894 12078 29946
rect 12130 29894 12142 29946
rect 12194 29894 12206 29946
rect 12258 29894 16950 29946
rect 17002 29894 17014 29946
rect 17066 29894 17078 29946
rect 17130 29894 17142 29946
rect 17194 29894 17206 29946
rect 17258 29894 21950 29946
rect 22002 29894 22014 29946
rect 22066 29894 22078 29946
rect 22130 29894 22142 29946
rect 22194 29894 22206 29946
rect 22258 29894 26950 29946
rect 27002 29894 27014 29946
rect 27066 29894 27078 29946
rect 27130 29894 27142 29946
rect 27194 29894 27206 29946
rect 27258 29894 31950 29946
rect 32002 29894 32014 29946
rect 32066 29894 32078 29946
rect 32130 29894 32142 29946
rect 32194 29894 32206 29946
rect 32258 29894 36950 29946
rect 37002 29894 37014 29946
rect 37066 29894 37078 29946
rect 37130 29894 37142 29946
rect 37194 29894 37206 29946
rect 37258 29894 40848 29946
rect 1104 29872 40848 29894
rect 3970 29792 3976 29844
rect 4028 29832 4034 29844
rect 8205 29835 8263 29841
rect 8205 29832 8217 29835
rect 4028 29804 8217 29832
rect 4028 29792 4034 29804
rect 8205 29801 8217 29804
rect 8251 29801 8263 29835
rect 8205 29795 8263 29801
rect 8478 29792 8484 29844
rect 8536 29832 8542 29844
rect 17402 29832 17408 29844
rect 8536 29804 17408 29832
rect 8536 29792 8542 29804
rect 17402 29792 17408 29804
rect 17460 29792 17466 29844
rect 18414 29792 18420 29844
rect 18472 29832 18478 29844
rect 31018 29832 31024 29844
rect 18472 29804 31024 29832
rect 18472 29792 18478 29804
rect 31018 29792 31024 29804
rect 31076 29792 31082 29844
rect 3878 29656 3884 29708
rect 3936 29696 3942 29708
rect 8021 29699 8079 29705
rect 8021 29696 8033 29699
rect 3936 29668 8033 29696
rect 3936 29656 3942 29668
rect 8021 29665 8033 29668
rect 8067 29696 8079 29699
rect 11606 29696 11612 29708
rect 8067 29668 11612 29696
rect 8067 29665 8079 29668
rect 8021 29659 8079 29665
rect 11606 29656 11612 29668
rect 11664 29656 11670 29708
rect 14182 29696 14188 29708
rect 12406 29668 14188 29696
rect 5997 29631 6055 29637
rect 5997 29597 6009 29631
rect 6043 29628 6055 29631
rect 6178 29628 6184 29640
rect 6043 29600 6184 29628
rect 6043 29597 6055 29600
rect 5997 29591 6055 29597
rect 6178 29588 6184 29600
rect 6236 29588 6242 29640
rect 8294 29588 8300 29640
rect 8352 29628 8358 29640
rect 12406 29628 12434 29668
rect 14182 29656 14188 29668
rect 14240 29656 14246 29708
rect 14274 29656 14280 29708
rect 14332 29696 14338 29708
rect 14461 29699 14519 29705
rect 14461 29696 14473 29699
rect 14332 29668 14473 29696
rect 14332 29656 14338 29668
rect 14461 29665 14473 29668
rect 14507 29665 14519 29699
rect 14461 29659 14519 29665
rect 8352 29600 12434 29628
rect 8352 29588 8358 29600
rect 13906 29588 13912 29640
rect 13964 29628 13970 29640
rect 14093 29631 14151 29637
rect 14093 29628 14105 29631
rect 13964 29600 14105 29628
rect 13964 29588 13970 29600
rect 14093 29597 14105 29600
rect 14139 29597 14151 29631
rect 15286 29628 15292 29640
rect 14093 29591 14151 29597
rect 14200 29600 15292 29628
rect 6086 29520 6092 29572
rect 6144 29560 6150 29572
rect 7745 29563 7803 29569
rect 6144 29532 6578 29560
rect 6144 29520 6150 29532
rect 7745 29529 7757 29563
rect 7791 29560 7803 29563
rect 14200 29560 14228 29600
rect 15286 29588 15292 29600
rect 15344 29588 15350 29640
rect 7791 29532 14228 29560
rect 7791 29529 7803 29532
rect 7745 29523 7803 29529
rect 6454 29452 6460 29504
rect 6512 29492 6518 29504
rect 8478 29492 8484 29504
rect 6512 29464 8484 29492
rect 6512 29452 6518 29464
rect 8478 29452 8484 29464
rect 8536 29452 8542 29504
rect 1104 29402 40848 29424
rect 1104 29350 2610 29402
rect 2662 29350 2674 29402
rect 2726 29350 2738 29402
rect 2790 29350 2802 29402
rect 2854 29350 2866 29402
rect 2918 29350 7610 29402
rect 7662 29350 7674 29402
rect 7726 29350 7738 29402
rect 7790 29350 7802 29402
rect 7854 29350 7866 29402
rect 7918 29350 12610 29402
rect 12662 29350 12674 29402
rect 12726 29350 12738 29402
rect 12790 29350 12802 29402
rect 12854 29350 12866 29402
rect 12918 29350 17610 29402
rect 17662 29350 17674 29402
rect 17726 29350 17738 29402
rect 17790 29350 17802 29402
rect 17854 29350 17866 29402
rect 17918 29350 22610 29402
rect 22662 29350 22674 29402
rect 22726 29350 22738 29402
rect 22790 29350 22802 29402
rect 22854 29350 22866 29402
rect 22918 29350 27610 29402
rect 27662 29350 27674 29402
rect 27726 29350 27738 29402
rect 27790 29350 27802 29402
rect 27854 29350 27866 29402
rect 27918 29350 32610 29402
rect 32662 29350 32674 29402
rect 32726 29350 32738 29402
rect 32790 29350 32802 29402
rect 32854 29350 32866 29402
rect 32918 29350 37610 29402
rect 37662 29350 37674 29402
rect 37726 29350 37738 29402
rect 37790 29350 37802 29402
rect 37854 29350 37866 29402
rect 37918 29350 40848 29402
rect 1104 29328 40848 29350
rect 15378 29288 15384 29300
rect 5920 29260 15384 29288
rect 5920 29229 5948 29260
rect 15378 29248 15384 29260
rect 15436 29248 15442 29300
rect 33686 29288 33692 29300
rect 17420 29260 33692 29288
rect 5905 29223 5963 29229
rect 5905 29189 5917 29223
rect 5951 29189 5963 29223
rect 14458 29220 14464 29232
rect 5905 29183 5963 29189
rect 7392 29192 14464 29220
rect 7392 29164 7420 29192
rect 14458 29180 14464 29192
rect 14516 29180 14522 29232
rect 17420 29229 17448 29260
rect 33686 29248 33692 29260
rect 33744 29248 33750 29300
rect 17405 29223 17463 29229
rect 17405 29189 17417 29223
rect 17451 29189 17463 29223
rect 17954 29220 17960 29232
rect 17405 29183 17463 29189
rect 17880 29192 17960 29220
rect 3878 29112 3884 29164
rect 3936 29112 3942 29164
rect 5258 29112 5264 29164
rect 5316 29112 5322 29164
rect 7285 29155 7343 29161
rect 7285 29121 7297 29155
rect 7331 29152 7343 29155
rect 7374 29152 7380 29164
rect 7331 29124 7380 29152
rect 7331 29121 7343 29124
rect 7285 29115 7343 29121
rect 7374 29112 7380 29124
rect 7432 29112 7438 29164
rect 12434 29112 12440 29164
rect 12492 29152 12498 29164
rect 16850 29152 16856 29164
rect 12492 29124 16856 29152
rect 12492 29112 12498 29124
rect 16850 29112 16856 29124
rect 16908 29152 16914 29164
rect 17037 29155 17095 29161
rect 17037 29152 17049 29155
rect 16908 29124 17049 29152
rect 16908 29112 16914 29124
rect 17037 29121 17049 29124
rect 17083 29121 17095 29155
rect 17037 29115 17095 29121
rect 17313 29155 17371 29161
rect 17313 29121 17325 29155
rect 17359 29152 17371 29155
rect 17880 29152 17908 29192
rect 17954 29180 17960 29192
rect 18012 29220 18018 29232
rect 18414 29220 18420 29232
rect 18012 29192 18420 29220
rect 18012 29180 18018 29192
rect 18414 29180 18420 29192
rect 18472 29180 18478 29232
rect 18506 29180 18512 29232
rect 18564 29180 18570 29232
rect 20714 29220 20720 29232
rect 19734 29192 20720 29220
rect 20714 29180 20720 29192
rect 20772 29180 20778 29232
rect 17359 29124 17908 29152
rect 20257 29155 20315 29161
rect 17359 29121 17371 29124
rect 17313 29115 17371 29121
rect 20257 29121 20269 29155
rect 20303 29152 20315 29155
rect 23014 29152 23020 29164
rect 20303 29124 23020 29152
rect 20303 29121 20315 29124
rect 20257 29115 20315 29121
rect 23014 29112 23020 29124
rect 23072 29112 23078 29164
rect 40218 29112 40224 29164
rect 40276 29152 40282 29164
rect 40313 29155 40371 29161
rect 40313 29152 40325 29155
rect 40276 29124 40325 29152
rect 40276 29112 40282 29124
rect 40313 29121 40325 29124
rect 40359 29121 40371 29155
rect 40313 29115 40371 29121
rect 3605 29087 3663 29093
rect 3605 29053 3617 29087
rect 3651 29084 3663 29087
rect 4157 29087 4215 29093
rect 4157 29084 4169 29087
rect 3651 29056 4169 29084
rect 3651 29053 3663 29056
rect 3605 29047 3663 29053
rect 4157 29053 4169 29056
rect 4203 29084 4215 29087
rect 4798 29084 4804 29096
rect 4203 29056 4804 29084
rect 4203 29053 4215 29056
rect 4157 29047 4215 29053
rect 4798 29044 4804 29056
rect 4856 29044 4862 29096
rect 6454 29044 6460 29096
rect 6512 29044 6518 29096
rect 18138 29044 18144 29096
rect 18196 29084 18202 29096
rect 18233 29087 18291 29093
rect 18233 29084 18245 29087
rect 18196 29056 18245 29084
rect 18196 29044 18202 29056
rect 18233 29053 18245 29056
rect 18279 29053 18291 29087
rect 26786 29084 26792 29096
rect 18233 29047 18291 29053
rect 26206 29056 26792 29084
rect 19518 28976 19524 29028
rect 19576 29016 19582 29028
rect 26206 29016 26234 29056
rect 26786 29044 26792 29056
rect 26844 29084 26850 29096
rect 39669 29087 39727 29093
rect 39669 29084 39681 29087
rect 26844 29056 39681 29084
rect 26844 29044 26850 29056
rect 39669 29053 39681 29056
rect 39715 29053 39727 29087
rect 39669 29047 39727 29053
rect 19576 28988 26234 29016
rect 19576 28976 19582 28988
rect 1104 28858 40848 28880
rect 1104 28806 1950 28858
rect 2002 28806 2014 28858
rect 2066 28806 2078 28858
rect 2130 28806 2142 28858
rect 2194 28806 2206 28858
rect 2258 28806 6950 28858
rect 7002 28806 7014 28858
rect 7066 28806 7078 28858
rect 7130 28806 7142 28858
rect 7194 28806 7206 28858
rect 7258 28806 11950 28858
rect 12002 28806 12014 28858
rect 12066 28806 12078 28858
rect 12130 28806 12142 28858
rect 12194 28806 12206 28858
rect 12258 28806 16950 28858
rect 17002 28806 17014 28858
rect 17066 28806 17078 28858
rect 17130 28806 17142 28858
rect 17194 28806 17206 28858
rect 17258 28806 21950 28858
rect 22002 28806 22014 28858
rect 22066 28806 22078 28858
rect 22130 28806 22142 28858
rect 22194 28806 22206 28858
rect 22258 28806 26950 28858
rect 27002 28806 27014 28858
rect 27066 28806 27078 28858
rect 27130 28806 27142 28858
rect 27194 28806 27206 28858
rect 27258 28806 31950 28858
rect 32002 28806 32014 28858
rect 32066 28806 32078 28858
rect 32130 28806 32142 28858
rect 32194 28806 32206 28858
rect 32258 28806 36950 28858
rect 37002 28806 37014 28858
rect 37066 28806 37078 28858
rect 37130 28806 37142 28858
rect 37194 28806 37206 28858
rect 37258 28806 40848 28858
rect 1104 28784 40848 28806
rect 17954 28636 17960 28688
rect 18012 28676 18018 28688
rect 19150 28676 19156 28688
rect 18012 28648 19156 28676
rect 18012 28636 18018 28648
rect 19150 28636 19156 28648
rect 19208 28676 19214 28688
rect 19208 28648 26234 28676
rect 19208 28636 19214 28648
rect 19245 28611 19303 28617
rect 19245 28577 19257 28611
rect 19291 28608 19303 28611
rect 19978 28608 19984 28620
rect 19291 28580 19984 28608
rect 19291 28577 19303 28580
rect 19245 28571 19303 28577
rect 19978 28568 19984 28580
rect 20036 28568 20042 28620
rect 4617 28543 4675 28549
rect 4617 28509 4629 28543
rect 4663 28540 4675 28543
rect 8294 28540 8300 28552
rect 4663 28512 8300 28540
rect 4663 28509 4675 28512
rect 4617 28503 4675 28509
rect 8294 28500 8300 28512
rect 8352 28500 8358 28552
rect 11514 28500 11520 28552
rect 11572 28540 11578 28552
rect 19613 28543 19671 28549
rect 19613 28540 19625 28543
rect 11572 28512 19625 28540
rect 11572 28500 11578 28512
rect 19613 28509 19625 28512
rect 19659 28509 19671 28543
rect 19613 28503 19671 28509
rect 11698 28432 11704 28484
rect 11756 28472 11762 28484
rect 19628 28472 19656 28503
rect 19794 28500 19800 28552
rect 19852 28500 19858 28552
rect 26206 28540 26234 28648
rect 30558 28636 30564 28688
rect 30616 28636 30622 28688
rect 29454 28568 29460 28620
rect 29512 28608 29518 28620
rect 29825 28611 29883 28617
rect 29825 28608 29837 28611
rect 29512 28580 29837 28608
rect 29512 28568 29518 28580
rect 29825 28577 29837 28580
rect 29871 28608 29883 28611
rect 33594 28608 33600 28620
rect 29871 28580 33600 28608
rect 29871 28577 29883 28580
rect 29825 28571 29883 28577
rect 33594 28568 33600 28580
rect 33652 28568 33658 28620
rect 30101 28543 30159 28549
rect 30101 28540 30113 28543
rect 26206 28512 30113 28540
rect 30101 28509 30113 28512
rect 30147 28509 30159 28543
rect 30101 28503 30159 28509
rect 30653 28543 30711 28549
rect 30653 28509 30665 28543
rect 30699 28540 30711 28543
rect 31570 28540 31576 28552
rect 30699 28512 31576 28540
rect 30699 28509 30711 28512
rect 30653 28503 30711 28509
rect 22002 28472 22008 28484
rect 11756 28444 19472 28472
rect 19628 28444 22008 28472
rect 11756 28432 11762 28444
rect 4709 28407 4767 28413
rect 4709 28373 4721 28407
rect 4755 28404 4767 28407
rect 8202 28404 8208 28416
rect 4755 28376 8208 28404
rect 4755 28373 4767 28376
rect 4709 28367 4767 28373
rect 8202 28364 8208 28376
rect 8260 28364 8266 28416
rect 8294 28364 8300 28416
rect 8352 28404 8358 28416
rect 17954 28404 17960 28416
rect 8352 28376 17960 28404
rect 8352 28364 8358 28376
rect 17954 28364 17960 28376
rect 18012 28364 18018 28416
rect 19334 28364 19340 28416
rect 19392 28364 19398 28416
rect 19444 28404 19472 28444
rect 22002 28432 22008 28444
rect 22060 28432 22066 28484
rect 30116 28472 30144 28503
rect 31570 28500 31576 28512
rect 31628 28500 31634 28552
rect 31846 28472 31852 28484
rect 30116 28444 31852 28472
rect 31846 28432 31852 28444
rect 31904 28432 31910 28484
rect 19794 28404 19800 28416
rect 19444 28376 19800 28404
rect 19794 28364 19800 28376
rect 19852 28404 19858 28416
rect 20438 28404 20444 28416
rect 19852 28376 20444 28404
rect 19852 28364 19858 28376
rect 20438 28364 20444 28376
rect 20496 28364 20502 28416
rect 1104 28314 40848 28336
rect 1104 28262 2610 28314
rect 2662 28262 2674 28314
rect 2726 28262 2738 28314
rect 2790 28262 2802 28314
rect 2854 28262 2866 28314
rect 2918 28262 7610 28314
rect 7662 28262 7674 28314
rect 7726 28262 7738 28314
rect 7790 28262 7802 28314
rect 7854 28262 7866 28314
rect 7918 28262 12610 28314
rect 12662 28262 12674 28314
rect 12726 28262 12738 28314
rect 12790 28262 12802 28314
rect 12854 28262 12866 28314
rect 12918 28262 17610 28314
rect 17662 28262 17674 28314
rect 17726 28262 17738 28314
rect 17790 28262 17802 28314
rect 17854 28262 17866 28314
rect 17918 28262 22610 28314
rect 22662 28262 22674 28314
rect 22726 28262 22738 28314
rect 22790 28262 22802 28314
rect 22854 28262 22866 28314
rect 22918 28262 27610 28314
rect 27662 28262 27674 28314
rect 27726 28262 27738 28314
rect 27790 28262 27802 28314
rect 27854 28262 27866 28314
rect 27918 28262 32610 28314
rect 32662 28262 32674 28314
rect 32726 28262 32738 28314
rect 32790 28262 32802 28314
rect 32854 28262 32866 28314
rect 32918 28262 37610 28314
rect 37662 28262 37674 28314
rect 37726 28262 37738 28314
rect 37790 28262 37802 28314
rect 37854 28262 37866 28314
rect 37918 28262 40848 28314
rect 1104 28240 40848 28262
rect 22005 28203 22063 28209
rect 22005 28169 22017 28203
rect 22051 28200 22063 28203
rect 29086 28200 29092 28212
rect 22051 28172 29092 28200
rect 22051 28169 22063 28172
rect 22005 28163 22063 28169
rect 29086 28160 29092 28172
rect 29144 28160 29150 28212
rect 29546 28160 29552 28212
rect 29604 28160 29610 28212
rect 31846 28160 31852 28212
rect 31904 28200 31910 28212
rect 32398 28200 32404 28212
rect 31904 28172 32404 28200
rect 31904 28160 31910 28172
rect 32398 28160 32404 28172
rect 32456 28160 32462 28212
rect 17494 28092 17500 28144
rect 17552 28132 17558 28144
rect 29270 28132 29276 28144
rect 17552 28104 29276 28132
rect 17552 28092 17558 28104
rect 29270 28092 29276 28104
rect 29328 28132 29334 28144
rect 29365 28135 29423 28141
rect 29365 28132 29377 28135
rect 29328 28104 29377 28132
rect 29328 28092 29334 28104
rect 29365 28101 29377 28104
rect 29411 28132 29423 28135
rect 29825 28135 29883 28141
rect 29825 28132 29837 28135
rect 29411 28104 29837 28132
rect 29411 28101 29423 28104
rect 29365 28095 29423 28101
rect 29825 28101 29837 28104
rect 29871 28101 29883 28135
rect 29825 28095 29883 28101
rect 20438 28024 20444 28076
rect 20496 28064 20502 28076
rect 21821 28067 21879 28073
rect 21821 28064 21833 28067
rect 20496 28036 21833 28064
rect 20496 28024 20502 28036
rect 21821 28033 21833 28036
rect 21867 28033 21879 28067
rect 21821 28027 21879 28033
rect 22002 28024 22008 28076
rect 22060 28064 22066 28076
rect 22281 28067 22339 28073
rect 22281 28064 22293 28067
rect 22060 28036 22293 28064
rect 22060 28024 22066 28036
rect 22281 28033 22293 28036
rect 22327 28064 22339 28067
rect 22327 28036 26096 28064
rect 22327 28033 22339 28036
rect 22281 28027 22339 28033
rect 9858 27888 9864 27940
rect 9916 27928 9922 27940
rect 10594 27928 10600 27940
rect 9916 27900 10600 27928
rect 9916 27888 9922 27900
rect 10594 27888 10600 27900
rect 10652 27928 10658 27940
rect 26068 27928 26096 28036
rect 29086 28024 29092 28076
rect 29144 28064 29150 28076
rect 29181 28067 29239 28073
rect 29181 28064 29193 28067
rect 29144 28036 29193 28064
rect 29144 28024 29150 28036
rect 29181 28033 29193 28036
rect 29227 28033 29239 28067
rect 29181 28027 29239 28033
rect 38562 27928 38568 27940
rect 10652 27900 22416 27928
rect 26068 27900 38568 27928
rect 10652 27888 10658 27900
rect 22388 27860 22416 27900
rect 38562 27888 38568 27900
rect 38620 27888 38626 27940
rect 28813 27863 28871 27869
rect 28813 27860 28825 27863
rect 22388 27832 28825 27860
rect 28813 27829 28825 27832
rect 28859 27860 28871 27863
rect 29086 27860 29092 27872
rect 28859 27832 29092 27860
rect 28859 27829 28871 27832
rect 28813 27823 28871 27829
rect 29086 27820 29092 27832
rect 29144 27820 29150 27872
rect 1104 27770 40848 27792
rect 1104 27718 1950 27770
rect 2002 27718 2014 27770
rect 2066 27718 2078 27770
rect 2130 27718 2142 27770
rect 2194 27718 2206 27770
rect 2258 27718 6950 27770
rect 7002 27718 7014 27770
rect 7066 27718 7078 27770
rect 7130 27718 7142 27770
rect 7194 27718 7206 27770
rect 7258 27718 11950 27770
rect 12002 27718 12014 27770
rect 12066 27718 12078 27770
rect 12130 27718 12142 27770
rect 12194 27718 12206 27770
rect 12258 27718 16950 27770
rect 17002 27718 17014 27770
rect 17066 27718 17078 27770
rect 17130 27718 17142 27770
rect 17194 27718 17206 27770
rect 17258 27718 21950 27770
rect 22002 27718 22014 27770
rect 22066 27718 22078 27770
rect 22130 27718 22142 27770
rect 22194 27718 22206 27770
rect 22258 27718 26950 27770
rect 27002 27718 27014 27770
rect 27066 27718 27078 27770
rect 27130 27718 27142 27770
rect 27194 27718 27206 27770
rect 27258 27718 31950 27770
rect 32002 27718 32014 27770
rect 32066 27718 32078 27770
rect 32130 27718 32142 27770
rect 32194 27718 32206 27770
rect 32258 27718 36950 27770
rect 37002 27718 37014 27770
rect 37066 27718 37078 27770
rect 37130 27718 37142 27770
rect 37194 27718 37206 27770
rect 37258 27718 40848 27770
rect 1104 27696 40848 27718
rect 17607 27659 17665 27665
rect 17607 27625 17619 27659
rect 17653 27656 17665 27659
rect 22462 27656 22468 27668
rect 17653 27628 22468 27656
rect 17653 27625 17665 27628
rect 17607 27619 17665 27625
rect 22462 27616 22468 27628
rect 22520 27616 22526 27668
rect 19978 27548 19984 27600
rect 20036 27588 20042 27600
rect 28994 27588 29000 27600
rect 20036 27560 29000 27588
rect 20036 27548 20042 27560
rect 28994 27548 29000 27560
rect 29052 27588 29058 27600
rect 31662 27588 31668 27600
rect 29052 27560 31668 27588
rect 29052 27548 29058 27560
rect 31662 27548 31668 27560
rect 31720 27548 31726 27600
rect 12342 27480 12348 27532
rect 12400 27520 12406 27532
rect 12400 27492 20300 27520
rect 12400 27480 12406 27492
rect 17865 27455 17923 27461
rect 17865 27421 17877 27455
rect 17911 27452 17923 27455
rect 18138 27452 18144 27464
rect 17911 27424 18144 27452
rect 17911 27421 17923 27424
rect 17865 27415 17923 27421
rect 18138 27412 18144 27424
rect 18196 27412 18202 27464
rect 19978 27412 19984 27464
rect 20036 27412 20042 27464
rect 20272 27461 20300 27492
rect 20438 27480 20444 27532
rect 20496 27480 20502 27532
rect 20257 27455 20315 27461
rect 20257 27421 20269 27455
rect 20303 27421 20315 27455
rect 20257 27415 20315 27421
rect 15838 27344 15844 27396
rect 15896 27344 15902 27396
rect 32490 27384 32496 27396
rect 17158 27356 17540 27384
rect 15565 27319 15623 27325
rect 15565 27285 15577 27319
rect 15611 27316 15623 27319
rect 17236 27316 17264 27356
rect 15611 27288 17264 27316
rect 17512 27316 17540 27356
rect 17696 27356 32496 27384
rect 17696 27316 17724 27356
rect 32490 27344 32496 27356
rect 32548 27344 32554 27396
rect 17512 27288 17724 27316
rect 20533 27319 20591 27325
rect 15611 27285 15623 27288
rect 15565 27279 15623 27285
rect 20533 27285 20545 27319
rect 20579 27316 20591 27319
rect 38010 27316 38016 27328
rect 20579 27288 38016 27316
rect 20579 27285 20591 27288
rect 20533 27279 20591 27285
rect 38010 27276 38016 27288
rect 38068 27276 38074 27328
rect 1104 27226 40848 27248
rect 1104 27174 2610 27226
rect 2662 27174 2674 27226
rect 2726 27174 2738 27226
rect 2790 27174 2802 27226
rect 2854 27174 2866 27226
rect 2918 27174 7610 27226
rect 7662 27174 7674 27226
rect 7726 27174 7738 27226
rect 7790 27174 7802 27226
rect 7854 27174 7866 27226
rect 7918 27174 12610 27226
rect 12662 27174 12674 27226
rect 12726 27174 12738 27226
rect 12790 27174 12802 27226
rect 12854 27174 12866 27226
rect 12918 27174 17610 27226
rect 17662 27174 17674 27226
rect 17726 27174 17738 27226
rect 17790 27174 17802 27226
rect 17854 27174 17866 27226
rect 17918 27174 22610 27226
rect 22662 27174 22674 27226
rect 22726 27174 22738 27226
rect 22790 27174 22802 27226
rect 22854 27174 22866 27226
rect 22918 27174 27610 27226
rect 27662 27174 27674 27226
rect 27726 27174 27738 27226
rect 27790 27174 27802 27226
rect 27854 27174 27866 27226
rect 27918 27174 32610 27226
rect 32662 27174 32674 27226
rect 32726 27174 32738 27226
rect 32790 27174 32802 27226
rect 32854 27174 32866 27226
rect 32918 27174 37610 27226
rect 37662 27174 37674 27226
rect 37726 27174 37738 27226
rect 37790 27174 37802 27226
rect 37854 27174 37866 27226
rect 37918 27174 40848 27226
rect 1104 27152 40848 27174
rect 8386 27072 8392 27124
rect 8444 27112 8450 27124
rect 14274 27112 14280 27124
rect 8444 27084 14280 27112
rect 8444 27072 8450 27084
rect 14274 27072 14280 27084
rect 14332 27112 14338 27124
rect 19978 27112 19984 27124
rect 14332 27084 19984 27112
rect 14332 27072 14338 27084
rect 19978 27072 19984 27084
rect 20036 27072 20042 27124
rect 8941 27047 8999 27053
rect 8941 27013 8953 27047
rect 8987 27044 8999 27047
rect 18046 27044 18052 27056
rect 8987 27016 18052 27044
rect 8987 27013 8999 27016
rect 8941 27007 8999 27013
rect 18046 27004 18052 27016
rect 18104 27004 18110 27056
rect 8662 26936 8668 26988
rect 8720 26976 8726 26988
rect 9125 26979 9183 26985
rect 9125 26976 9137 26979
rect 8720 26948 9137 26976
rect 8720 26936 8726 26948
rect 9125 26945 9137 26948
rect 9171 26945 9183 26979
rect 9125 26939 9183 26945
rect 9214 26732 9220 26784
rect 9272 26732 9278 26784
rect 1104 26682 40848 26704
rect 1104 26630 1950 26682
rect 2002 26630 2014 26682
rect 2066 26630 2078 26682
rect 2130 26630 2142 26682
rect 2194 26630 2206 26682
rect 2258 26630 6950 26682
rect 7002 26630 7014 26682
rect 7066 26630 7078 26682
rect 7130 26630 7142 26682
rect 7194 26630 7206 26682
rect 7258 26630 11950 26682
rect 12002 26630 12014 26682
rect 12066 26630 12078 26682
rect 12130 26630 12142 26682
rect 12194 26630 12206 26682
rect 12258 26630 16950 26682
rect 17002 26630 17014 26682
rect 17066 26630 17078 26682
rect 17130 26630 17142 26682
rect 17194 26630 17206 26682
rect 17258 26630 21950 26682
rect 22002 26630 22014 26682
rect 22066 26630 22078 26682
rect 22130 26630 22142 26682
rect 22194 26630 22206 26682
rect 22258 26630 26950 26682
rect 27002 26630 27014 26682
rect 27066 26630 27078 26682
rect 27130 26630 27142 26682
rect 27194 26630 27206 26682
rect 27258 26630 31950 26682
rect 32002 26630 32014 26682
rect 32066 26630 32078 26682
rect 32130 26630 32142 26682
rect 32194 26630 32206 26682
rect 32258 26630 36950 26682
rect 37002 26630 37014 26682
rect 37066 26630 37078 26682
rect 37130 26630 37142 26682
rect 37194 26630 37206 26682
rect 37258 26630 40848 26682
rect 1104 26608 40848 26630
rect 1104 26138 40848 26160
rect 1104 26086 2610 26138
rect 2662 26086 2674 26138
rect 2726 26086 2738 26138
rect 2790 26086 2802 26138
rect 2854 26086 2866 26138
rect 2918 26086 7610 26138
rect 7662 26086 7674 26138
rect 7726 26086 7738 26138
rect 7790 26086 7802 26138
rect 7854 26086 7866 26138
rect 7918 26086 12610 26138
rect 12662 26086 12674 26138
rect 12726 26086 12738 26138
rect 12790 26086 12802 26138
rect 12854 26086 12866 26138
rect 12918 26086 17610 26138
rect 17662 26086 17674 26138
rect 17726 26086 17738 26138
rect 17790 26086 17802 26138
rect 17854 26086 17866 26138
rect 17918 26086 22610 26138
rect 22662 26086 22674 26138
rect 22726 26086 22738 26138
rect 22790 26086 22802 26138
rect 22854 26086 22866 26138
rect 22918 26086 27610 26138
rect 27662 26086 27674 26138
rect 27726 26086 27738 26138
rect 27790 26086 27802 26138
rect 27854 26086 27866 26138
rect 27918 26086 32610 26138
rect 32662 26086 32674 26138
rect 32726 26086 32738 26138
rect 32790 26086 32802 26138
rect 32854 26086 32866 26138
rect 32918 26086 37610 26138
rect 37662 26086 37674 26138
rect 37726 26086 37738 26138
rect 37790 26086 37802 26138
rect 37854 26086 37866 26138
rect 37918 26086 40848 26138
rect 1104 26064 40848 26086
rect 32401 26027 32459 26033
rect 32401 25993 32413 26027
rect 32447 26024 32459 26027
rect 36630 26024 36636 26036
rect 32447 25996 36636 26024
rect 32447 25993 32459 25996
rect 32401 25987 32459 25993
rect 36630 25984 36636 25996
rect 36688 25984 36694 26036
rect 31846 25916 31852 25968
rect 31904 25956 31910 25968
rect 32284 25959 32342 25965
rect 32284 25956 32296 25959
rect 31904 25928 32296 25956
rect 31904 25916 31910 25928
rect 32284 25925 32296 25928
rect 32330 25925 32342 25959
rect 32284 25919 32342 25925
rect 32769 25891 32827 25897
rect 32769 25857 32781 25891
rect 32815 25888 32827 25891
rect 32950 25888 32956 25900
rect 32815 25860 32956 25888
rect 32815 25857 32827 25860
rect 32769 25851 32827 25857
rect 32950 25848 32956 25860
rect 33008 25848 33014 25900
rect 32493 25823 32551 25829
rect 32493 25789 32505 25823
rect 32539 25820 32551 25823
rect 33042 25820 33048 25832
rect 32539 25792 33048 25820
rect 32539 25789 32551 25792
rect 32493 25783 32551 25789
rect 33042 25780 33048 25792
rect 33100 25780 33106 25832
rect 32125 25755 32183 25761
rect 32125 25721 32137 25755
rect 32171 25752 32183 25755
rect 32306 25752 32312 25764
rect 32171 25724 32312 25752
rect 32171 25721 32183 25724
rect 32125 25715 32183 25721
rect 32306 25712 32312 25724
rect 32364 25712 32370 25764
rect 1104 25594 40848 25616
rect 1104 25542 1950 25594
rect 2002 25542 2014 25594
rect 2066 25542 2078 25594
rect 2130 25542 2142 25594
rect 2194 25542 2206 25594
rect 2258 25542 6950 25594
rect 7002 25542 7014 25594
rect 7066 25542 7078 25594
rect 7130 25542 7142 25594
rect 7194 25542 7206 25594
rect 7258 25542 11950 25594
rect 12002 25542 12014 25594
rect 12066 25542 12078 25594
rect 12130 25542 12142 25594
rect 12194 25542 12206 25594
rect 12258 25542 16950 25594
rect 17002 25542 17014 25594
rect 17066 25542 17078 25594
rect 17130 25542 17142 25594
rect 17194 25542 17206 25594
rect 17258 25542 21950 25594
rect 22002 25542 22014 25594
rect 22066 25542 22078 25594
rect 22130 25542 22142 25594
rect 22194 25542 22206 25594
rect 22258 25542 26950 25594
rect 27002 25542 27014 25594
rect 27066 25542 27078 25594
rect 27130 25542 27142 25594
rect 27194 25542 27206 25594
rect 27258 25542 31950 25594
rect 32002 25542 32014 25594
rect 32066 25542 32078 25594
rect 32130 25542 32142 25594
rect 32194 25542 32206 25594
rect 32258 25542 36950 25594
rect 37002 25542 37014 25594
rect 37066 25542 37078 25594
rect 37130 25542 37142 25594
rect 37194 25542 37206 25594
rect 37258 25542 40848 25594
rect 1104 25520 40848 25542
rect 9582 25440 9588 25492
rect 9640 25480 9646 25492
rect 9640 25452 22094 25480
rect 9640 25440 9646 25452
rect 11606 25304 11612 25356
rect 11664 25344 11670 25356
rect 11885 25347 11943 25353
rect 11885 25344 11897 25347
rect 11664 25316 11897 25344
rect 11664 25304 11670 25316
rect 11885 25313 11897 25316
rect 11931 25313 11943 25347
rect 11885 25307 11943 25313
rect 13909 25347 13967 25353
rect 13909 25313 13921 25347
rect 13955 25344 13967 25347
rect 14090 25344 14096 25356
rect 13955 25316 14096 25344
rect 13955 25313 13967 25316
rect 13909 25307 13967 25313
rect 14090 25304 14096 25316
rect 14148 25344 14154 25356
rect 14826 25344 14832 25356
rect 14148 25316 14832 25344
rect 14148 25304 14154 25316
rect 14826 25304 14832 25316
rect 14884 25304 14890 25356
rect 15838 25304 15844 25356
rect 15896 25344 15902 25356
rect 22066 25344 22094 25452
rect 28629 25347 28687 25353
rect 28629 25344 28641 25347
rect 15896 25316 17632 25344
rect 22066 25316 28641 25344
rect 15896 25304 15902 25316
rect 17604 25276 17632 25316
rect 28629 25313 28641 25316
rect 28675 25313 28687 25347
rect 28629 25307 28687 25313
rect 28813 25279 28871 25285
rect 28813 25276 28825 25279
rect 13294 25248 17356 25276
rect 17604 25248 28825 25276
rect 11609 25211 11667 25217
rect 11609 25177 11621 25211
rect 11655 25208 11667 25211
rect 12161 25211 12219 25217
rect 12161 25208 12173 25211
rect 11655 25180 12173 25208
rect 11655 25177 11667 25180
rect 11609 25171 11667 25177
rect 12161 25177 12173 25180
rect 12207 25208 12219 25211
rect 17328 25208 17356 25248
rect 28813 25245 28825 25248
rect 28859 25245 28871 25279
rect 29362 25276 29368 25288
rect 28813 25239 28871 25245
rect 28920 25248 29368 25276
rect 26142 25208 26148 25220
rect 12207 25180 12434 25208
rect 17328 25180 26148 25208
rect 12207 25177 12219 25180
rect 12161 25171 12219 25177
rect 12406 25140 12434 25180
rect 26142 25168 26148 25180
rect 26200 25168 26206 25220
rect 28920 25140 28948 25248
rect 29362 25236 29368 25248
rect 29420 25236 29426 25288
rect 29086 25168 29092 25220
rect 29144 25168 29150 25220
rect 12406 25112 28948 25140
rect 28994 25100 29000 25152
rect 29052 25140 29058 25152
rect 29270 25140 29276 25152
rect 29052 25112 29276 25140
rect 29052 25100 29058 25112
rect 29270 25100 29276 25112
rect 29328 25100 29334 25152
rect 1104 25050 40848 25072
rect 1104 24998 2610 25050
rect 2662 24998 2674 25050
rect 2726 24998 2738 25050
rect 2790 24998 2802 25050
rect 2854 24998 2866 25050
rect 2918 24998 7610 25050
rect 7662 24998 7674 25050
rect 7726 24998 7738 25050
rect 7790 24998 7802 25050
rect 7854 24998 7866 25050
rect 7918 24998 12610 25050
rect 12662 24998 12674 25050
rect 12726 24998 12738 25050
rect 12790 24998 12802 25050
rect 12854 24998 12866 25050
rect 12918 24998 17610 25050
rect 17662 24998 17674 25050
rect 17726 24998 17738 25050
rect 17790 24998 17802 25050
rect 17854 24998 17866 25050
rect 17918 24998 22610 25050
rect 22662 24998 22674 25050
rect 22726 24998 22738 25050
rect 22790 24998 22802 25050
rect 22854 24998 22866 25050
rect 22918 24998 27610 25050
rect 27662 24998 27674 25050
rect 27726 24998 27738 25050
rect 27790 24998 27802 25050
rect 27854 24998 27866 25050
rect 27918 24998 32610 25050
rect 32662 24998 32674 25050
rect 32726 24998 32738 25050
rect 32790 24998 32802 25050
rect 32854 24998 32866 25050
rect 32918 24998 37610 25050
rect 37662 24998 37674 25050
rect 37726 24998 37738 25050
rect 37790 24998 37802 25050
rect 37854 24998 37866 25050
rect 37918 24998 40848 25050
rect 1104 24976 40848 24998
rect 24210 24828 24216 24880
rect 24268 24828 24274 24880
rect 5718 24760 5724 24812
rect 5776 24800 5782 24812
rect 6730 24800 6736 24812
rect 5776 24772 6736 24800
rect 5776 24760 5782 24772
rect 6730 24760 6736 24772
rect 6788 24760 6794 24812
rect 18138 24760 18144 24812
rect 18196 24800 18202 24812
rect 23474 24800 23480 24812
rect 18196 24772 23480 24800
rect 18196 24760 18202 24772
rect 23474 24760 23480 24772
rect 23532 24760 23538 24812
rect 23014 24692 23020 24744
rect 23072 24732 23078 24744
rect 23753 24735 23811 24741
rect 23753 24732 23765 24735
rect 23072 24704 23765 24732
rect 23072 24692 23078 24704
rect 23753 24701 23765 24704
rect 23799 24701 23811 24735
rect 23753 24695 23811 24701
rect 25501 24735 25559 24741
rect 25501 24701 25513 24735
rect 25547 24732 25559 24735
rect 31202 24732 31208 24744
rect 25547 24704 31208 24732
rect 25547 24701 25559 24704
rect 25501 24695 25559 24701
rect 6730 24556 6736 24608
rect 6788 24596 6794 24608
rect 25516 24596 25544 24695
rect 31202 24692 31208 24704
rect 31260 24692 31266 24744
rect 6788 24568 25544 24596
rect 6788 24556 6794 24568
rect 1104 24506 40848 24528
rect 1104 24454 1950 24506
rect 2002 24454 2014 24506
rect 2066 24454 2078 24506
rect 2130 24454 2142 24506
rect 2194 24454 2206 24506
rect 2258 24454 6950 24506
rect 7002 24454 7014 24506
rect 7066 24454 7078 24506
rect 7130 24454 7142 24506
rect 7194 24454 7206 24506
rect 7258 24454 11950 24506
rect 12002 24454 12014 24506
rect 12066 24454 12078 24506
rect 12130 24454 12142 24506
rect 12194 24454 12206 24506
rect 12258 24454 16950 24506
rect 17002 24454 17014 24506
rect 17066 24454 17078 24506
rect 17130 24454 17142 24506
rect 17194 24454 17206 24506
rect 17258 24454 21950 24506
rect 22002 24454 22014 24506
rect 22066 24454 22078 24506
rect 22130 24454 22142 24506
rect 22194 24454 22206 24506
rect 22258 24454 26950 24506
rect 27002 24454 27014 24506
rect 27066 24454 27078 24506
rect 27130 24454 27142 24506
rect 27194 24454 27206 24506
rect 27258 24454 31950 24506
rect 32002 24454 32014 24506
rect 32066 24454 32078 24506
rect 32130 24454 32142 24506
rect 32194 24454 32206 24506
rect 32258 24454 36950 24506
rect 37002 24454 37014 24506
rect 37066 24454 37078 24506
rect 37130 24454 37142 24506
rect 37194 24454 37206 24506
rect 37258 24454 40848 24506
rect 1104 24432 40848 24454
rect 15562 24352 15568 24404
rect 15620 24392 15626 24404
rect 24210 24392 24216 24404
rect 15620 24364 24216 24392
rect 15620 24352 15626 24364
rect 24210 24352 24216 24364
rect 24268 24352 24274 24404
rect 27338 24284 27344 24336
rect 27396 24324 27402 24336
rect 34977 24327 35035 24333
rect 34977 24324 34989 24327
rect 27396 24296 34989 24324
rect 27396 24284 27402 24296
rect 34977 24293 34989 24296
rect 35023 24293 35035 24327
rect 34977 24287 35035 24293
rect 24118 24216 24124 24268
rect 24176 24256 24182 24268
rect 35713 24259 35771 24265
rect 35713 24256 35725 24259
rect 24176 24228 35725 24256
rect 24176 24216 24182 24228
rect 35713 24225 35725 24228
rect 35759 24225 35771 24259
rect 35713 24219 35771 24225
rect 3418 24148 3424 24200
rect 3476 24188 3482 24200
rect 3476 24160 26234 24188
rect 3476 24148 3482 24160
rect 14274 24080 14280 24132
rect 14332 24120 14338 24132
rect 14550 24120 14556 24132
rect 14332 24092 14556 24120
rect 14332 24080 14338 24092
rect 14550 24080 14556 24092
rect 14608 24080 14614 24132
rect 26206 24120 26234 24160
rect 34882 24148 34888 24200
rect 34940 24148 34946 24200
rect 35437 24191 35495 24197
rect 35437 24157 35449 24191
rect 35483 24157 35495 24191
rect 35437 24151 35495 24157
rect 35452 24120 35480 24151
rect 26206 24092 35480 24120
rect 1104 23962 40848 23984
rect 1104 23910 2610 23962
rect 2662 23910 2674 23962
rect 2726 23910 2738 23962
rect 2790 23910 2802 23962
rect 2854 23910 2866 23962
rect 2918 23910 7610 23962
rect 7662 23910 7674 23962
rect 7726 23910 7738 23962
rect 7790 23910 7802 23962
rect 7854 23910 7866 23962
rect 7918 23910 12610 23962
rect 12662 23910 12674 23962
rect 12726 23910 12738 23962
rect 12790 23910 12802 23962
rect 12854 23910 12866 23962
rect 12918 23910 17610 23962
rect 17662 23910 17674 23962
rect 17726 23910 17738 23962
rect 17790 23910 17802 23962
rect 17854 23910 17866 23962
rect 17918 23910 22610 23962
rect 22662 23910 22674 23962
rect 22726 23910 22738 23962
rect 22790 23910 22802 23962
rect 22854 23910 22866 23962
rect 22918 23910 27610 23962
rect 27662 23910 27674 23962
rect 27726 23910 27738 23962
rect 27790 23910 27802 23962
rect 27854 23910 27866 23962
rect 27918 23910 32610 23962
rect 32662 23910 32674 23962
rect 32726 23910 32738 23962
rect 32790 23910 32802 23962
rect 32854 23910 32866 23962
rect 32918 23910 37610 23962
rect 37662 23910 37674 23962
rect 37726 23910 37738 23962
rect 37790 23910 37802 23962
rect 37854 23910 37866 23962
rect 37918 23910 40848 23962
rect 1104 23888 40848 23910
rect 26206 23820 33640 23848
rect 9674 23740 9680 23792
rect 9732 23780 9738 23792
rect 26206 23780 26234 23820
rect 9732 23752 26234 23780
rect 9732 23740 9738 23752
rect 33226 23740 33232 23792
rect 33284 23780 33290 23792
rect 33612 23789 33640 23820
rect 33413 23783 33471 23789
rect 33413 23780 33425 23783
rect 33284 23752 33425 23780
rect 33284 23740 33290 23752
rect 33413 23749 33425 23752
rect 33459 23749 33471 23783
rect 33413 23743 33471 23749
rect 33597 23783 33655 23789
rect 33597 23749 33609 23783
rect 33643 23780 33655 23783
rect 33873 23783 33931 23789
rect 33873 23780 33885 23783
rect 33643 23752 33885 23780
rect 33643 23749 33655 23752
rect 33597 23743 33655 23749
rect 33873 23749 33885 23752
rect 33919 23749 33931 23783
rect 33873 23743 33931 23749
rect 21726 23672 21732 23724
rect 21784 23712 21790 23724
rect 22005 23715 22063 23721
rect 22005 23712 22017 23715
rect 21784 23684 22017 23712
rect 21784 23672 21790 23684
rect 22005 23681 22017 23684
rect 22051 23681 22063 23715
rect 22005 23675 22063 23681
rect 2314 23536 2320 23588
rect 2372 23576 2378 23588
rect 33229 23579 33287 23585
rect 33229 23576 33241 23579
rect 2372 23548 33241 23576
rect 2372 23536 2378 23548
rect 33229 23545 33241 23548
rect 33275 23545 33287 23579
rect 33229 23539 33287 23545
rect 21818 23468 21824 23520
rect 21876 23508 21882 23520
rect 21913 23511 21971 23517
rect 21913 23508 21925 23511
rect 21876 23480 21925 23508
rect 21876 23468 21882 23480
rect 21913 23477 21925 23480
rect 21959 23477 21971 23511
rect 21913 23471 21971 23477
rect 32861 23511 32919 23517
rect 32861 23477 32873 23511
rect 32907 23508 32919 23511
rect 33410 23508 33416 23520
rect 32907 23480 33416 23508
rect 32907 23477 32919 23480
rect 32861 23471 32919 23477
rect 33410 23468 33416 23480
rect 33468 23468 33474 23520
rect 1104 23418 40848 23440
rect 1104 23366 1950 23418
rect 2002 23366 2014 23418
rect 2066 23366 2078 23418
rect 2130 23366 2142 23418
rect 2194 23366 2206 23418
rect 2258 23366 6950 23418
rect 7002 23366 7014 23418
rect 7066 23366 7078 23418
rect 7130 23366 7142 23418
rect 7194 23366 7206 23418
rect 7258 23366 11950 23418
rect 12002 23366 12014 23418
rect 12066 23366 12078 23418
rect 12130 23366 12142 23418
rect 12194 23366 12206 23418
rect 12258 23366 16950 23418
rect 17002 23366 17014 23418
rect 17066 23366 17078 23418
rect 17130 23366 17142 23418
rect 17194 23366 17206 23418
rect 17258 23366 21950 23418
rect 22002 23366 22014 23418
rect 22066 23366 22078 23418
rect 22130 23366 22142 23418
rect 22194 23366 22206 23418
rect 22258 23366 26950 23418
rect 27002 23366 27014 23418
rect 27066 23366 27078 23418
rect 27130 23366 27142 23418
rect 27194 23366 27206 23418
rect 27258 23366 31950 23418
rect 32002 23366 32014 23418
rect 32066 23366 32078 23418
rect 32130 23366 32142 23418
rect 32194 23366 32206 23418
rect 32258 23366 36950 23418
rect 37002 23366 37014 23418
rect 37066 23366 37078 23418
rect 37130 23366 37142 23418
rect 37194 23366 37206 23418
rect 37258 23366 40848 23418
rect 1104 23344 40848 23366
rect 10321 23239 10379 23245
rect 10321 23205 10333 23239
rect 10367 23236 10379 23239
rect 19610 23236 19616 23248
rect 10367 23208 19616 23236
rect 10367 23205 10379 23208
rect 10321 23199 10379 23205
rect 19610 23196 19616 23208
rect 19668 23196 19674 23248
rect 10229 23103 10287 23109
rect 10229 23069 10241 23103
rect 10275 23100 10287 23103
rect 10318 23100 10324 23112
rect 10275 23072 10324 23100
rect 10275 23069 10287 23072
rect 10229 23063 10287 23069
rect 10318 23060 10324 23072
rect 10376 23060 10382 23112
rect 14182 23060 14188 23112
rect 14240 23100 14246 23112
rect 16482 23100 16488 23112
rect 14240 23072 16488 23100
rect 14240 23060 14246 23072
rect 16482 23060 16488 23072
rect 16540 23060 16546 23112
rect 3234 22992 3240 23044
rect 3292 23032 3298 23044
rect 25038 23032 25044 23044
rect 3292 23004 25044 23032
rect 3292 22992 3298 23004
rect 25038 22992 25044 23004
rect 25096 22992 25102 23044
rect 5626 22924 5632 22976
rect 5684 22964 5690 22976
rect 9858 22964 9864 22976
rect 5684 22936 9864 22964
rect 5684 22924 5690 22936
rect 9858 22924 9864 22936
rect 9916 22924 9922 22976
rect 16577 22967 16635 22973
rect 16577 22933 16589 22967
rect 16623 22964 16635 22967
rect 38654 22964 38660 22976
rect 16623 22936 38660 22964
rect 16623 22933 16635 22936
rect 16577 22927 16635 22933
rect 38654 22924 38660 22936
rect 38712 22924 38718 22976
rect 1104 22874 40848 22896
rect 1104 22822 2610 22874
rect 2662 22822 2674 22874
rect 2726 22822 2738 22874
rect 2790 22822 2802 22874
rect 2854 22822 2866 22874
rect 2918 22822 7610 22874
rect 7662 22822 7674 22874
rect 7726 22822 7738 22874
rect 7790 22822 7802 22874
rect 7854 22822 7866 22874
rect 7918 22822 12610 22874
rect 12662 22822 12674 22874
rect 12726 22822 12738 22874
rect 12790 22822 12802 22874
rect 12854 22822 12866 22874
rect 12918 22822 17610 22874
rect 17662 22822 17674 22874
rect 17726 22822 17738 22874
rect 17790 22822 17802 22874
rect 17854 22822 17866 22874
rect 17918 22822 22610 22874
rect 22662 22822 22674 22874
rect 22726 22822 22738 22874
rect 22790 22822 22802 22874
rect 22854 22822 22866 22874
rect 22918 22822 27610 22874
rect 27662 22822 27674 22874
rect 27726 22822 27738 22874
rect 27790 22822 27802 22874
rect 27854 22822 27866 22874
rect 27918 22822 32610 22874
rect 32662 22822 32674 22874
rect 32726 22822 32738 22874
rect 32790 22822 32802 22874
rect 32854 22822 32866 22874
rect 32918 22822 37610 22874
rect 37662 22822 37674 22874
rect 37726 22822 37738 22874
rect 37790 22822 37802 22874
rect 37854 22822 37866 22874
rect 37918 22822 40848 22874
rect 1104 22800 40848 22822
rect 3234 22720 3240 22772
rect 3292 22720 3298 22772
rect 6822 22760 6828 22772
rect 6748 22732 6828 22760
rect 6748 22701 6776 22732
rect 6822 22720 6828 22732
rect 6880 22720 6886 22772
rect 6914 22720 6920 22772
rect 6972 22760 6978 22772
rect 19334 22760 19340 22772
rect 6972 22732 19340 22760
rect 6972 22720 6978 22732
rect 19334 22720 19340 22732
rect 19392 22720 19398 22772
rect 6725 22695 6783 22701
rect 6725 22661 6737 22695
rect 6771 22661 6783 22695
rect 6725 22655 6783 22661
rect 7101 22695 7159 22701
rect 7101 22661 7113 22695
rect 7147 22692 7159 22695
rect 7282 22692 7288 22704
rect 7147 22664 7288 22692
rect 7147 22661 7159 22664
rect 7101 22655 7159 22661
rect 7282 22652 7288 22664
rect 7340 22652 7346 22704
rect 24578 22652 24584 22704
rect 24636 22652 24642 22704
rect 3234 22584 3240 22636
rect 3292 22584 3298 22636
rect 3510 22584 3516 22636
rect 3568 22584 3574 22636
rect 6549 22627 6607 22633
rect 6549 22624 6561 22627
rect 6288 22596 6561 22624
rect 3053 22559 3111 22565
rect 3053 22525 3065 22559
rect 3099 22556 3111 22559
rect 5626 22556 5632 22568
rect 3099 22528 5632 22556
rect 3099 22525 3111 22528
rect 3053 22519 3111 22525
rect 5626 22516 5632 22528
rect 5684 22516 5690 22568
rect 6178 22448 6184 22500
rect 6236 22488 6242 22500
rect 6288 22488 6316 22596
rect 6549 22593 6561 22596
rect 6595 22593 6607 22627
rect 6549 22587 6607 22593
rect 6641 22627 6699 22633
rect 6641 22593 6653 22627
rect 6687 22624 6699 22627
rect 8294 22624 8300 22636
rect 6687 22596 8300 22624
rect 6687 22593 6699 22596
rect 6641 22587 6699 22593
rect 8294 22584 8300 22596
rect 8352 22584 8358 22636
rect 6365 22559 6423 22565
rect 6365 22525 6377 22559
rect 6411 22556 6423 22559
rect 8662 22556 8668 22568
rect 6411 22528 8668 22556
rect 6411 22525 6423 22528
rect 6365 22519 6423 22525
rect 8662 22516 8668 22528
rect 8720 22516 8726 22568
rect 7469 22491 7527 22497
rect 7469 22488 7481 22491
rect 6236 22460 7481 22488
rect 6236 22448 6242 22460
rect 7469 22457 7481 22460
rect 7515 22488 7527 22491
rect 36170 22488 36176 22500
rect 7515 22460 36176 22488
rect 7515 22457 7527 22460
rect 7469 22451 7527 22457
rect 36170 22448 36176 22460
rect 36228 22448 36234 22500
rect 24670 22380 24676 22432
rect 24728 22420 24734 22432
rect 25869 22423 25927 22429
rect 25869 22420 25881 22423
rect 24728 22392 25881 22420
rect 24728 22380 24734 22392
rect 25869 22389 25881 22392
rect 25915 22389 25927 22423
rect 25869 22383 25927 22389
rect 1104 22330 40848 22352
rect 1104 22278 1950 22330
rect 2002 22278 2014 22330
rect 2066 22278 2078 22330
rect 2130 22278 2142 22330
rect 2194 22278 2206 22330
rect 2258 22278 6950 22330
rect 7002 22278 7014 22330
rect 7066 22278 7078 22330
rect 7130 22278 7142 22330
rect 7194 22278 7206 22330
rect 7258 22278 11950 22330
rect 12002 22278 12014 22330
rect 12066 22278 12078 22330
rect 12130 22278 12142 22330
rect 12194 22278 12206 22330
rect 12258 22278 16950 22330
rect 17002 22278 17014 22330
rect 17066 22278 17078 22330
rect 17130 22278 17142 22330
rect 17194 22278 17206 22330
rect 17258 22278 21950 22330
rect 22002 22278 22014 22330
rect 22066 22278 22078 22330
rect 22130 22278 22142 22330
rect 22194 22278 22206 22330
rect 22258 22278 26950 22330
rect 27002 22278 27014 22330
rect 27066 22278 27078 22330
rect 27130 22278 27142 22330
rect 27194 22278 27206 22330
rect 27258 22278 31950 22330
rect 32002 22278 32014 22330
rect 32066 22278 32078 22330
rect 32130 22278 32142 22330
rect 32194 22278 32206 22330
rect 32258 22278 36950 22330
rect 37002 22278 37014 22330
rect 37066 22278 37078 22330
rect 37130 22278 37142 22330
rect 37194 22278 37206 22330
rect 37258 22278 40848 22330
rect 1104 22256 40848 22278
rect 6914 22176 6920 22228
rect 6972 22216 6978 22228
rect 7282 22216 7288 22228
rect 6972 22188 7288 22216
rect 6972 22176 6978 22188
rect 7282 22176 7288 22188
rect 7340 22176 7346 22228
rect 9582 22176 9588 22228
rect 9640 22216 9646 22228
rect 9769 22219 9827 22225
rect 9769 22216 9781 22219
rect 9640 22188 9781 22216
rect 9640 22176 9646 22188
rect 9769 22185 9781 22188
rect 9815 22216 9827 22219
rect 11606 22216 11612 22228
rect 9815 22188 11612 22216
rect 9815 22185 9827 22188
rect 9769 22179 9827 22185
rect 11606 22176 11612 22188
rect 11664 22176 11670 22228
rect 3510 22040 3516 22092
rect 3568 22080 3574 22092
rect 7282 22080 7288 22092
rect 3568 22052 7288 22080
rect 3568 22040 3574 22052
rect 7282 22040 7288 22052
rect 7340 22080 7346 22092
rect 8386 22080 8392 22092
rect 7340 22052 8392 22080
rect 7340 22040 7346 22052
rect 8386 22040 8392 22052
rect 8444 22040 8450 22092
rect 11054 21904 11060 21956
rect 11112 21904 11118 21956
rect 23382 21904 23388 21956
rect 23440 21944 23446 21956
rect 24670 21944 24676 21956
rect 23440 21916 24676 21944
rect 23440 21904 23446 21916
rect 24670 21904 24676 21916
rect 24728 21904 24734 21956
rect 1104 21786 40848 21808
rect 1104 21734 2610 21786
rect 2662 21734 2674 21786
rect 2726 21734 2738 21786
rect 2790 21734 2802 21786
rect 2854 21734 2866 21786
rect 2918 21734 7610 21786
rect 7662 21734 7674 21786
rect 7726 21734 7738 21786
rect 7790 21734 7802 21786
rect 7854 21734 7866 21786
rect 7918 21734 12610 21786
rect 12662 21734 12674 21786
rect 12726 21734 12738 21786
rect 12790 21734 12802 21786
rect 12854 21734 12866 21786
rect 12918 21734 17610 21786
rect 17662 21734 17674 21786
rect 17726 21734 17738 21786
rect 17790 21734 17802 21786
rect 17854 21734 17866 21786
rect 17918 21734 22610 21786
rect 22662 21734 22674 21786
rect 22726 21734 22738 21786
rect 22790 21734 22802 21786
rect 22854 21734 22866 21786
rect 22918 21734 27610 21786
rect 27662 21734 27674 21786
rect 27726 21734 27738 21786
rect 27790 21734 27802 21786
rect 27854 21734 27866 21786
rect 27918 21734 32610 21786
rect 32662 21734 32674 21786
rect 32726 21734 32738 21786
rect 32790 21734 32802 21786
rect 32854 21734 32866 21786
rect 32918 21734 37610 21786
rect 37662 21734 37674 21786
rect 37726 21734 37738 21786
rect 37790 21734 37802 21786
rect 37854 21734 37866 21786
rect 37918 21734 40848 21786
rect 1104 21712 40848 21734
rect 22370 21564 22376 21616
rect 22428 21604 22434 21616
rect 22833 21607 22891 21613
rect 22833 21604 22845 21607
rect 22428 21576 22845 21604
rect 22428 21564 22434 21576
rect 22833 21573 22845 21576
rect 22879 21573 22891 21607
rect 27522 21604 27528 21616
rect 24058 21576 27528 21604
rect 22833 21567 22891 21573
rect 27522 21564 27528 21576
rect 27580 21564 27586 21616
rect 31110 21564 31116 21616
rect 31168 21604 31174 21616
rect 31662 21604 31668 21616
rect 31168 21576 31668 21604
rect 31168 21564 31174 21576
rect 31662 21564 31668 21576
rect 31720 21604 31726 21616
rect 31720 21576 32720 21604
rect 31720 21564 31726 21576
rect 22554 21496 22560 21548
rect 22612 21496 22618 21548
rect 32692 21545 32720 21576
rect 32677 21539 32735 21545
rect 32677 21505 32689 21539
rect 32723 21505 32735 21539
rect 32677 21499 32735 21505
rect 33505 21539 33563 21545
rect 33505 21505 33517 21539
rect 33551 21536 33563 21539
rect 37366 21536 37372 21548
rect 33551 21508 37372 21536
rect 33551 21505 33563 21508
rect 33505 21499 33563 21505
rect 37366 21496 37372 21508
rect 37424 21496 37430 21548
rect 24581 21471 24639 21477
rect 22066 21440 23888 21468
rect 6914 21292 6920 21344
rect 6972 21332 6978 21344
rect 22066 21332 22094 21440
rect 6972 21304 22094 21332
rect 6972 21292 6978 21304
rect 22554 21292 22560 21344
rect 22612 21332 22618 21344
rect 23382 21332 23388 21344
rect 22612 21304 23388 21332
rect 22612 21292 22618 21304
rect 23382 21292 23388 21304
rect 23440 21292 23446 21344
rect 23860 21332 23888 21440
rect 24581 21437 24593 21471
rect 24627 21468 24639 21471
rect 28994 21468 29000 21480
rect 24627 21440 29000 21468
rect 24627 21437 24639 21440
rect 24581 21431 24639 21437
rect 28994 21428 29000 21440
rect 29052 21428 29058 21480
rect 33873 21471 33931 21477
rect 31754 21360 31760 21412
rect 31812 21400 31818 21412
rect 32493 21403 32551 21409
rect 32493 21400 32505 21403
rect 31812 21372 32505 21400
rect 31812 21360 31818 21372
rect 32493 21369 32505 21372
rect 32539 21369 32551 21403
rect 32493 21363 32551 21369
rect 32398 21332 32404 21344
rect 23860 21304 32404 21332
rect 32398 21292 32404 21304
rect 32456 21332 32462 21344
rect 32600 21332 32628 21454
rect 33873 21437 33885 21471
rect 33919 21468 33931 21471
rect 36630 21468 36636 21480
rect 33919 21440 36636 21468
rect 33919 21437 33931 21440
rect 33873 21431 33931 21437
rect 36630 21428 36636 21440
rect 36688 21428 36694 21480
rect 32456 21304 32628 21332
rect 32456 21292 32462 21304
rect 1104 21242 40848 21264
rect 1104 21190 1950 21242
rect 2002 21190 2014 21242
rect 2066 21190 2078 21242
rect 2130 21190 2142 21242
rect 2194 21190 2206 21242
rect 2258 21190 6950 21242
rect 7002 21190 7014 21242
rect 7066 21190 7078 21242
rect 7130 21190 7142 21242
rect 7194 21190 7206 21242
rect 7258 21190 11950 21242
rect 12002 21190 12014 21242
rect 12066 21190 12078 21242
rect 12130 21190 12142 21242
rect 12194 21190 12206 21242
rect 12258 21190 16950 21242
rect 17002 21190 17014 21242
rect 17066 21190 17078 21242
rect 17130 21190 17142 21242
rect 17194 21190 17206 21242
rect 17258 21190 21950 21242
rect 22002 21190 22014 21242
rect 22066 21190 22078 21242
rect 22130 21190 22142 21242
rect 22194 21190 22206 21242
rect 22258 21190 26950 21242
rect 27002 21190 27014 21242
rect 27066 21190 27078 21242
rect 27130 21190 27142 21242
rect 27194 21190 27206 21242
rect 27258 21190 31950 21242
rect 32002 21190 32014 21242
rect 32066 21190 32078 21242
rect 32130 21190 32142 21242
rect 32194 21190 32206 21242
rect 32258 21190 36950 21242
rect 37002 21190 37014 21242
rect 37066 21190 37078 21242
rect 37130 21190 37142 21242
rect 37194 21190 37206 21242
rect 37258 21190 40848 21242
rect 1104 21168 40848 21190
rect 1104 20698 40848 20720
rect 1104 20646 2610 20698
rect 2662 20646 2674 20698
rect 2726 20646 2738 20698
rect 2790 20646 2802 20698
rect 2854 20646 2866 20698
rect 2918 20646 7610 20698
rect 7662 20646 7674 20698
rect 7726 20646 7738 20698
rect 7790 20646 7802 20698
rect 7854 20646 7866 20698
rect 7918 20646 12610 20698
rect 12662 20646 12674 20698
rect 12726 20646 12738 20698
rect 12790 20646 12802 20698
rect 12854 20646 12866 20698
rect 12918 20646 17610 20698
rect 17662 20646 17674 20698
rect 17726 20646 17738 20698
rect 17790 20646 17802 20698
rect 17854 20646 17866 20698
rect 17918 20646 22610 20698
rect 22662 20646 22674 20698
rect 22726 20646 22738 20698
rect 22790 20646 22802 20698
rect 22854 20646 22866 20698
rect 22918 20646 27610 20698
rect 27662 20646 27674 20698
rect 27726 20646 27738 20698
rect 27790 20646 27802 20698
rect 27854 20646 27866 20698
rect 27918 20646 32610 20698
rect 32662 20646 32674 20698
rect 32726 20646 32738 20698
rect 32790 20646 32802 20698
rect 32854 20646 32866 20698
rect 32918 20646 37610 20698
rect 37662 20646 37674 20698
rect 37726 20646 37738 20698
rect 37790 20646 37802 20698
rect 37854 20646 37866 20698
rect 37918 20646 40848 20698
rect 1104 20624 40848 20646
rect 2685 20587 2743 20593
rect 2685 20553 2697 20587
rect 2731 20584 2743 20587
rect 2731 20556 4384 20584
rect 2731 20553 2743 20556
rect 2685 20547 2743 20553
rect 2961 20519 3019 20525
rect 2961 20485 2973 20519
rect 3007 20516 3019 20519
rect 3418 20516 3424 20528
rect 3007 20488 3424 20516
rect 3007 20485 3019 20488
rect 2961 20479 3019 20485
rect 3418 20476 3424 20488
rect 3476 20476 3482 20528
rect 4356 20516 4384 20556
rect 40402 20516 40408 20528
rect 4278 20488 40408 20516
rect 40402 20476 40408 20488
rect 40460 20476 40466 20528
rect 4709 20383 4767 20389
rect 4709 20349 4721 20383
rect 4755 20380 4767 20383
rect 4985 20383 5043 20389
rect 4755 20352 4936 20380
rect 4755 20349 4767 20352
rect 4709 20343 4767 20349
rect 4908 20244 4936 20352
rect 4985 20349 4997 20383
rect 5031 20380 5043 20383
rect 6638 20380 6644 20392
rect 5031 20352 6644 20380
rect 5031 20349 5043 20352
rect 4985 20343 5043 20349
rect 6638 20340 6644 20352
rect 6696 20340 6702 20392
rect 5353 20247 5411 20253
rect 5353 20244 5365 20247
rect 4908 20216 5365 20244
rect 5353 20213 5365 20216
rect 5399 20244 5411 20247
rect 39574 20244 39580 20256
rect 5399 20216 39580 20244
rect 5399 20213 5411 20216
rect 5353 20207 5411 20213
rect 39574 20204 39580 20216
rect 39632 20204 39638 20256
rect 1104 20154 40848 20176
rect 1104 20102 1950 20154
rect 2002 20102 2014 20154
rect 2066 20102 2078 20154
rect 2130 20102 2142 20154
rect 2194 20102 2206 20154
rect 2258 20102 6950 20154
rect 7002 20102 7014 20154
rect 7066 20102 7078 20154
rect 7130 20102 7142 20154
rect 7194 20102 7206 20154
rect 7258 20102 11950 20154
rect 12002 20102 12014 20154
rect 12066 20102 12078 20154
rect 12130 20102 12142 20154
rect 12194 20102 12206 20154
rect 12258 20102 16950 20154
rect 17002 20102 17014 20154
rect 17066 20102 17078 20154
rect 17130 20102 17142 20154
rect 17194 20102 17206 20154
rect 17258 20102 21950 20154
rect 22002 20102 22014 20154
rect 22066 20102 22078 20154
rect 22130 20102 22142 20154
rect 22194 20102 22206 20154
rect 22258 20102 26950 20154
rect 27002 20102 27014 20154
rect 27066 20102 27078 20154
rect 27130 20102 27142 20154
rect 27194 20102 27206 20154
rect 27258 20102 31950 20154
rect 32002 20102 32014 20154
rect 32066 20102 32078 20154
rect 32130 20102 32142 20154
rect 32194 20102 32206 20154
rect 32258 20102 36950 20154
rect 37002 20102 37014 20154
rect 37066 20102 37078 20154
rect 37130 20102 37142 20154
rect 37194 20102 37206 20154
rect 37258 20102 40848 20154
rect 1104 20080 40848 20102
rect 22005 20043 22063 20049
rect 22005 20009 22017 20043
rect 22051 20040 22063 20043
rect 23014 20040 23020 20052
rect 22051 20012 23020 20040
rect 22051 20009 22063 20012
rect 22005 20003 22063 20009
rect 23014 20000 23020 20012
rect 23072 20000 23078 20052
rect 19245 19907 19303 19913
rect 19245 19873 19257 19907
rect 19291 19904 19303 19907
rect 19426 19904 19432 19916
rect 19291 19876 19432 19904
rect 19291 19873 19303 19876
rect 19245 19867 19303 19873
rect 19426 19864 19432 19876
rect 19484 19864 19490 19916
rect 20990 19864 20996 19916
rect 21048 19864 21054 19916
rect 21269 19907 21327 19913
rect 21269 19873 21281 19907
rect 21315 19904 21327 19907
rect 23382 19904 23388 19916
rect 21315 19876 23388 19904
rect 21315 19873 21327 19876
rect 21269 19867 21327 19873
rect 23382 19864 23388 19876
rect 23440 19864 23446 19916
rect 8202 19796 8208 19848
rect 8260 19836 8266 19848
rect 21821 19839 21879 19845
rect 8260 19808 19918 19836
rect 8260 19796 8266 19808
rect 21821 19805 21833 19839
rect 21867 19836 21879 19839
rect 24394 19836 24400 19848
rect 21867 19808 24400 19836
rect 21867 19805 21879 19808
rect 21821 19799 21879 19805
rect 24394 19796 24400 19808
rect 24452 19796 24458 19848
rect 1104 19610 40848 19632
rect 1104 19558 2610 19610
rect 2662 19558 2674 19610
rect 2726 19558 2738 19610
rect 2790 19558 2802 19610
rect 2854 19558 2866 19610
rect 2918 19558 7610 19610
rect 7662 19558 7674 19610
rect 7726 19558 7738 19610
rect 7790 19558 7802 19610
rect 7854 19558 7866 19610
rect 7918 19558 12610 19610
rect 12662 19558 12674 19610
rect 12726 19558 12738 19610
rect 12790 19558 12802 19610
rect 12854 19558 12866 19610
rect 12918 19558 17610 19610
rect 17662 19558 17674 19610
rect 17726 19558 17738 19610
rect 17790 19558 17802 19610
rect 17854 19558 17866 19610
rect 17918 19558 22610 19610
rect 22662 19558 22674 19610
rect 22726 19558 22738 19610
rect 22790 19558 22802 19610
rect 22854 19558 22866 19610
rect 22918 19558 27610 19610
rect 27662 19558 27674 19610
rect 27726 19558 27738 19610
rect 27790 19558 27802 19610
rect 27854 19558 27866 19610
rect 27918 19558 32610 19610
rect 32662 19558 32674 19610
rect 32726 19558 32738 19610
rect 32790 19558 32802 19610
rect 32854 19558 32866 19610
rect 32918 19558 37610 19610
rect 37662 19558 37674 19610
rect 37726 19558 37738 19610
rect 37790 19558 37802 19610
rect 37854 19558 37866 19610
rect 37918 19558 40848 19610
rect 1104 19536 40848 19558
rect 6638 19456 6644 19508
rect 6696 19496 6702 19508
rect 9582 19496 9588 19508
rect 6696 19468 9588 19496
rect 6696 19456 6702 19468
rect 9582 19456 9588 19468
rect 9640 19456 9646 19508
rect 30834 19428 30840 19440
rect 8142 19400 30840 19428
rect 30834 19388 30840 19400
rect 30892 19388 30898 19440
rect 6638 19320 6644 19372
rect 6696 19320 6702 19372
rect 8662 19320 8668 19372
rect 8720 19320 8726 19372
rect 1854 19252 1860 19304
rect 1912 19292 1918 19304
rect 6917 19295 6975 19301
rect 6917 19292 6929 19295
rect 1912 19264 6929 19292
rect 1912 19252 1918 19264
rect 6917 19261 6929 19264
rect 6963 19261 6975 19295
rect 6917 19255 6975 19261
rect 1104 19066 40848 19088
rect 1104 19014 1950 19066
rect 2002 19014 2014 19066
rect 2066 19014 2078 19066
rect 2130 19014 2142 19066
rect 2194 19014 2206 19066
rect 2258 19014 6950 19066
rect 7002 19014 7014 19066
rect 7066 19014 7078 19066
rect 7130 19014 7142 19066
rect 7194 19014 7206 19066
rect 7258 19014 11950 19066
rect 12002 19014 12014 19066
rect 12066 19014 12078 19066
rect 12130 19014 12142 19066
rect 12194 19014 12206 19066
rect 12258 19014 16950 19066
rect 17002 19014 17014 19066
rect 17066 19014 17078 19066
rect 17130 19014 17142 19066
rect 17194 19014 17206 19066
rect 17258 19014 21950 19066
rect 22002 19014 22014 19066
rect 22066 19014 22078 19066
rect 22130 19014 22142 19066
rect 22194 19014 22206 19066
rect 22258 19014 26950 19066
rect 27002 19014 27014 19066
rect 27066 19014 27078 19066
rect 27130 19014 27142 19066
rect 27194 19014 27206 19066
rect 27258 19014 31950 19066
rect 32002 19014 32014 19066
rect 32066 19014 32078 19066
rect 32130 19014 32142 19066
rect 32194 19014 32206 19066
rect 32258 19014 36950 19066
rect 37002 19014 37014 19066
rect 37066 19014 37078 19066
rect 37130 19014 37142 19066
rect 37194 19014 37206 19066
rect 37258 19014 40848 19066
rect 1104 18992 40848 19014
rect 6886 18856 9720 18884
rect 6886 18816 6914 18856
rect 3436 18788 6914 18816
rect 3436 18757 3464 18788
rect 9582 18776 9588 18828
rect 9640 18776 9646 18828
rect 9692 18816 9720 18856
rect 25958 18816 25964 18828
rect 9692 18788 25964 18816
rect 25958 18776 25964 18788
rect 26016 18776 26022 18828
rect 3145 18751 3203 18757
rect 3145 18717 3157 18751
rect 3191 18748 3203 18751
rect 3421 18751 3479 18757
rect 3421 18748 3433 18751
rect 3191 18720 3433 18748
rect 3191 18717 3203 18720
rect 3145 18711 3203 18717
rect 3421 18717 3433 18720
rect 3467 18717 3479 18751
rect 10994 18734 22094 18748
rect 3421 18711 3479 18717
rect 10980 18720 22094 18734
rect 9858 18640 9864 18692
rect 9916 18640 9922 18692
rect 3602 18572 3608 18624
rect 3660 18572 3666 18624
rect 9309 18615 9367 18621
rect 9309 18581 9321 18615
rect 9355 18612 9367 18615
rect 10980 18612 11008 18720
rect 11609 18683 11667 18689
rect 11609 18649 11621 18683
rect 11655 18680 11667 18683
rect 17310 18680 17316 18692
rect 11655 18652 17316 18680
rect 11655 18649 11667 18652
rect 11609 18643 11667 18649
rect 17310 18640 17316 18652
rect 17368 18640 17374 18692
rect 22066 18680 22094 18720
rect 39850 18680 39856 18692
rect 22066 18652 39856 18680
rect 39850 18640 39856 18652
rect 39908 18640 39914 18692
rect 9355 18584 11008 18612
rect 9355 18581 9367 18584
rect 9309 18575 9367 18581
rect 1104 18522 40848 18544
rect 1104 18470 2610 18522
rect 2662 18470 2674 18522
rect 2726 18470 2738 18522
rect 2790 18470 2802 18522
rect 2854 18470 2866 18522
rect 2918 18470 7610 18522
rect 7662 18470 7674 18522
rect 7726 18470 7738 18522
rect 7790 18470 7802 18522
rect 7854 18470 7866 18522
rect 7918 18470 12610 18522
rect 12662 18470 12674 18522
rect 12726 18470 12738 18522
rect 12790 18470 12802 18522
rect 12854 18470 12866 18522
rect 12918 18470 17610 18522
rect 17662 18470 17674 18522
rect 17726 18470 17738 18522
rect 17790 18470 17802 18522
rect 17854 18470 17866 18522
rect 17918 18470 22610 18522
rect 22662 18470 22674 18522
rect 22726 18470 22738 18522
rect 22790 18470 22802 18522
rect 22854 18470 22866 18522
rect 22918 18470 27610 18522
rect 27662 18470 27674 18522
rect 27726 18470 27738 18522
rect 27790 18470 27802 18522
rect 27854 18470 27866 18522
rect 27918 18470 32610 18522
rect 32662 18470 32674 18522
rect 32726 18470 32738 18522
rect 32790 18470 32802 18522
rect 32854 18470 32866 18522
rect 32918 18470 37610 18522
rect 37662 18470 37674 18522
rect 37726 18470 37738 18522
rect 37790 18470 37802 18522
rect 37854 18470 37866 18522
rect 37918 18470 40848 18522
rect 1104 18448 40848 18470
rect 3602 18368 3608 18420
rect 3660 18408 3666 18420
rect 9858 18408 9864 18420
rect 3660 18380 9864 18408
rect 3660 18368 3666 18380
rect 9858 18368 9864 18380
rect 9916 18368 9922 18420
rect 36630 18368 36636 18420
rect 36688 18368 36694 18420
rect 33410 18300 33416 18352
rect 33468 18340 33474 18352
rect 36449 18343 36507 18349
rect 36449 18340 36461 18343
rect 33468 18312 36461 18340
rect 33468 18300 33474 18312
rect 36449 18309 36461 18312
rect 36495 18309 36507 18343
rect 36449 18303 36507 18309
rect 36909 18275 36967 18281
rect 36909 18272 36921 18275
rect 31726 18244 36921 18272
rect 24118 18164 24124 18216
rect 24176 18204 24182 18216
rect 31726 18204 31754 18244
rect 36909 18241 36921 18244
rect 36955 18241 36967 18275
rect 36909 18235 36967 18241
rect 24176 18176 31754 18204
rect 24176 18164 24182 18176
rect 9214 18096 9220 18148
rect 9272 18136 9278 18148
rect 26786 18136 26792 18148
rect 9272 18108 26792 18136
rect 9272 18096 9278 18108
rect 26786 18096 26792 18108
rect 26844 18096 26850 18148
rect 26970 18096 26976 18148
rect 27028 18136 27034 18148
rect 27028 18108 36032 18136
rect 27028 18096 27034 18108
rect 1670 18028 1676 18080
rect 1728 18068 1734 18080
rect 24118 18068 24124 18080
rect 1728 18040 24124 18068
rect 1728 18028 1734 18040
rect 24118 18028 24124 18040
rect 24176 18028 24182 18080
rect 36004 18068 36032 18108
rect 36173 18071 36231 18077
rect 36173 18068 36185 18071
rect 36004 18040 36185 18068
rect 36173 18037 36185 18040
rect 36219 18068 36231 18071
rect 36633 18071 36691 18077
rect 36633 18068 36645 18071
rect 36219 18040 36645 18068
rect 36219 18037 36231 18040
rect 36173 18031 36231 18037
rect 36633 18037 36645 18040
rect 36679 18037 36691 18071
rect 36633 18031 36691 18037
rect 1104 17978 40848 18000
rect 1104 17926 1950 17978
rect 2002 17926 2014 17978
rect 2066 17926 2078 17978
rect 2130 17926 2142 17978
rect 2194 17926 2206 17978
rect 2258 17926 6950 17978
rect 7002 17926 7014 17978
rect 7066 17926 7078 17978
rect 7130 17926 7142 17978
rect 7194 17926 7206 17978
rect 7258 17926 11950 17978
rect 12002 17926 12014 17978
rect 12066 17926 12078 17978
rect 12130 17926 12142 17978
rect 12194 17926 12206 17978
rect 12258 17926 16950 17978
rect 17002 17926 17014 17978
rect 17066 17926 17078 17978
rect 17130 17926 17142 17978
rect 17194 17926 17206 17978
rect 17258 17926 21950 17978
rect 22002 17926 22014 17978
rect 22066 17926 22078 17978
rect 22130 17926 22142 17978
rect 22194 17926 22206 17978
rect 22258 17926 26950 17978
rect 27002 17926 27014 17978
rect 27066 17926 27078 17978
rect 27130 17926 27142 17978
rect 27194 17926 27206 17978
rect 27258 17926 31950 17978
rect 32002 17926 32014 17978
rect 32066 17926 32078 17978
rect 32130 17926 32142 17978
rect 32194 17926 32206 17978
rect 32258 17926 36950 17978
rect 37002 17926 37014 17978
rect 37066 17926 37078 17978
rect 37130 17926 37142 17978
rect 37194 17926 37206 17978
rect 37258 17926 40848 17978
rect 1104 17904 40848 17926
rect 20806 17824 20812 17876
rect 20864 17864 20870 17876
rect 21174 17864 21180 17876
rect 20864 17836 21180 17864
rect 20864 17824 20870 17836
rect 21174 17824 21180 17836
rect 21232 17864 21238 17876
rect 36446 17864 36452 17876
rect 21232 17836 36452 17864
rect 21232 17824 21238 17836
rect 36446 17824 36452 17836
rect 36504 17824 36510 17876
rect 3878 17620 3884 17672
rect 3936 17660 3942 17672
rect 3936 17632 16574 17660
rect 3936 17620 3942 17632
rect 3326 17552 3332 17604
rect 3384 17592 3390 17604
rect 8662 17592 8668 17604
rect 3384 17564 8668 17592
rect 3384 17552 3390 17564
rect 8662 17552 8668 17564
rect 8720 17592 8726 17604
rect 9122 17592 9128 17604
rect 8720 17564 9128 17592
rect 8720 17552 8726 17564
rect 9122 17552 9128 17564
rect 9180 17552 9186 17604
rect 2958 17484 2964 17536
rect 3016 17524 3022 17536
rect 7466 17524 7472 17536
rect 3016 17496 7472 17524
rect 3016 17484 3022 17496
rect 7466 17484 7472 17496
rect 7524 17484 7530 17536
rect 16546 17524 16574 17632
rect 18506 17552 18512 17604
rect 18564 17592 18570 17604
rect 38194 17592 38200 17604
rect 18564 17564 38200 17592
rect 18564 17552 18570 17564
rect 38194 17552 38200 17564
rect 38252 17552 38258 17604
rect 36538 17524 36544 17536
rect 16546 17496 36544 17524
rect 36538 17484 36544 17496
rect 36596 17484 36602 17536
rect 1104 17434 40848 17456
rect 1104 17382 2610 17434
rect 2662 17382 2674 17434
rect 2726 17382 2738 17434
rect 2790 17382 2802 17434
rect 2854 17382 2866 17434
rect 2918 17382 7610 17434
rect 7662 17382 7674 17434
rect 7726 17382 7738 17434
rect 7790 17382 7802 17434
rect 7854 17382 7866 17434
rect 7918 17382 12610 17434
rect 12662 17382 12674 17434
rect 12726 17382 12738 17434
rect 12790 17382 12802 17434
rect 12854 17382 12866 17434
rect 12918 17382 17610 17434
rect 17662 17382 17674 17434
rect 17726 17382 17738 17434
rect 17790 17382 17802 17434
rect 17854 17382 17866 17434
rect 17918 17382 22610 17434
rect 22662 17382 22674 17434
rect 22726 17382 22738 17434
rect 22790 17382 22802 17434
rect 22854 17382 22866 17434
rect 22918 17382 27610 17434
rect 27662 17382 27674 17434
rect 27726 17382 27738 17434
rect 27790 17382 27802 17434
rect 27854 17382 27866 17434
rect 27918 17382 32610 17434
rect 32662 17382 32674 17434
rect 32726 17382 32738 17434
rect 32790 17382 32802 17434
rect 32854 17382 32866 17434
rect 32918 17382 37610 17434
rect 37662 17382 37674 17434
rect 37726 17382 37738 17434
rect 37790 17382 37802 17434
rect 37854 17382 37866 17434
rect 37918 17382 40848 17434
rect 1104 17360 40848 17382
rect 3326 17280 3332 17332
rect 3384 17280 3390 17332
rect 3620 17292 6914 17320
rect 2869 17255 2927 17261
rect 2869 17221 2881 17255
rect 2915 17252 2927 17255
rect 2958 17252 2964 17264
rect 2915 17224 2964 17252
rect 2915 17221 2927 17224
rect 2869 17215 2927 17221
rect 2958 17212 2964 17224
rect 3016 17212 3022 17264
rect 3620 17261 3648 17292
rect 3237 17255 3295 17261
rect 3237 17221 3249 17255
rect 3283 17252 3295 17255
rect 3605 17255 3663 17261
rect 3283 17224 3556 17252
rect 3283 17221 3295 17224
rect 3237 17215 3295 17221
rect 3421 17187 3479 17193
rect 3421 17153 3433 17187
rect 3467 17153 3479 17187
rect 3528 17184 3556 17224
rect 3605 17221 3617 17255
rect 3651 17221 3663 17255
rect 3605 17215 3663 17221
rect 3878 17212 3884 17264
rect 3936 17252 3942 17264
rect 4525 17255 4583 17261
rect 4525 17252 4537 17255
rect 3936 17224 4537 17252
rect 3936 17212 3942 17224
rect 4525 17221 4537 17224
rect 4571 17221 4583 17255
rect 4525 17215 4583 17221
rect 4709 17255 4767 17261
rect 4709 17221 4721 17255
rect 4755 17252 4767 17255
rect 6454 17252 6460 17264
rect 4755 17224 6460 17252
rect 4755 17221 4767 17224
rect 4709 17215 4767 17221
rect 6454 17212 6460 17224
rect 6512 17212 6518 17264
rect 6178 17184 6184 17196
rect 3528 17156 6184 17184
rect 3421 17147 3479 17153
rect 3436 17116 3464 17147
rect 6178 17144 6184 17156
rect 6236 17144 6242 17196
rect 5718 17116 5724 17128
rect 3436 17088 5724 17116
rect 5718 17076 5724 17088
rect 5776 17076 5782 17128
rect 6886 17116 6914 17292
rect 18414 17280 18420 17332
rect 18472 17320 18478 17332
rect 18598 17320 18604 17332
rect 18472 17292 18604 17320
rect 18472 17280 18478 17292
rect 18598 17280 18604 17292
rect 18656 17320 18662 17332
rect 18693 17323 18751 17329
rect 18693 17320 18705 17323
rect 18656 17292 18705 17320
rect 18656 17280 18662 17292
rect 18693 17289 18705 17292
rect 18739 17289 18751 17323
rect 18693 17283 18751 17289
rect 18782 17280 18788 17332
rect 18840 17280 18846 17332
rect 31573 17323 31631 17329
rect 31573 17289 31585 17323
rect 31619 17320 31631 17323
rect 33962 17320 33968 17332
rect 31619 17292 33968 17320
rect 31619 17289 31631 17292
rect 31573 17283 31631 17289
rect 33962 17280 33968 17292
rect 34020 17280 34026 17332
rect 18506 17212 18512 17264
rect 18564 17212 18570 17264
rect 18874 17212 18880 17264
rect 18932 17212 18938 17264
rect 19245 17255 19303 17261
rect 19245 17221 19257 17255
rect 19291 17252 19303 17255
rect 20438 17252 20444 17264
rect 19291 17224 20444 17252
rect 19291 17221 19303 17224
rect 19245 17215 19303 17221
rect 20438 17212 20444 17224
rect 20496 17212 20502 17264
rect 28718 17212 28724 17264
rect 28776 17212 28782 17264
rect 28902 17212 28908 17264
rect 28960 17212 28966 17264
rect 28994 17212 29000 17264
rect 29052 17252 29058 17264
rect 29052 17224 31616 17252
rect 29052 17212 29058 17224
rect 19518 17144 19524 17196
rect 19576 17144 19582 17196
rect 29086 17144 29092 17196
rect 29144 17184 29150 17196
rect 31588 17193 31616 17224
rect 31389 17187 31447 17193
rect 31389 17184 31401 17187
rect 29144 17156 31401 17184
rect 29144 17144 29150 17156
rect 31389 17153 31401 17156
rect 31435 17153 31447 17187
rect 31389 17147 31447 17153
rect 31573 17187 31631 17193
rect 31573 17153 31585 17187
rect 31619 17153 31631 17187
rect 31573 17147 31631 17153
rect 21726 17116 21732 17128
rect 6886 17088 21732 17116
rect 21726 17076 21732 17088
rect 21784 17076 21790 17128
rect 4341 17051 4399 17057
rect 4341 17017 4353 17051
rect 4387 17048 4399 17051
rect 15654 17048 15660 17060
rect 4387 17020 15660 17048
rect 4387 17017 4399 17020
rect 4341 17011 4399 17017
rect 15654 17008 15660 17020
rect 15712 17008 15718 17060
rect 1670 16940 1676 16992
rect 1728 16980 1734 16992
rect 3878 16980 3884 16992
rect 1728 16952 3884 16980
rect 1728 16940 1734 16952
rect 3878 16940 3884 16952
rect 3936 16940 3942 16992
rect 4522 16940 4528 16992
rect 4580 16940 4586 16992
rect 17310 16940 17316 16992
rect 17368 16980 17374 16992
rect 19429 16983 19487 16989
rect 19429 16980 19441 16983
rect 17368 16952 19441 16980
rect 17368 16940 17374 16952
rect 19429 16949 19441 16952
rect 19475 16949 19487 16983
rect 19429 16943 19487 16949
rect 28534 16940 28540 16992
rect 28592 16940 28598 16992
rect 1104 16890 40848 16912
rect 1104 16838 1950 16890
rect 2002 16838 2014 16890
rect 2066 16838 2078 16890
rect 2130 16838 2142 16890
rect 2194 16838 2206 16890
rect 2258 16838 6950 16890
rect 7002 16838 7014 16890
rect 7066 16838 7078 16890
rect 7130 16838 7142 16890
rect 7194 16838 7206 16890
rect 7258 16838 11950 16890
rect 12002 16838 12014 16890
rect 12066 16838 12078 16890
rect 12130 16838 12142 16890
rect 12194 16838 12206 16890
rect 12258 16838 16950 16890
rect 17002 16838 17014 16890
rect 17066 16838 17078 16890
rect 17130 16838 17142 16890
rect 17194 16838 17206 16890
rect 17258 16838 21950 16890
rect 22002 16838 22014 16890
rect 22066 16838 22078 16890
rect 22130 16838 22142 16890
rect 22194 16838 22206 16890
rect 22258 16838 26950 16890
rect 27002 16838 27014 16890
rect 27066 16838 27078 16890
rect 27130 16838 27142 16890
rect 27194 16838 27206 16890
rect 27258 16838 31950 16890
rect 32002 16838 32014 16890
rect 32066 16838 32078 16890
rect 32130 16838 32142 16890
rect 32194 16838 32206 16890
rect 32258 16838 36950 16890
rect 37002 16838 37014 16890
rect 37066 16838 37078 16890
rect 37130 16838 37142 16890
rect 37194 16838 37206 16890
rect 37258 16838 40848 16890
rect 1104 16816 40848 16838
rect 4522 16736 4528 16788
rect 4580 16776 4586 16788
rect 28534 16776 28540 16788
rect 4580 16748 28540 16776
rect 4580 16736 4586 16748
rect 28534 16736 28540 16748
rect 28592 16736 28598 16788
rect 14274 16600 14280 16652
rect 14332 16600 14338 16652
rect 15749 16643 15807 16649
rect 15749 16609 15761 16643
rect 15795 16640 15807 16643
rect 21174 16640 21180 16652
rect 15795 16612 21180 16640
rect 15795 16609 15807 16612
rect 15749 16603 15807 16609
rect 21174 16600 21180 16612
rect 21232 16600 21238 16652
rect 23382 16600 23388 16652
rect 23440 16640 23446 16652
rect 30834 16640 30840 16652
rect 23440 16612 30840 16640
rect 23440 16600 23446 16612
rect 30834 16600 30840 16612
rect 30892 16600 30898 16652
rect 31110 16600 31116 16652
rect 31168 16600 31174 16652
rect 14734 16532 14740 16584
rect 14792 16532 14798 16584
rect 15010 16532 15016 16584
rect 15068 16532 15074 16584
rect 15197 16575 15255 16581
rect 15197 16541 15209 16575
rect 15243 16572 15255 16575
rect 15470 16572 15476 16584
rect 15243 16544 15476 16572
rect 15243 16541 15255 16544
rect 15197 16535 15255 16541
rect 15470 16532 15476 16544
rect 15528 16532 15534 16584
rect 15565 16575 15623 16581
rect 15565 16541 15577 16575
rect 15611 16572 15623 16575
rect 32861 16575 32919 16581
rect 15611 16544 16574 16572
rect 15611 16541 15623 16544
rect 15565 16535 15623 16541
rect 16546 16436 16574 16544
rect 32861 16541 32873 16575
rect 32907 16572 32919 16575
rect 34974 16572 34980 16584
rect 32907 16544 34980 16572
rect 32907 16541 32919 16544
rect 32861 16535 32919 16541
rect 34974 16532 34980 16544
rect 35032 16532 35038 16584
rect 18690 16464 18696 16516
rect 18748 16504 18754 16516
rect 18748 16476 31602 16504
rect 18748 16464 18754 16476
rect 39758 16436 39764 16448
rect 16546 16408 39764 16436
rect 39758 16396 39764 16408
rect 39816 16396 39822 16448
rect 1104 16346 40848 16368
rect 1104 16294 2610 16346
rect 2662 16294 2674 16346
rect 2726 16294 2738 16346
rect 2790 16294 2802 16346
rect 2854 16294 2866 16346
rect 2918 16294 7610 16346
rect 7662 16294 7674 16346
rect 7726 16294 7738 16346
rect 7790 16294 7802 16346
rect 7854 16294 7866 16346
rect 7918 16294 12610 16346
rect 12662 16294 12674 16346
rect 12726 16294 12738 16346
rect 12790 16294 12802 16346
rect 12854 16294 12866 16346
rect 12918 16294 17610 16346
rect 17662 16294 17674 16346
rect 17726 16294 17738 16346
rect 17790 16294 17802 16346
rect 17854 16294 17866 16346
rect 17918 16294 22610 16346
rect 22662 16294 22674 16346
rect 22726 16294 22738 16346
rect 22790 16294 22802 16346
rect 22854 16294 22866 16346
rect 22918 16294 27610 16346
rect 27662 16294 27674 16346
rect 27726 16294 27738 16346
rect 27790 16294 27802 16346
rect 27854 16294 27866 16346
rect 27918 16294 32610 16346
rect 32662 16294 32674 16346
rect 32726 16294 32738 16346
rect 32790 16294 32802 16346
rect 32854 16294 32866 16346
rect 32918 16294 37610 16346
rect 37662 16294 37674 16346
rect 37726 16294 37738 16346
rect 37790 16294 37802 16346
rect 37854 16294 37866 16346
rect 37918 16294 40848 16346
rect 1104 16272 40848 16294
rect 15010 16192 15016 16244
rect 15068 16232 15074 16244
rect 20898 16232 20904 16244
rect 15068 16204 20904 16232
rect 15068 16192 15074 16204
rect 20898 16192 20904 16204
rect 20956 16192 20962 16244
rect 22738 15852 22744 15904
rect 22796 15892 22802 15904
rect 23290 15892 23296 15904
rect 22796 15864 23296 15892
rect 22796 15852 22802 15864
rect 23290 15852 23296 15864
rect 23348 15892 23354 15904
rect 38194 15892 38200 15904
rect 23348 15864 38200 15892
rect 23348 15852 23354 15864
rect 38194 15852 38200 15864
rect 38252 15852 38258 15904
rect 1104 15802 40848 15824
rect 1104 15750 1950 15802
rect 2002 15750 2014 15802
rect 2066 15750 2078 15802
rect 2130 15750 2142 15802
rect 2194 15750 2206 15802
rect 2258 15750 6950 15802
rect 7002 15750 7014 15802
rect 7066 15750 7078 15802
rect 7130 15750 7142 15802
rect 7194 15750 7206 15802
rect 7258 15750 11950 15802
rect 12002 15750 12014 15802
rect 12066 15750 12078 15802
rect 12130 15750 12142 15802
rect 12194 15750 12206 15802
rect 12258 15750 16950 15802
rect 17002 15750 17014 15802
rect 17066 15750 17078 15802
rect 17130 15750 17142 15802
rect 17194 15750 17206 15802
rect 17258 15750 21950 15802
rect 22002 15750 22014 15802
rect 22066 15750 22078 15802
rect 22130 15750 22142 15802
rect 22194 15750 22206 15802
rect 22258 15750 26950 15802
rect 27002 15750 27014 15802
rect 27066 15750 27078 15802
rect 27130 15750 27142 15802
rect 27194 15750 27206 15802
rect 27258 15750 31950 15802
rect 32002 15750 32014 15802
rect 32066 15750 32078 15802
rect 32130 15750 32142 15802
rect 32194 15750 32206 15802
rect 32258 15750 36950 15802
rect 37002 15750 37014 15802
rect 37066 15750 37078 15802
rect 37130 15750 37142 15802
rect 37194 15750 37206 15802
rect 37258 15750 40848 15802
rect 1104 15728 40848 15750
rect 14090 15444 14096 15496
rect 14148 15444 14154 15496
rect 14366 15444 14372 15496
rect 14424 15444 14430 15496
rect 22738 15416 22744 15428
rect 14200 15388 22744 15416
rect 14200 15360 14228 15388
rect 22738 15376 22744 15388
rect 22796 15376 22802 15428
rect 14182 15308 14188 15360
rect 14240 15308 14246 15360
rect 14553 15351 14611 15357
rect 14553 15317 14565 15351
rect 14599 15348 14611 15351
rect 33226 15348 33232 15360
rect 14599 15320 33232 15348
rect 14599 15317 14611 15320
rect 14553 15311 14611 15317
rect 33226 15308 33232 15320
rect 33284 15308 33290 15360
rect 1104 15258 40848 15280
rect 1104 15206 2610 15258
rect 2662 15206 2674 15258
rect 2726 15206 2738 15258
rect 2790 15206 2802 15258
rect 2854 15206 2866 15258
rect 2918 15206 7610 15258
rect 7662 15206 7674 15258
rect 7726 15206 7738 15258
rect 7790 15206 7802 15258
rect 7854 15206 7866 15258
rect 7918 15206 12610 15258
rect 12662 15206 12674 15258
rect 12726 15206 12738 15258
rect 12790 15206 12802 15258
rect 12854 15206 12866 15258
rect 12918 15206 17610 15258
rect 17662 15206 17674 15258
rect 17726 15206 17738 15258
rect 17790 15206 17802 15258
rect 17854 15206 17866 15258
rect 17918 15206 22610 15258
rect 22662 15206 22674 15258
rect 22726 15206 22738 15258
rect 22790 15206 22802 15258
rect 22854 15206 22866 15258
rect 22918 15206 27610 15258
rect 27662 15206 27674 15258
rect 27726 15206 27738 15258
rect 27790 15206 27802 15258
rect 27854 15206 27866 15258
rect 27918 15206 32610 15258
rect 32662 15206 32674 15258
rect 32726 15206 32738 15258
rect 32790 15206 32802 15258
rect 32854 15206 32866 15258
rect 32918 15206 37610 15258
rect 37662 15206 37674 15258
rect 37726 15206 37738 15258
rect 37790 15206 37802 15258
rect 37854 15206 37866 15258
rect 37918 15206 40848 15258
rect 1104 15184 40848 15206
rect 31202 15036 31208 15088
rect 31260 15076 31266 15088
rect 32309 15079 32367 15085
rect 32309 15076 32321 15079
rect 31260 15048 32321 15076
rect 31260 15036 31266 15048
rect 32309 15045 32321 15048
rect 32355 15045 32367 15079
rect 32309 15039 32367 15045
rect 32398 15036 32404 15088
rect 32456 15076 32462 15088
rect 32493 15079 32551 15085
rect 32493 15076 32505 15079
rect 32456 15048 32505 15076
rect 32456 15036 32462 15048
rect 32493 15045 32505 15048
rect 32539 15045 32551 15079
rect 32493 15039 32551 15045
rect 38010 14968 38016 15020
rect 38068 14968 38074 15020
rect 38194 14968 38200 15020
rect 38252 14968 38258 15020
rect 33318 14832 33324 14884
rect 33376 14872 33382 14884
rect 38105 14875 38163 14881
rect 38105 14872 38117 14875
rect 33376 14844 38117 14872
rect 33376 14832 33382 14844
rect 38105 14841 38117 14844
rect 38151 14841 38163 14875
rect 38105 14835 38163 14841
rect 24762 14764 24768 14816
rect 24820 14804 24826 14816
rect 32217 14807 32275 14813
rect 32217 14804 32229 14807
rect 24820 14776 32229 14804
rect 24820 14764 24826 14776
rect 32217 14773 32229 14776
rect 32263 14773 32275 14807
rect 32217 14767 32275 14773
rect 1104 14714 40848 14736
rect 1104 14662 1950 14714
rect 2002 14662 2014 14714
rect 2066 14662 2078 14714
rect 2130 14662 2142 14714
rect 2194 14662 2206 14714
rect 2258 14662 6950 14714
rect 7002 14662 7014 14714
rect 7066 14662 7078 14714
rect 7130 14662 7142 14714
rect 7194 14662 7206 14714
rect 7258 14662 11950 14714
rect 12002 14662 12014 14714
rect 12066 14662 12078 14714
rect 12130 14662 12142 14714
rect 12194 14662 12206 14714
rect 12258 14662 16950 14714
rect 17002 14662 17014 14714
rect 17066 14662 17078 14714
rect 17130 14662 17142 14714
rect 17194 14662 17206 14714
rect 17258 14662 21950 14714
rect 22002 14662 22014 14714
rect 22066 14662 22078 14714
rect 22130 14662 22142 14714
rect 22194 14662 22206 14714
rect 22258 14662 26950 14714
rect 27002 14662 27014 14714
rect 27066 14662 27078 14714
rect 27130 14662 27142 14714
rect 27194 14662 27206 14714
rect 27258 14662 31950 14714
rect 32002 14662 32014 14714
rect 32066 14662 32078 14714
rect 32130 14662 32142 14714
rect 32194 14662 32206 14714
rect 32258 14662 36950 14714
rect 37002 14662 37014 14714
rect 37066 14662 37078 14714
rect 37130 14662 37142 14714
rect 37194 14662 37206 14714
rect 37258 14662 40848 14714
rect 1104 14640 40848 14662
rect 31018 14356 31024 14408
rect 31076 14396 31082 14408
rect 38565 14399 38623 14405
rect 38565 14396 38577 14399
rect 31076 14368 38577 14396
rect 31076 14356 31082 14368
rect 38565 14365 38577 14368
rect 38611 14365 38623 14399
rect 38565 14359 38623 14365
rect 38930 14356 38936 14408
rect 38988 14356 38994 14408
rect 18598 14288 18604 14340
rect 18656 14328 18662 14340
rect 38749 14331 38807 14337
rect 38749 14328 38761 14331
rect 18656 14300 38761 14328
rect 18656 14288 18662 14300
rect 38749 14297 38761 14300
rect 38795 14297 38807 14331
rect 38749 14291 38807 14297
rect 1104 14170 40848 14192
rect 1104 14118 2610 14170
rect 2662 14118 2674 14170
rect 2726 14118 2738 14170
rect 2790 14118 2802 14170
rect 2854 14118 2866 14170
rect 2918 14118 7610 14170
rect 7662 14118 7674 14170
rect 7726 14118 7738 14170
rect 7790 14118 7802 14170
rect 7854 14118 7866 14170
rect 7918 14118 12610 14170
rect 12662 14118 12674 14170
rect 12726 14118 12738 14170
rect 12790 14118 12802 14170
rect 12854 14118 12866 14170
rect 12918 14118 17610 14170
rect 17662 14118 17674 14170
rect 17726 14118 17738 14170
rect 17790 14118 17802 14170
rect 17854 14118 17866 14170
rect 17918 14118 22610 14170
rect 22662 14118 22674 14170
rect 22726 14118 22738 14170
rect 22790 14118 22802 14170
rect 22854 14118 22866 14170
rect 22918 14118 27610 14170
rect 27662 14118 27674 14170
rect 27726 14118 27738 14170
rect 27790 14118 27802 14170
rect 27854 14118 27866 14170
rect 27918 14118 32610 14170
rect 32662 14118 32674 14170
rect 32726 14118 32738 14170
rect 32790 14118 32802 14170
rect 32854 14118 32866 14170
rect 32918 14118 37610 14170
rect 37662 14118 37674 14170
rect 37726 14118 37738 14170
rect 37790 14118 37802 14170
rect 37854 14118 37866 14170
rect 37918 14118 40848 14170
rect 1104 14096 40848 14118
rect 9766 14016 9772 14068
rect 9824 14056 9830 14068
rect 28537 14059 28595 14065
rect 28537 14056 28549 14059
rect 9824 14028 28549 14056
rect 9824 14016 9830 14028
rect 28537 14025 28549 14028
rect 28583 14025 28595 14059
rect 28537 14019 28595 14025
rect 8018 13948 8024 14000
rect 8076 13988 8082 14000
rect 14645 13991 14703 13997
rect 8076 13960 13386 13988
rect 8076 13948 8082 13960
rect 14645 13957 14657 13991
rect 14691 13988 14703 13991
rect 18598 13988 18604 14000
rect 14691 13960 18604 13988
rect 14691 13957 14703 13960
rect 14645 13951 14703 13957
rect 18598 13948 18604 13960
rect 18656 13948 18662 14000
rect 28629 13923 28687 13929
rect 28629 13889 28641 13923
rect 28675 13920 28687 13923
rect 29730 13920 29736 13932
rect 28675 13892 29736 13920
rect 28675 13889 28687 13892
rect 28629 13883 28687 13889
rect 29730 13880 29736 13892
rect 29788 13880 29794 13932
rect 9582 13812 9588 13864
rect 9640 13852 9646 13864
rect 12621 13855 12679 13861
rect 12621 13852 12633 13855
rect 9640 13824 12633 13852
rect 9640 13812 9646 13824
rect 12621 13821 12633 13824
rect 12667 13821 12679 13855
rect 12621 13815 12679 13821
rect 12884 13719 12942 13725
rect 12884 13685 12896 13719
rect 12930 13716 12942 13719
rect 13630 13716 13636 13728
rect 12930 13688 13636 13716
rect 12930 13685 12942 13688
rect 12884 13679 12942 13685
rect 13630 13676 13636 13688
rect 13688 13676 13694 13728
rect 1104 13626 40848 13648
rect 1104 13574 1950 13626
rect 2002 13574 2014 13626
rect 2066 13574 2078 13626
rect 2130 13574 2142 13626
rect 2194 13574 2206 13626
rect 2258 13574 6950 13626
rect 7002 13574 7014 13626
rect 7066 13574 7078 13626
rect 7130 13574 7142 13626
rect 7194 13574 7206 13626
rect 7258 13574 11950 13626
rect 12002 13574 12014 13626
rect 12066 13574 12078 13626
rect 12130 13574 12142 13626
rect 12194 13574 12206 13626
rect 12258 13574 16950 13626
rect 17002 13574 17014 13626
rect 17066 13574 17078 13626
rect 17130 13574 17142 13626
rect 17194 13574 17206 13626
rect 17258 13574 21950 13626
rect 22002 13574 22014 13626
rect 22066 13574 22078 13626
rect 22130 13574 22142 13626
rect 22194 13574 22206 13626
rect 22258 13574 26950 13626
rect 27002 13574 27014 13626
rect 27066 13574 27078 13626
rect 27130 13574 27142 13626
rect 27194 13574 27206 13626
rect 27258 13574 31950 13626
rect 32002 13574 32014 13626
rect 32066 13574 32078 13626
rect 32130 13574 32142 13626
rect 32194 13574 32206 13626
rect 32258 13574 36950 13626
rect 37002 13574 37014 13626
rect 37066 13574 37078 13626
rect 37130 13574 37142 13626
rect 37194 13574 37206 13626
rect 37258 13574 40848 13626
rect 1104 13552 40848 13574
rect 27522 13472 27528 13524
rect 27580 13512 27586 13524
rect 27985 13515 28043 13521
rect 27985 13512 27997 13515
rect 27580 13484 27997 13512
rect 27580 13472 27586 13484
rect 27985 13481 27997 13484
rect 28031 13481 28043 13515
rect 27985 13475 28043 13481
rect 34882 13336 34888 13388
rect 34940 13376 34946 13388
rect 36541 13379 36599 13385
rect 36541 13376 36553 13379
rect 34940 13348 36553 13376
rect 34940 13336 34946 13348
rect 36541 13345 36553 13348
rect 36587 13345 36599 13379
rect 39666 13376 39672 13388
rect 36541 13339 36599 13345
rect 36740 13348 39672 13376
rect 15838 13268 15844 13320
rect 15896 13308 15902 13320
rect 16482 13308 16488 13320
rect 15896 13280 16488 13308
rect 15896 13268 15902 13280
rect 16482 13268 16488 13280
rect 16540 13308 16546 13320
rect 36740 13317 36768 13348
rect 39666 13336 39672 13348
rect 39724 13336 39730 13388
rect 28077 13311 28135 13317
rect 28077 13308 28089 13311
rect 16540 13280 28089 13308
rect 16540 13268 16546 13280
rect 28077 13277 28089 13280
rect 28123 13277 28135 13311
rect 28077 13271 28135 13277
rect 36725 13311 36783 13317
rect 36725 13277 36737 13311
rect 36771 13277 36783 13311
rect 36725 13271 36783 13277
rect 36817 13311 36875 13317
rect 36817 13277 36829 13311
rect 36863 13277 36875 13311
rect 36817 13271 36875 13277
rect 36446 13200 36452 13252
rect 36504 13240 36510 13252
rect 36832 13240 36860 13271
rect 36504 13212 36860 13240
rect 36504 13200 36510 13212
rect 1104 13082 40848 13104
rect 1104 13030 2610 13082
rect 2662 13030 2674 13082
rect 2726 13030 2738 13082
rect 2790 13030 2802 13082
rect 2854 13030 2866 13082
rect 2918 13030 7610 13082
rect 7662 13030 7674 13082
rect 7726 13030 7738 13082
rect 7790 13030 7802 13082
rect 7854 13030 7866 13082
rect 7918 13030 12610 13082
rect 12662 13030 12674 13082
rect 12726 13030 12738 13082
rect 12790 13030 12802 13082
rect 12854 13030 12866 13082
rect 12918 13030 17610 13082
rect 17662 13030 17674 13082
rect 17726 13030 17738 13082
rect 17790 13030 17802 13082
rect 17854 13030 17866 13082
rect 17918 13030 22610 13082
rect 22662 13030 22674 13082
rect 22726 13030 22738 13082
rect 22790 13030 22802 13082
rect 22854 13030 22866 13082
rect 22918 13030 27610 13082
rect 27662 13030 27674 13082
rect 27726 13030 27738 13082
rect 27790 13030 27802 13082
rect 27854 13030 27866 13082
rect 27918 13030 32610 13082
rect 32662 13030 32674 13082
rect 32726 13030 32738 13082
rect 32790 13030 32802 13082
rect 32854 13030 32866 13082
rect 32918 13030 37610 13082
rect 37662 13030 37674 13082
rect 37726 13030 37738 13082
rect 37790 13030 37802 13082
rect 37854 13030 37866 13082
rect 37918 13030 40848 13082
rect 1104 13008 40848 13030
rect 1104 12538 40848 12560
rect 1104 12486 1950 12538
rect 2002 12486 2014 12538
rect 2066 12486 2078 12538
rect 2130 12486 2142 12538
rect 2194 12486 2206 12538
rect 2258 12486 6950 12538
rect 7002 12486 7014 12538
rect 7066 12486 7078 12538
rect 7130 12486 7142 12538
rect 7194 12486 7206 12538
rect 7258 12486 11950 12538
rect 12002 12486 12014 12538
rect 12066 12486 12078 12538
rect 12130 12486 12142 12538
rect 12194 12486 12206 12538
rect 12258 12486 16950 12538
rect 17002 12486 17014 12538
rect 17066 12486 17078 12538
rect 17130 12486 17142 12538
rect 17194 12486 17206 12538
rect 17258 12486 21950 12538
rect 22002 12486 22014 12538
rect 22066 12486 22078 12538
rect 22130 12486 22142 12538
rect 22194 12486 22206 12538
rect 22258 12486 26950 12538
rect 27002 12486 27014 12538
rect 27066 12486 27078 12538
rect 27130 12486 27142 12538
rect 27194 12486 27206 12538
rect 27258 12486 31950 12538
rect 32002 12486 32014 12538
rect 32066 12486 32078 12538
rect 32130 12486 32142 12538
rect 32194 12486 32206 12538
rect 32258 12486 36950 12538
rect 37002 12486 37014 12538
rect 37066 12486 37078 12538
rect 37130 12486 37142 12538
rect 37194 12486 37206 12538
rect 37258 12486 40848 12538
rect 1104 12464 40848 12486
rect 4801 12223 4859 12229
rect 4801 12189 4813 12223
rect 4847 12220 4859 12223
rect 18046 12220 18052 12232
rect 4847 12192 18052 12220
rect 4847 12189 4859 12192
rect 4801 12183 4859 12189
rect 18046 12180 18052 12192
rect 18104 12220 18110 12232
rect 18598 12220 18604 12232
rect 18104 12192 18604 12220
rect 18104 12180 18110 12192
rect 18598 12180 18604 12192
rect 18656 12180 18662 12232
rect 18782 12180 18788 12232
rect 18840 12220 18846 12232
rect 23569 12223 23627 12229
rect 23569 12220 23581 12223
rect 18840 12192 23581 12220
rect 18840 12180 18846 12192
rect 23569 12189 23581 12192
rect 23615 12189 23627 12223
rect 23569 12183 23627 12189
rect 4706 12044 4712 12096
rect 4764 12044 4770 12096
rect 23584 12084 23612 12183
rect 23750 12180 23756 12232
rect 23808 12180 23814 12232
rect 23937 12155 23995 12161
rect 23937 12121 23949 12155
rect 23983 12152 23995 12155
rect 38470 12152 38476 12164
rect 23983 12124 38476 12152
rect 23983 12121 23995 12124
rect 23937 12115 23995 12121
rect 38470 12112 38476 12124
rect 38528 12112 38534 12164
rect 25774 12084 25780 12096
rect 23584 12056 25780 12084
rect 25774 12044 25780 12056
rect 25832 12044 25838 12096
rect 1104 11994 40848 12016
rect 1104 11942 2610 11994
rect 2662 11942 2674 11994
rect 2726 11942 2738 11994
rect 2790 11942 2802 11994
rect 2854 11942 2866 11994
rect 2918 11942 7610 11994
rect 7662 11942 7674 11994
rect 7726 11942 7738 11994
rect 7790 11942 7802 11994
rect 7854 11942 7866 11994
rect 7918 11942 12610 11994
rect 12662 11942 12674 11994
rect 12726 11942 12738 11994
rect 12790 11942 12802 11994
rect 12854 11942 12866 11994
rect 12918 11942 17610 11994
rect 17662 11942 17674 11994
rect 17726 11942 17738 11994
rect 17790 11942 17802 11994
rect 17854 11942 17866 11994
rect 17918 11942 22610 11994
rect 22662 11942 22674 11994
rect 22726 11942 22738 11994
rect 22790 11942 22802 11994
rect 22854 11942 22866 11994
rect 22918 11942 27610 11994
rect 27662 11942 27674 11994
rect 27726 11942 27738 11994
rect 27790 11942 27802 11994
rect 27854 11942 27866 11994
rect 27918 11942 32610 11994
rect 32662 11942 32674 11994
rect 32726 11942 32738 11994
rect 32790 11942 32802 11994
rect 32854 11942 32866 11994
rect 32918 11942 37610 11994
rect 37662 11942 37674 11994
rect 37726 11942 37738 11994
rect 37790 11942 37802 11994
rect 37854 11942 37866 11994
rect 37918 11942 40848 11994
rect 1104 11920 40848 11942
rect 1104 11450 40848 11472
rect 1104 11398 1950 11450
rect 2002 11398 2014 11450
rect 2066 11398 2078 11450
rect 2130 11398 2142 11450
rect 2194 11398 2206 11450
rect 2258 11398 6950 11450
rect 7002 11398 7014 11450
rect 7066 11398 7078 11450
rect 7130 11398 7142 11450
rect 7194 11398 7206 11450
rect 7258 11398 11950 11450
rect 12002 11398 12014 11450
rect 12066 11398 12078 11450
rect 12130 11398 12142 11450
rect 12194 11398 12206 11450
rect 12258 11398 16950 11450
rect 17002 11398 17014 11450
rect 17066 11398 17078 11450
rect 17130 11398 17142 11450
rect 17194 11398 17206 11450
rect 17258 11398 21950 11450
rect 22002 11398 22014 11450
rect 22066 11398 22078 11450
rect 22130 11398 22142 11450
rect 22194 11398 22206 11450
rect 22258 11398 26950 11450
rect 27002 11398 27014 11450
rect 27066 11398 27078 11450
rect 27130 11398 27142 11450
rect 27194 11398 27206 11450
rect 27258 11398 31950 11450
rect 32002 11398 32014 11450
rect 32066 11398 32078 11450
rect 32130 11398 32142 11450
rect 32194 11398 32206 11450
rect 32258 11398 36950 11450
rect 37002 11398 37014 11450
rect 37066 11398 37078 11450
rect 37130 11398 37142 11450
rect 37194 11398 37206 11450
rect 37258 11398 40848 11450
rect 1104 11376 40848 11398
rect 29638 11228 29644 11280
rect 29696 11268 29702 11280
rect 29696 11240 31248 11268
rect 29696 11228 29702 11240
rect 30834 11160 30840 11212
rect 30892 11200 30898 11212
rect 31113 11203 31171 11209
rect 31113 11200 31125 11203
rect 30892 11172 31125 11200
rect 30892 11160 30898 11172
rect 31113 11169 31125 11172
rect 31159 11169 31171 11203
rect 31220 11200 31248 11240
rect 31220 11172 32536 11200
rect 31113 11163 31171 11169
rect 32508 11118 32536 11172
rect 33042 11160 33048 11212
rect 33100 11200 33106 11212
rect 33137 11203 33195 11209
rect 33137 11200 33149 11203
rect 33100 11172 33149 11200
rect 33100 11160 33106 11172
rect 33137 11169 33149 11172
rect 33183 11169 33195 11203
rect 33137 11163 33195 11169
rect 6546 11024 6552 11076
rect 6604 11064 6610 11076
rect 30745 11067 30803 11073
rect 30745 11064 30757 11067
rect 6604 11036 30757 11064
rect 6604 11024 6610 11036
rect 30745 11033 30757 11036
rect 30791 11064 30803 11067
rect 31389 11067 31447 11073
rect 31389 11064 31401 11067
rect 30791 11036 31401 11064
rect 30791 11033 30803 11036
rect 30745 11027 30803 11033
rect 31389 11033 31401 11036
rect 31435 11033 31447 11067
rect 31389 11027 31447 11033
rect 1104 10906 40848 10928
rect 1104 10854 2610 10906
rect 2662 10854 2674 10906
rect 2726 10854 2738 10906
rect 2790 10854 2802 10906
rect 2854 10854 2866 10906
rect 2918 10854 7610 10906
rect 7662 10854 7674 10906
rect 7726 10854 7738 10906
rect 7790 10854 7802 10906
rect 7854 10854 7866 10906
rect 7918 10854 12610 10906
rect 12662 10854 12674 10906
rect 12726 10854 12738 10906
rect 12790 10854 12802 10906
rect 12854 10854 12866 10906
rect 12918 10854 17610 10906
rect 17662 10854 17674 10906
rect 17726 10854 17738 10906
rect 17790 10854 17802 10906
rect 17854 10854 17866 10906
rect 17918 10854 22610 10906
rect 22662 10854 22674 10906
rect 22726 10854 22738 10906
rect 22790 10854 22802 10906
rect 22854 10854 22866 10906
rect 22918 10854 27610 10906
rect 27662 10854 27674 10906
rect 27726 10854 27738 10906
rect 27790 10854 27802 10906
rect 27854 10854 27866 10906
rect 27918 10854 32610 10906
rect 32662 10854 32674 10906
rect 32726 10854 32738 10906
rect 32790 10854 32802 10906
rect 32854 10854 32866 10906
rect 32918 10854 37610 10906
rect 37662 10854 37674 10906
rect 37726 10854 37738 10906
rect 37790 10854 37802 10906
rect 37854 10854 37866 10906
rect 37918 10854 40848 10906
rect 1104 10832 40848 10854
rect 33778 10792 33784 10804
rect 6886 10764 33784 10792
rect 5445 10659 5503 10665
rect 5445 10625 5457 10659
rect 5491 10656 5503 10659
rect 5721 10659 5779 10665
rect 5721 10656 5733 10659
rect 5491 10628 5733 10656
rect 5491 10625 5503 10628
rect 5445 10619 5503 10625
rect 5721 10625 5733 10628
rect 5767 10656 5779 10659
rect 6886 10656 6914 10764
rect 33778 10752 33784 10764
rect 33836 10752 33842 10804
rect 24673 10727 24731 10733
rect 24673 10693 24685 10727
rect 24719 10724 24731 10727
rect 36354 10724 36360 10736
rect 24719 10696 36360 10724
rect 24719 10693 24731 10696
rect 24673 10687 24731 10693
rect 36354 10684 36360 10696
rect 36412 10684 36418 10736
rect 5767 10628 6914 10656
rect 32953 10659 33011 10665
rect 5767 10625 5779 10628
rect 5721 10619 5779 10625
rect 32953 10625 32965 10659
rect 32999 10656 33011 10659
rect 33134 10656 33140 10668
rect 32999 10628 33140 10656
rect 32999 10625 33011 10628
rect 32953 10619 33011 10625
rect 33134 10616 33140 10628
rect 33192 10616 33198 10668
rect 33597 10659 33655 10665
rect 33597 10625 33609 10659
rect 33643 10656 33655 10659
rect 36446 10656 36452 10668
rect 33643 10628 36452 10656
rect 33643 10625 33655 10628
rect 33597 10619 33655 10625
rect 36446 10616 36452 10628
rect 36504 10616 36510 10668
rect 3142 10548 3148 10600
rect 3200 10588 3206 10600
rect 32125 10591 32183 10597
rect 32125 10588 32137 10591
rect 3200 10560 32137 10588
rect 3200 10548 3206 10560
rect 32125 10557 32137 10560
rect 32171 10557 32183 10591
rect 32125 10551 32183 10557
rect 5905 10523 5963 10529
rect 5905 10489 5917 10523
rect 5951 10520 5963 10523
rect 22370 10520 22376 10532
rect 5951 10492 22376 10520
rect 5951 10489 5963 10492
rect 5905 10483 5963 10489
rect 22370 10480 22376 10492
rect 22428 10480 22434 10532
rect 24857 10523 24915 10529
rect 24857 10489 24869 10523
rect 24903 10520 24915 10523
rect 38378 10520 38384 10532
rect 24903 10492 38384 10520
rect 24903 10489 24915 10492
rect 24857 10483 24915 10489
rect 38378 10480 38384 10492
rect 38436 10480 38442 10532
rect 1104 10362 40848 10384
rect 1104 10310 1950 10362
rect 2002 10310 2014 10362
rect 2066 10310 2078 10362
rect 2130 10310 2142 10362
rect 2194 10310 2206 10362
rect 2258 10310 6950 10362
rect 7002 10310 7014 10362
rect 7066 10310 7078 10362
rect 7130 10310 7142 10362
rect 7194 10310 7206 10362
rect 7258 10310 11950 10362
rect 12002 10310 12014 10362
rect 12066 10310 12078 10362
rect 12130 10310 12142 10362
rect 12194 10310 12206 10362
rect 12258 10310 16950 10362
rect 17002 10310 17014 10362
rect 17066 10310 17078 10362
rect 17130 10310 17142 10362
rect 17194 10310 17206 10362
rect 17258 10310 21950 10362
rect 22002 10310 22014 10362
rect 22066 10310 22078 10362
rect 22130 10310 22142 10362
rect 22194 10310 22206 10362
rect 22258 10310 26950 10362
rect 27002 10310 27014 10362
rect 27066 10310 27078 10362
rect 27130 10310 27142 10362
rect 27194 10310 27206 10362
rect 27258 10310 31950 10362
rect 32002 10310 32014 10362
rect 32066 10310 32078 10362
rect 32130 10310 32142 10362
rect 32194 10310 32206 10362
rect 32258 10310 36950 10362
rect 37002 10310 37014 10362
rect 37066 10310 37078 10362
rect 37130 10310 37142 10362
rect 37194 10310 37206 10362
rect 37258 10310 40848 10362
rect 1104 10288 40848 10310
rect 1104 9818 40848 9840
rect 1104 9766 2610 9818
rect 2662 9766 2674 9818
rect 2726 9766 2738 9818
rect 2790 9766 2802 9818
rect 2854 9766 2866 9818
rect 2918 9766 7610 9818
rect 7662 9766 7674 9818
rect 7726 9766 7738 9818
rect 7790 9766 7802 9818
rect 7854 9766 7866 9818
rect 7918 9766 12610 9818
rect 12662 9766 12674 9818
rect 12726 9766 12738 9818
rect 12790 9766 12802 9818
rect 12854 9766 12866 9818
rect 12918 9766 17610 9818
rect 17662 9766 17674 9818
rect 17726 9766 17738 9818
rect 17790 9766 17802 9818
rect 17854 9766 17866 9818
rect 17918 9766 22610 9818
rect 22662 9766 22674 9818
rect 22726 9766 22738 9818
rect 22790 9766 22802 9818
rect 22854 9766 22866 9818
rect 22918 9766 27610 9818
rect 27662 9766 27674 9818
rect 27726 9766 27738 9818
rect 27790 9766 27802 9818
rect 27854 9766 27866 9818
rect 27918 9766 32610 9818
rect 32662 9766 32674 9818
rect 32726 9766 32738 9818
rect 32790 9766 32802 9818
rect 32854 9766 32866 9818
rect 32918 9766 37610 9818
rect 37662 9766 37674 9818
rect 37726 9766 37738 9818
rect 37790 9766 37802 9818
rect 37854 9766 37866 9818
rect 37918 9766 40848 9818
rect 1104 9744 40848 9766
rect 7009 9639 7067 9645
rect 7009 9605 7021 9639
rect 7055 9636 7067 9639
rect 7558 9636 7564 9648
rect 7055 9608 7564 9636
rect 7055 9605 7067 9608
rect 7009 9599 7067 9605
rect 7558 9596 7564 9608
rect 7616 9596 7622 9648
rect 17310 9636 17316 9648
rect 8786 9608 17316 9636
rect 17310 9596 17316 9608
rect 17368 9596 17374 9648
rect 19518 9596 19524 9648
rect 19576 9636 19582 9648
rect 19978 9636 19984 9648
rect 19576 9608 19984 9636
rect 19576 9596 19582 9608
rect 19978 9596 19984 9608
rect 20036 9596 20042 9648
rect 9309 9571 9367 9577
rect 9309 9537 9321 9571
rect 9355 9568 9367 9571
rect 10410 9568 10416 9580
rect 9355 9540 10416 9568
rect 9355 9537 9367 9540
rect 9309 9531 9367 9537
rect 10410 9528 10416 9540
rect 10468 9528 10474 9580
rect 13722 9528 13728 9580
rect 13780 9568 13786 9580
rect 14553 9571 14611 9577
rect 14553 9568 14565 9571
rect 13780 9540 14565 9568
rect 13780 9528 13786 9540
rect 14553 9537 14565 9540
rect 14599 9568 14611 9571
rect 19536 9568 19564 9596
rect 14599 9540 19564 9568
rect 14599 9537 14611 9540
rect 14553 9531 14611 9537
rect 7285 9503 7343 9509
rect 7285 9469 7297 9503
rect 7331 9469 7343 9503
rect 7285 9463 7343 9469
rect 7300 9364 7328 9463
rect 9582 9364 9588 9376
rect 7300 9336 9588 9364
rect 9582 9324 9588 9336
rect 9640 9324 9646 9376
rect 14645 9367 14703 9373
rect 14645 9333 14657 9367
rect 14691 9364 14703 9367
rect 38838 9364 38844 9376
rect 14691 9336 38844 9364
rect 14691 9333 14703 9336
rect 14645 9327 14703 9333
rect 38838 9324 38844 9336
rect 38896 9324 38902 9376
rect 1104 9274 40848 9296
rect 1104 9222 1950 9274
rect 2002 9222 2014 9274
rect 2066 9222 2078 9274
rect 2130 9222 2142 9274
rect 2194 9222 2206 9274
rect 2258 9222 6950 9274
rect 7002 9222 7014 9274
rect 7066 9222 7078 9274
rect 7130 9222 7142 9274
rect 7194 9222 7206 9274
rect 7258 9222 11950 9274
rect 12002 9222 12014 9274
rect 12066 9222 12078 9274
rect 12130 9222 12142 9274
rect 12194 9222 12206 9274
rect 12258 9222 16950 9274
rect 17002 9222 17014 9274
rect 17066 9222 17078 9274
rect 17130 9222 17142 9274
rect 17194 9222 17206 9274
rect 17258 9222 21950 9274
rect 22002 9222 22014 9274
rect 22066 9222 22078 9274
rect 22130 9222 22142 9274
rect 22194 9222 22206 9274
rect 22258 9222 26950 9274
rect 27002 9222 27014 9274
rect 27066 9222 27078 9274
rect 27130 9222 27142 9274
rect 27194 9222 27206 9274
rect 27258 9222 31950 9274
rect 32002 9222 32014 9274
rect 32066 9222 32078 9274
rect 32130 9222 32142 9274
rect 32194 9222 32206 9274
rect 32258 9222 36950 9274
rect 37002 9222 37014 9274
rect 37066 9222 37078 9274
rect 37130 9222 37142 9274
rect 37194 9222 37206 9274
rect 37258 9222 40848 9274
rect 1104 9200 40848 9222
rect 7377 9163 7435 9169
rect 7377 9129 7389 9163
rect 7423 9160 7435 9163
rect 7558 9160 7564 9172
rect 7423 9132 7564 9160
rect 7423 9129 7435 9132
rect 7377 9123 7435 9129
rect 7558 9120 7564 9132
rect 7616 9120 7622 9172
rect 22462 9120 22468 9172
rect 22520 9160 22526 9172
rect 22741 9163 22799 9169
rect 22741 9160 22753 9163
rect 22520 9132 22753 9160
rect 22520 9120 22526 9132
rect 22741 9129 22753 9132
rect 22787 9129 22799 9163
rect 22741 9123 22799 9129
rect 33226 9120 33232 9172
rect 33284 9160 33290 9172
rect 37277 9163 37335 9169
rect 37277 9160 37289 9163
rect 33284 9132 37289 9160
rect 33284 9120 33290 9132
rect 37277 9129 37289 9132
rect 37323 9129 37335 9163
rect 37277 9123 37335 9129
rect 9306 8916 9312 8968
rect 9364 8956 9370 8968
rect 22925 8959 22983 8965
rect 22925 8956 22937 8959
rect 9364 8928 22937 8956
rect 9364 8916 9370 8928
rect 22925 8925 22937 8928
rect 22971 8925 22983 8959
rect 36909 8959 36967 8965
rect 36909 8956 36921 8959
rect 22925 8919 22983 8925
rect 26206 8928 36921 8956
rect 14090 8780 14096 8832
rect 14148 8820 14154 8832
rect 26206 8820 26234 8928
rect 36909 8925 36921 8928
rect 36955 8956 36967 8959
rect 37553 8959 37611 8965
rect 37553 8956 37565 8959
rect 36955 8928 37565 8956
rect 36955 8925 36967 8928
rect 36909 8919 36967 8925
rect 37553 8925 37565 8928
rect 37599 8956 37611 8959
rect 38010 8956 38016 8968
rect 37599 8928 38016 8956
rect 37599 8925 37611 8928
rect 37553 8919 37611 8925
rect 38010 8916 38016 8928
rect 38068 8916 38074 8968
rect 37369 8891 37427 8897
rect 37369 8857 37381 8891
rect 37415 8888 37427 8891
rect 38194 8888 38200 8900
rect 37415 8860 38200 8888
rect 37415 8857 37427 8860
rect 37369 8851 37427 8857
rect 38194 8848 38200 8860
rect 38252 8848 38258 8900
rect 14148 8792 26234 8820
rect 14148 8780 14154 8792
rect 1104 8730 40848 8752
rect 1104 8678 2610 8730
rect 2662 8678 2674 8730
rect 2726 8678 2738 8730
rect 2790 8678 2802 8730
rect 2854 8678 2866 8730
rect 2918 8678 7610 8730
rect 7662 8678 7674 8730
rect 7726 8678 7738 8730
rect 7790 8678 7802 8730
rect 7854 8678 7866 8730
rect 7918 8678 12610 8730
rect 12662 8678 12674 8730
rect 12726 8678 12738 8730
rect 12790 8678 12802 8730
rect 12854 8678 12866 8730
rect 12918 8678 17610 8730
rect 17662 8678 17674 8730
rect 17726 8678 17738 8730
rect 17790 8678 17802 8730
rect 17854 8678 17866 8730
rect 17918 8678 22610 8730
rect 22662 8678 22674 8730
rect 22726 8678 22738 8730
rect 22790 8678 22802 8730
rect 22854 8678 22866 8730
rect 22918 8678 27610 8730
rect 27662 8678 27674 8730
rect 27726 8678 27738 8730
rect 27790 8678 27802 8730
rect 27854 8678 27866 8730
rect 27918 8678 32610 8730
rect 32662 8678 32674 8730
rect 32726 8678 32738 8730
rect 32790 8678 32802 8730
rect 32854 8678 32866 8730
rect 32918 8678 37610 8730
rect 37662 8678 37674 8730
rect 37726 8678 37738 8730
rect 37790 8678 37802 8730
rect 37854 8678 37866 8730
rect 37918 8678 40848 8730
rect 1104 8656 40848 8678
rect 1104 8186 40848 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 6950 8186
rect 7002 8134 7014 8186
rect 7066 8134 7078 8186
rect 7130 8134 7142 8186
rect 7194 8134 7206 8186
rect 7258 8134 11950 8186
rect 12002 8134 12014 8186
rect 12066 8134 12078 8186
rect 12130 8134 12142 8186
rect 12194 8134 12206 8186
rect 12258 8134 16950 8186
rect 17002 8134 17014 8186
rect 17066 8134 17078 8186
rect 17130 8134 17142 8186
rect 17194 8134 17206 8186
rect 17258 8134 21950 8186
rect 22002 8134 22014 8186
rect 22066 8134 22078 8186
rect 22130 8134 22142 8186
rect 22194 8134 22206 8186
rect 22258 8134 26950 8186
rect 27002 8134 27014 8186
rect 27066 8134 27078 8186
rect 27130 8134 27142 8186
rect 27194 8134 27206 8186
rect 27258 8134 31950 8186
rect 32002 8134 32014 8186
rect 32066 8134 32078 8186
rect 32130 8134 32142 8186
rect 32194 8134 32206 8186
rect 32258 8134 36950 8186
rect 37002 8134 37014 8186
rect 37066 8134 37078 8186
rect 37130 8134 37142 8186
rect 37194 8134 37206 8186
rect 37258 8134 40848 8186
rect 1104 8112 40848 8134
rect 9033 8075 9091 8081
rect 9033 8041 9045 8075
rect 9079 8072 9091 8075
rect 9490 8072 9496 8084
rect 9079 8044 9496 8072
rect 9079 8041 9091 8044
rect 9033 8035 9091 8041
rect 9490 8032 9496 8044
rect 9548 8032 9554 8084
rect 13630 8032 13636 8084
rect 13688 8072 13694 8084
rect 18693 8075 18751 8081
rect 18693 8072 18705 8075
rect 13688 8044 18705 8072
rect 13688 8032 13694 8044
rect 18693 8041 18705 8044
rect 18739 8041 18751 8075
rect 18693 8035 18751 8041
rect 8941 7871 8999 7877
rect 8941 7837 8953 7871
rect 8987 7868 8999 7871
rect 13722 7868 13728 7880
rect 8987 7840 13728 7868
rect 8987 7837 8999 7840
rect 8941 7831 8999 7837
rect 13722 7828 13728 7840
rect 13780 7828 13786 7880
rect 18417 7871 18475 7877
rect 18417 7837 18429 7871
rect 18463 7868 18475 7871
rect 18874 7868 18880 7880
rect 18463 7840 18880 7868
rect 18463 7837 18475 7840
rect 18417 7831 18475 7837
rect 18874 7828 18880 7840
rect 18932 7828 18938 7880
rect 1104 7642 40848 7664
rect 1104 7590 2610 7642
rect 2662 7590 2674 7642
rect 2726 7590 2738 7642
rect 2790 7590 2802 7642
rect 2854 7590 2866 7642
rect 2918 7590 7610 7642
rect 7662 7590 7674 7642
rect 7726 7590 7738 7642
rect 7790 7590 7802 7642
rect 7854 7590 7866 7642
rect 7918 7590 12610 7642
rect 12662 7590 12674 7642
rect 12726 7590 12738 7642
rect 12790 7590 12802 7642
rect 12854 7590 12866 7642
rect 12918 7590 17610 7642
rect 17662 7590 17674 7642
rect 17726 7590 17738 7642
rect 17790 7590 17802 7642
rect 17854 7590 17866 7642
rect 17918 7590 22610 7642
rect 22662 7590 22674 7642
rect 22726 7590 22738 7642
rect 22790 7590 22802 7642
rect 22854 7590 22866 7642
rect 22918 7590 27610 7642
rect 27662 7590 27674 7642
rect 27726 7590 27738 7642
rect 27790 7590 27802 7642
rect 27854 7590 27866 7642
rect 27918 7590 32610 7642
rect 32662 7590 32674 7642
rect 32726 7590 32738 7642
rect 32790 7590 32802 7642
rect 32854 7590 32866 7642
rect 32918 7590 37610 7642
rect 37662 7590 37674 7642
rect 37726 7590 37738 7642
rect 37790 7590 37802 7642
rect 37854 7590 37866 7642
rect 37918 7590 40848 7642
rect 1104 7568 40848 7590
rect 1104 7098 40848 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 6950 7098
rect 7002 7046 7014 7098
rect 7066 7046 7078 7098
rect 7130 7046 7142 7098
rect 7194 7046 7206 7098
rect 7258 7046 11950 7098
rect 12002 7046 12014 7098
rect 12066 7046 12078 7098
rect 12130 7046 12142 7098
rect 12194 7046 12206 7098
rect 12258 7046 16950 7098
rect 17002 7046 17014 7098
rect 17066 7046 17078 7098
rect 17130 7046 17142 7098
rect 17194 7046 17206 7098
rect 17258 7046 21950 7098
rect 22002 7046 22014 7098
rect 22066 7046 22078 7098
rect 22130 7046 22142 7098
rect 22194 7046 22206 7098
rect 22258 7046 26950 7098
rect 27002 7046 27014 7098
rect 27066 7046 27078 7098
rect 27130 7046 27142 7098
rect 27194 7046 27206 7098
rect 27258 7046 31950 7098
rect 32002 7046 32014 7098
rect 32066 7046 32078 7098
rect 32130 7046 32142 7098
rect 32194 7046 32206 7098
rect 32258 7046 36950 7098
rect 37002 7046 37014 7098
rect 37066 7046 37078 7098
rect 37130 7046 37142 7098
rect 37194 7046 37206 7098
rect 37258 7046 40848 7098
rect 1104 7024 40848 7046
rect 1104 6554 40848 6576
rect 1104 6502 2610 6554
rect 2662 6502 2674 6554
rect 2726 6502 2738 6554
rect 2790 6502 2802 6554
rect 2854 6502 2866 6554
rect 2918 6502 7610 6554
rect 7662 6502 7674 6554
rect 7726 6502 7738 6554
rect 7790 6502 7802 6554
rect 7854 6502 7866 6554
rect 7918 6502 12610 6554
rect 12662 6502 12674 6554
rect 12726 6502 12738 6554
rect 12790 6502 12802 6554
rect 12854 6502 12866 6554
rect 12918 6502 17610 6554
rect 17662 6502 17674 6554
rect 17726 6502 17738 6554
rect 17790 6502 17802 6554
rect 17854 6502 17866 6554
rect 17918 6502 22610 6554
rect 22662 6502 22674 6554
rect 22726 6502 22738 6554
rect 22790 6502 22802 6554
rect 22854 6502 22866 6554
rect 22918 6502 27610 6554
rect 27662 6502 27674 6554
rect 27726 6502 27738 6554
rect 27790 6502 27802 6554
rect 27854 6502 27866 6554
rect 27918 6502 32610 6554
rect 32662 6502 32674 6554
rect 32726 6502 32738 6554
rect 32790 6502 32802 6554
rect 32854 6502 32866 6554
rect 32918 6502 37610 6554
rect 37662 6502 37674 6554
rect 37726 6502 37738 6554
rect 37790 6502 37802 6554
rect 37854 6502 37866 6554
rect 37918 6502 40848 6554
rect 1104 6480 40848 6502
rect 1104 6010 40848 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 6950 6010
rect 7002 5958 7014 6010
rect 7066 5958 7078 6010
rect 7130 5958 7142 6010
rect 7194 5958 7206 6010
rect 7258 5958 11950 6010
rect 12002 5958 12014 6010
rect 12066 5958 12078 6010
rect 12130 5958 12142 6010
rect 12194 5958 12206 6010
rect 12258 5958 16950 6010
rect 17002 5958 17014 6010
rect 17066 5958 17078 6010
rect 17130 5958 17142 6010
rect 17194 5958 17206 6010
rect 17258 5958 21950 6010
rect 22002 5958 22014 6010
rect 22066 5958 22078 6010
rect 22130 5958 22142 6010
rect 22194 5958 22206 6010
rect 22258 5958 26950 6010
rect 27002 5958 27014 6010
rect 27066 5958 27078 6010
rect 27130 5958 27142 6010
rect 27194 5958 27206 6010
rect 27258 5958 31950 6010
rect 32002 5958 32014 6010
rect 32066 5958 32078 6010
rect 32130 5958 32142 6010
rect 32194 5958 32206 6010
rect 32258 5958 36950 6010
rect 37002 5958 37014 6010
rect 37066 5958 37078 6010
rect 37130 5958 37142 6010
rect 37194 5958 37206 6010
rect 37258 5958 40848 6010
rect 1104 5936 40848 5958
rect 1104 5466 40848 5488
rect 1104 5414 2610 5466
rect 2662 5414 2674 5466
rect 2726 5414 2738 5466
rect 2790 5414 2802 5466
rect 2854 5414 2866 5466
rect 2918 5414 7610 5466
rect 7662 5414 7674 5466
rect 7726 5414 7738 5466
rect 7790 5414 7802 5466
rect 7854 5414 7866 5466
rect 7918 5414 12610 5466
rect 12662 5414 12674 5466
rect 12726 5414 12738 5466
rect 12790 5414 12802 5466
rect 12854 5414 12866 5466
rect 12918 5414 17610 5466
rect 17662 5414 17674 5466
rect 17726 5414 17738 5466
rect 17790 5414 17802 5466
rect 17854 5414 17866 5466
rect 17918 5414 22610 5466
rect 22662 5414 22674 5466
rect 22726 5414 22738 5466
rect 22790 5414 22802 5466
rect 22854 5414 22866 5466
rect 22918 5414 27610 5466
rect 27662 5414 27674 5466
rect 27726 5414 27738 5466
rect 27790 5414 27802 5466
rect 27854 5414 27866 5466
rect 27918 5414 32610 5466
rect 32662 5414 32674 5466
rect 32726 5414 32738 5466
rect 32790 5414 32802 5466
rect 32854 5414 32866 5466
rect 32918 5414 37610 5466
rect 37662 5414 37674 5466
rect 37726 5414 37738 5466
rect 37790 5414 37802 5466
rect 37854 5414 37866 5466
rect 37918 5414 40848 5466
rect 1104 5392 40848 5414
rect 19978 5176 19984 5228
rect 20036 5216 20042 5228
rect 21177 5219 21235 5225
rect 21177 5216 21189 5219
rect 20036 5188 21189 5216
rect 20036 5176 20042 5188
rect 21177 5185 21189 5188
rect 21223 5185 21235 5219
rect 21177 5179 21235 5185
rect 6086 4972 6092 5024
rect 6144 5012 6150 5024
rect 21085 5015 21143 5021
rect 21085 5012 21097 5015
rect 6144 4984 21097 5012
rect 6144 4972 6150 4984
rect 21085 4981 21097 4984
rect 21131 4981 21143 5015
rect 21085 4975 21143 4981
rect 1104 4922 40848 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 6950 4922
rect 7002 4870 7014 4922
rect 7066 4870 7078 4922
rect 7130 4870 7142 4922
rect 7194 4870 7206 4922
rect 7258 4870 11950 4922
rect 12002 4870 12014 4922
rect 12066 4870 12078 4922
rect 12130 4870 12142 4922
rect 12194 4870 12206 4922
rect 12258 4870 16950 4922
rect 17002 4870 17014 4922
rect 17066 4870 17078 4922
rect 17130 4870 17142 4922
rect 17194 4870 17206 4922
rect 17258 4870 21950 4922
rect 22002 4870 22014 4922
rect 22066 4870 22078 4922
rect 22130 4870 22142 4922
rect 22194 4870 22206 4922
rect 22258 4870 26950 4922
rect 27002 4870 27014 4922
rect 27066 4870 27078 4922
rect 27130 4870 27142 4922
rect 27194 4870 27206 4922
rect 27258 4870 31950 4922
rect 32002 4870 32014 4922
rect 32066 4870 32078 4922
rect 32130 4870 32142 4922
rect 32194 4870 32206 4922
rect 32258 4870 36950 4922
rect 37002 4870 37014 4922
rect 37066 4870 37078 4922
rect 37130 4870 37142 4922
rect 37194 4870 37206 4922
rect 37258 4870 40848 4922
rect 1104 4848 40848 4870
rect 25593 4811 25651 4817
rect 25593 4777 25605 4811
rect 25639 4777 25651 4811
rect 25593 4771 25651 4777
rect 25608 4740 25636 4771
rect 26050 4768 26056 4820
rect 26108 4768 26114 4820
rect 28902 4740 28908 4752
rect 25608 4712 28908 4740
rect 28902 4700 28908 4712
rect 28960 4700 28966 4752
rect 15838 4672 15844 4684
rect 1872 4644 15844 4672
rect 1872 4613 1900 4644
rect 15838 4632 15844 4644
rect 15896 4632 15902 4684
rect 1857 4607 1915 4613
rect 1857 4573 1869 4607
rect 1903 4573 1915 4607
rect 1857 4567 1915 4573
rect 6270 4564 6276 4616
rect 6328 4564 6334 4616
rect 25774 4564 25780 4616
rect 25832 4564 25838 4616
rect 1765 4539 1823 4545
rect 1765 4505 1777 4539
rect 1811 4536 1823 4539
rect 1811 4508 6914 4536
rect 1811 4505 1823 4508
rect 1765 4499 1823 4505
rect 6178 4428 6184 4480
rect 6236 4428 6242 4480
rect 6886 4468 6914 4508
rect 23750 4496 23756 4548
rect 23808 4536 23814 4548
rect 25869 4539 25927 4545
rect 25869 4536 25881 4539
rect 23808 4508 25881 4536
rect 23808 4496 23814 4508
rect 25869 4505 25881 4508
rect 25915 4505 25927 4539
rect 25869 4499 25927 4505
rect 38746 4468 38752 4480
rect 6886 4440 38752 4468
rect 38746 4428 38752 4440
rect 38804 4428 38810 4480
rect 1104 4378 40848 4400
rect 1104 4326 2610 4378
rect 2662 4326 2674 4378
rect 2726 4326 2738 4378
rect 2790 4326 2802 4378
rect 2854 4326 2866 4378
rect 2918 4326 7610 4378
rect 7662 4326 7674 4378
rect 7726 4326 7738 4378
rect 7790 4326 7802 4378
rect 7854 4326 7866 4378
rect 7918 4326 12610 4378
rect 12662 4326 12674 4378
rect 12726 4326 12738 4378
rect 12790 4326 12802 4378
rect 12854 4326 12866 4378
rect 12918 4326 17610 4378
rect 17662 4326 17674 4378
rect 17726 4326 17738 4378
rect 17790 4326 17802 4378
rect 17854 4326 17866 4378
rect 17918 4326 22610 4378
rect 22662 4326 22674 4378
rect 22726 4326 22738 4378
rect 22790 4326 22802 4378
rect 22854 4326 22866 4378
rect 22918 4326 27610 4378
rect 27662 4326 27674 4378
rect 27726 4326 27738 4378
rect 27790 4326 27802 4378
rect 27854 4326 27866 4378
rect 27918 4326 32610 4378
rect 32662 4326 32674 4378
rect 32726 4326 32738 4378
rect 32790 4326 32802 4378
rect 32854 4326 32866 4378
rect 32918 4326 37610 4378
rect 37662 4326 37674 4378
rect 37726 4326 37738 4378
rect 37790 4326 37802 4378
rect 37854 4326 37866 4378
rect 37918 4326 40848 4378
rect 1104 4304 40848 4326
rect 2498 3952 2504 4004
rect 2556 3992 2562 4004
rect 14274 3992 14280 4004
rect 2556 3964 14280 3992
rect 2556 3952 2562 3964
rect 14274 3952 14280 3964
rect 14332 3952 14338 4004
rect 2866 3884 2872 3936
rect 2924 3924 2930 3936
rect 12342 3924 12348 3936
rect 2924 3896 12348 3924
rect 2924 3884 2930 3896
rect 12342 3884 12348 3896
rect 12400 3884 12406 3936
rect 1104 3834 40848 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 6950 3834
rect 7002 3782 7014 3834
rect 7066 3782 7078 3834
rect 7130 3782 7142 3834
rect 7194 3782 7206 3834
rect 7258 3782 11950 3834
rect 12002 3782 12014 3834
rect 12066 3782 12078 3834
rect 12130 3782 12142 3834
rect 12194 3782 12206 3834
rect 12258 3782 16950 3834
rect 17002 3782 17014 3834
rect 17066 3782 17078 3834
rect 17130 3782 17142 3834
rect 17194 3782 17206 3834
rect 17258 3782 21950 3834
rect 22002 3782 22014 3834
rect 22066 3782 22078 3834
rect 22130 3782 22142 3834
rect 22194 3782 22206 3834
rect 22258 3782 26950 3834
rect 27002 3782 27014 3834
rect 27066 3782 27078 3834
rect 27130 3782 27142 3834
rect 27194 3782 27206 3834
rect 27258 3782 31950 3834
rect 32002 3782 32014 3834
rect 32066 3782 32078 3834
rect 32130 3782 32142 3834
rect 32194 3782 32206 3834
rect 32258 3782 36950 3834
rect 37002 3782 37014 3834
rect 37066 3782 37078 3834
rect 37130 3782 37142 3834
rect 37194 3782 37206 3834
rect 37258 3782 40848 3834
rect 1104 3760 40848 3782
rect 8478 3680 8484 3732
rect 8536 3720 8542 3732
rect 29454 3720 29460 3732
rect 8536 3692 29460 3720
rect 8536 3680 8542 3692
rect 29454 3680 29460 3692
rect 29512 3680 29518 3732
rect 3050 3612 3056 3664
rect 3108 3612 3114 3664
rect 7101 3655 7159 3661
rect 7101 3652 7113 3655
rect 6886 3624 7113 3652
rect 1670 3544 1676 3596
rect 1728 3544 1734 3596
rect 6886 3584 6914 3624
rect 7101 3621 7113 3624
rect 7147 3652 7159 3655
rect 13906 3652 13912 3664
rect 7147 3624 13912 3652
rect 7147 3621 7159 3624
rect 7101 3615 7159 3621
rect 13906 3612 13912 3624
rect 13964 3612 13970 3664
rect 2990 3556 6914 3584
rect 2225 3519 2283 3525
rect 2225 3485 2237 3519
rect 2271 3485 2283 3519
rect 2225 3479 2283 3485
rect 2240 3448 2268 3479
rect 2866 3476 2872 3528
rect 2924 3476 2930 3528
rect 7193 3519 7251 3525
rect 7193 3485 7205 3519
rect 7239 3516 7251 3519
rect 7374 3516 7380 3528
rect 7239 3488 7380 3516
rect 7239 3485 7251 3488
rect 7193 3479 7251 3485
rect 7374 3476 7380 3488
rect 7432 3476 7438 3528
rect 6178 3448 6184 3460
rect 2240 3420 6184 3448
rect 6178 3408 6184 3420
rect 6236 3408 6242 3460
rect 6362 3340 6368 3392
rect 6420 3380 6426 3392
rect 7006 3380 7012 3392
rect 6420 3352 7012 3380
rect 6420 3340 6426 3352
rect 7006 3340 7012 3352
rect 7064 3340 7070 3392
rect 9490 3340 9496 3392
rect 9548 3380 9554 3392
rect 14366 3380 14372 3392
rect 9548 3352 14372 3380
rect 9548 3340 9554 3352
rect 14366 3340 14372 3352
rect 14424 3340 14430 3392
rect 1104 3290 40848 3312
rect 1104 3238 2610 3290
rect 2662 3238 2674 3290
rect 2726 3238 2738 3290
rect 2790 3238 2802 3290
rect 2854 3238 2866 3290
rect 2918 3238 7610 3290
rect 7662 3238 7674 3290
rect 7726 3238 7738 3290
rect 7790 3238 7802 3290
rect 7854 3238 7866 3290
rect 7918 3238 12610 3290
rect 12662 3238 12674 3290
rect 12726 3238 12738 3290
rect 12790 3238 12802 3290
rect 12854 3238 12866 3290
rect 12918 3238 17610 3290
rect 17662 3238 17674 3290
rect 17726 3238 17738 3290
rect 17790 3238 17802 3290
rect 17854 3238 17866 3290
rect 17918 3238 22610 3290
rect 22662 3238 22674 3290
rect 22726 3238 22738 3290
rect 22790 3238 22802 3290
rect 22854 3238 22866 3290
rect 22918 3238 27610 3290
rect 27662 3238 27674 3290
rect 27726 3238 27738 3290
rect 27790 3238 27802 3290
rect 27854 3238 27866 3290
rect 27918 3238 32610 3290
rect 32662 3238 32674 3290
rect 32726 3238 32738 3290
rect 32790 3238 32802 3290
rect 32854 3238 32866 3290
rect 32918 3238 37610 3290
rect 37662 3238 37674 3290
rect 37726 3238 37738 3290
rect 37790 3238 37802 3290
rect 37854 3238 37866 3290
rect 37918 3238 40848 3290
rect 1104 3216 40848 3238
rect 4706 3136 4712 3188
rect 4764 3176 4770 3188
rect 14829 3179 14887 3185
rect 14829 3176 14841 3179
rect 4764 3148 14841 3176
rect 4764 3136 4770 3148
rect 14829 3145 14841 3148
rect 14875 3145 14887 3179
rect 14829 3139 14887 3145
rect 7006 3068 7012 3120
rect 7064 3108 7070 3120
rect 14645 3111 14703 3117
rect 14645 3108 14657 3111
rect 7064 3080 14657 3108
rect 7064 3068 7070 3080
rect 14645 3077 14657 3080
rect 14691 3077 14703 3111
rect 14645 3071 14703 3077
rect 7282 3000 7288 3052
rect 7340 3040 7346 3052
rect 7561 3043 7619 3049
rect 7561 3040 7573 3043
rect 7340 3012 7573 3040
rect 7340 3000 7346 3012
rect 7561 3009 7573 3012
rect 7607 3009 7619 3043
rect 7561 3003 7619 3009
rect 8110 3000 8116 3052
rect 8168 3000 8174 3052
rect 8478 3000 8484 3052
rect 8536 3000 8542 3052
rect 8754 3000 8760 3052
rect 8812 3000 8818 3052
rect 9033 3043 9091 3049
rect 9033 3009 9045 3043
rect 9079 3040 9091 3043
rect 9079 3012 9444 3040
rect 9079 3009 9091 3012
rect 9033 3003 9091 3009
rect 8294 2932 8300 2984
rect 8352 2932 8358 2984
rect 9416 2904 9444 3012
rect 9490 3000 9496 3052
rect 9548 3000 9554 3052
rect 9861 3043 9919 3049
rect 9861 3009 9873 3043
rect 9907 3009 9919 3043
rect 9861 3003 9919 3009
rect 10137 3043 10195 3049
rect 10137 3009 10149 3043
rect 10183 3040 10195 3043
rect 14090 3040 14096 3052
rect 10183 3012 14096 3040
rect 10183 3009 10195 3012
rect 10137 3003 10195 3009
rect 9766 2932 9772 2984
rect 9824 2932 9830 2984
rect 9876 2972 9904 3003
rect 14090 3000 14096 3012
rect 14148 3000 14154 3052
rect 14274 3000 14280 3052
rect 14332 3000 14338 3052
rect 21818 3040 21824 3052
rect 16546 3012 21824 3040
rect 14182 2972 14188 2984
rect 9876 2944 14188 2972
rect 14182 2932 14188 2944
rect 14240 2932 14246 2984
rect 16546 2904 16574 3012
rect 21818 3000 21824 3012
rect 21876 3000 21882 3052
rect 29178 3000 29184 3052
rect 29236 3040 29242 3052
rect 30653 3043 30711 3049
rect 30653 3040 30665 3043
rect 29236 3012 30665 3040
rect 29236 3000 29242 3012
rect 30653 3009 30665 3012
rect 30699 3009 30711 3043
rect 30653 3003 30711 3009
rect 30929 3043 30987 3049
rect 30929 3009 30941 3043
rect 30975 3040 30987 3043
rect 38286 3040 38292 3052
rect 30975 3012 38292 3040
rect 30975 3009 30987 3012
rect 30929 3003 30987 3009
rect 38286 3000 38292 3012
rect 38344 3000 38350 3052
rect 9416 2876 16574 2904
rect 14274 2796 14280 2848
rect 14332 2836 14338 2848
rect 14829 2839 14887 2845
rect 14829 2836 14841 2839
rect 14332 2808 14841 2836
rect 14332 2796 14338 2808
rect 14829 2805 14841 2808
rect 14875 2805 14887 2839
rect 14829 2799 14887 2805
rect 15013 2839 15071 2845
rect 15013 2805 15025 2839
rect 15059 2836 15071 2839
rect 21634 2836 21640 2848
rect 15059 2808 21640 2836
rect 15059 2805 15071 2808
rect 15013 2799 15071 2805
rect 21634 2796 21640 2808
rect 21692 2796 21698 2848
rect 1104 2746 40848 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 6950 2746
rect 7002 2694 7014 2746
rect 7066 2694 7078 2746
rect 7130 2694 7142 2746
rect 7194 2694 7206 2746
rect 7258 2694 11950 2746
rect 12002 2694 12014 2746
rect 12066 2694 12078 2746
rect 12130 2694 12142 2746
rect 12194 2694 12206 2746
rect 12258 2694 16950 2746
rect 17002 2694 17014 2746
rect 17066 2694 17078 2746
rect 17130 2694 17142 2746
rect 17194 2694 17206 2746
rect 17258 2694 21950 2746
rect 22002 2694 22014 2746
rect 22066 2694 22078 2746
rect 22130 2694 22142 2746
rect 22194 2694 22206 2746
rect 22258 2694 26950 2746
rect 27002 2694 27014 2746
rect 27066 2694 27078 2746
rect 27130 2694 27142 2746
rect 27194 2694 27206 2746
rect 27258 2694 31950 2746
rect 32002 2694 32014 2746
rect 32066 2694 32078 2746
rect 32130 2694 32142 2746
rect 32194 2694 32206 2746
rect 32258 2694 36950 2746
rect 37002 2694 37014 2746
rect 37066 2694 37078 2746
rect 37130 2694 37142 2746
rect 37194 2694 37206 2746
rect 37258 2694 40848 2746
rect 1104 2672 40848 2694
rect 36630 2592 36636 2644
rect 36688 2632 36694 2644
rect 36817 2635 36875 2641
rect 36817 2632 36829 2635
rect 36688 2604 36829 2632
rect 36688 2592 36694 2604
rect 36817 2601 36829 2604
rect 36863 2601 36875 2635
rect 36817 2595 36875 2601
rect 15194 2524 15200 2576
rect 15252 2564 15258 2576
rect 39393 2567 39451 2573
rect 39393 2564 39405 2567
rect 15252 2536 39405 2564
rect 15252 2524 15258 2536
rect 39393 2533 39405 2536
rect 39439 2533 39451 2567
rect 39393 2527 39451 2533
rect 18598 2456 18604 2508
rect 18656 2496 18662 2508
rect 30834 2496 30840 2508
rect 18656 2468 30840 2496
rect 18656 2456 18662 2468
rect 30834 2456 30840 2468
rect 30892 2456 30898 2508
rect 30944 2468 36952 2496
rect 2498 2388 2504 2440
rect 2556 2428 2562 2440
rect 2685 2431 2743 2437
rect 2685 2428 2697 2431
rect 2556 2400 2697 2428
rect 2556 2388 2562 2400
rect 2685 2397 2697 2400
rect 2731 2397 2743 2431
rect 2685 2391 2743 2397
rect 9122 2388 9128 2440
rect 9180 2428 9186 2440
rect 30944 2428 30972 2468
rect 9180 2400 30972 2428
rect 9180 2388 9186 2400
rect 31110 2388 31116 2440
rect 31168 2428 31174 2440
rect 36924 2437 36952 2468
rect 36725 2431 36783 2437
rect 36725 2428 36737 2431
rect 31168 2400 36737 2428
rect 31168 2388 31174 2400
rect 36725 2397 36737 2400
rect 36771 2397 36783 2431
rect 36725 2391 36783 2397
rect 36909 2431 36967 2437
rect 36909 2397 36921 2431
rect 36955 2397 36967 2431
rect 36909 2391 36967 2397
rect 39298 2388 39304 2440
rect 39356 2428 39362 2440
rect 39853 2431 39911 2437
rect 39853 2428 39865 2431
rect 39356 2400 39865 2428
rect 39356 2388 39362 2400
rect 39853 2397 39865 2400
rect 39899 2397 39911 2431
rect 39853 2391 39911 2397
rect 10226 2320 10232 2372
rect 10284 2360 10290 2372
rect 39209 2363 39267 2369
rect 39209 2360 39221 2363
rect 10284 2332 35894 2360
rect 10284 2320 10290 2332
rect 7929 2295 7987 2301
rect 7929 2261 7941 2295
rect 7975 2292 7987 2295
rect 8018 2292 8024 2304
rect 7975 2264 8024 2292
rect 7975 2261 7987 2264
rect 7929 2255 7987 2261
rect 8018 2252 8024 2264
rect 8076 2252 8082 2304
rect 13078 2252 13084 2304
rect 13136 2292 13142 2304
rect 13173 2295 13231 2301
rect 13173 2292 13185 2295
rect 13136 2264 13185 2292
rect 13136 2252 13142 2264
rect 13173 2261 13185 2264
rect 13219 2261 13231 2295
rect 13173 2255 13231 2261
rect 18322 2252 18328 2304
rect 18380 2292 18386 2304
rect 18417 2295 18475 2301
rect 18417 2292 18429 2295
rect 18380 2264 18429 2292
rect 18380 2252 18386 2264
rect 18417 2261 18429 2264
rect 18463 2261 18475 2295
rect 18417 2255 18475 2261
rect 23566 2252 23572 2304
rect 23624 2292 23630 2304
rect 23661 2295 23719 2301
rect 23661 2292 23673 2295
rect 23624 2264 23673 2292
rect 23624 2252 23630 2264
rect 23661 2261 23673 2264
rect 23707 2261 23719 2295
rect 23661 2255 23719 2261
rect 28810 2252 28816 2304
rect 28868 2292 28874 2304
rect 28905 2295 28963 2301
rect 28905 2292 28917 2295
rect 28868 2264 28917 2292
rect 28868 2252 28874 2264
rect 28905 2261 28917 2264
rect 28951 2261 28963 2295
rect 28905 2255 28963 2261
rect 34054 2252 34060 2304
rect 34112 2292 34118 2304
rect 34149 2295 34207 2301
rect 34149 2292 34161 2295
rect 34112 2264 34161 2292
rect 34112 2252 34118 2264
rect 34149 2261 34161 2264
rect 34195 2261 34207 2295
rect 35866 2292 35894 2332
rect 38764 2332 39221 2360
rect 38764 2301 38792 2332
rect 39209 2329 39221 2332
rect 39255 2329 39267 2363
rect 39209 2323 39267 2329
rect 38749 2295 38807 2301
rect 38749 2292 38761 2295
rect 35866 2264 38761 2292
rect 34149 2255 34207 2261
rect 38749 2261 38761 2264
rect 38795 2261 38807 2295
rect 38749 2255 38807 2261
rect 1104 2202 40848 2224
rect 1104 2150 2610 2202
rect 2662 2150 2674 2202
rect 2726 2150 2738 2202
rect 2790 2150 2802 2202
rect 2854 2150 2866 2202
rect 2918 2150 7610 2202
rect 7662 2150 7674 2202
rect 7726 2150 7738 2202
rect 7790 2150 7802 2202
rect 7854 2150 7866 2202
rect 7918 2150 12610 2202
rect 12662 2150 12674 2202
rect 12726 2150 12738 2202
rect 12790 2150 12802 2202
rect 12854 2150 12866 2202
rect 12918 2150 17610 2202
rect 17662 2150 17674 2202
rect 17726 2150 17738 2202
rect 17790 2150 17802 2202
rect 17854 2150 17866 2202
rect 17918 2150 22610 2202
rect 22662 2150 22674 2202
rect 22726 2150 22738 2202
rect 22790 2150 22802 2202
rect 22854 2150 22866 2202
rect 22918 2150 27610 2202
rect 27662 2150 27674 2202
rect 27726 2150 27738 2202
rect 27790 2150 27802 2202
rect 27854 2150 27866 2202
rect 27918 2150 32610 2202
rect 32662 2150 32674 2202
rect 32726 2150 32738 2202
rect 32790 2150 32802 2202
rect 32854 2150 32866 2202
rect 32918 2150 37610 2202
rect 37662 2150 37674 2202
rect 37726 2150 37738 2202
rect 37790 2150 37802 2202
rect 37854 2150 37866 2202
rect 37918 2150 40848 2202
rect 1104 2128 40848 2150
<< via1 >>
rect 2610 69606 2662 69658
rect 2674 69606 2726 69658
rect 2738 69606 2790 69658
rect 2802 69606 2854 69658
rect 2866 69606 2918 69658
rect 7610 69606 7662 69658
rect 7674 69606 7726 69658
rect 7738 69606 7790 69658
rect 7802 69606 7854 69658
rect 7866 69606 7918 69658
rect 12610 69606 12662 69658
rect 12674 69606 12726 69658
rect 12738 69606 12790 69658
rect 12802 69606 12854 69658
rect 12866 69606 12918 69658
rect 17610 69606 17662 69658
rect 17674 69606 17726 69658
rect 17738 69606 17790 69658
rect 17802 69606 17854 69658
rect 17866 69606 17918 69658
rect 22610 69606 22662 69658
rect 22674 69606 22726 69658
rect 22738 69606 22790 69658
rect 22802 69606 22854 69658
rect 22866 69606 22918 69658
rect 27610 69606 27662 69658
rect 27674 69606 27726 69658
rect 27738 69606 27790 69658
rect 27802 69606 27854 69658
rect 27866 69606 27918 69658
rect 32610 69606 32662 69658
rect 32674 69606 32726 69658
rect 32738 69606 32790 69658
rect 32802 69606 32854 69658
rect 32866 69606 32918 69658
rect 37610 69606 37662 69658
rect 37674 69606 37726 69658
rect 37738 69606 37790 69658
rect 37802 69606 37854 69658
rect 37866 69606 37918 69658
rect 3056 69547 3108 69556
rect 3056 69513 3065 69547
rect 3065 69513 3099 69547
rect 3099 69513 3108 69547
rect 3056 69504 3108 69513
rect 8944 69504 8996 69556
rect 15016 69547 15068 69556
rect 15016 69513 15025 69547
rect 15025 69513 15059 69547
rect 15059 69513 15068 69547
rect 15016 69504 15068 69513
rect 20996 69547 21048 69556
rect 20996 69513 21005 69547
rect 21005 69513 21039 69547
rect 21039 69513 21048 69547
rect 20996 69504 21048 69513
rect 26976 69547 27028 69556
rect 26976 69513 26985 69547
rect 26985 69513 27019 69547
rect 27019 69513 27028 69547
rect 26976 69504 27028 69513
rect 32956 69547 33008 69556
rect 32956 69513 32965 69547
rect 32965 69513 32999 69547
rect 32999 69513 33008 69547
rect 32956 69504 33008 69513
rect 38936 69547 38988 69556
rect 38936 69513 38945 69547
rect 38945 69513 38979 69547
rect 38979 69513 38988 69547
rect 38936 69504 38988 69513
rect 3332 69368 3384 69420
rect 9220 69411 9272 69420
rect 9220 69377 9229 69411
rect 9229 69377 9263 69411
rect 9263 69377 9272 69411
rect 9220 69368 9272 69377
rect 15200 69411 15252 69420
rect 15200 69377 15209 69411
rect 15209 69377 15243 69411
rect 15243 69377 15252 69411
rect 15200 69368 15252 69377
rect 21180 69411 21232 69420
rect 21180 69377 21189 69411
rect 21189 69377 21223 69411
rect 21223 69377 21232 69411
rect 21180 69368 21232 69377
rect 27344 69368 27396 69420
rect 33140 69411 33192 69420
rect 33140 69377 33149 69411
rect 33149 69377 33183 69411
rect 33183 69377 33192 69411
rect 33140 69368 33192 69377
rect 39120 69411 39172 69420
rect 39120 69377 39129 69411
rect 39129 69377 39163 69411
rect 39163 69377 39172 69411
rect 39120 69368 39172 69377
rect 1950 69062 2002 69114
rect 2014 69062 2066 69114
rect 2078 69062 2130 69114
rect 2142 69062 2194 69114
rect 2206 69062 2258 69114
rect 6950 69062 7002 69114
rect 7014 69062 7066 69114
rect 7078 69062 7130 69114
rect 7142 69062 7194 69114
rect 7206 69062 7258 69114
rect 11950 69062 12002 69114
rect 12014 69062 12066 69114
rect 12078 69062 12130 69114
rect 12142 69062 12194 69114
rect 12206 69062 12258 69114
rect 16950 69062 17002 69114
rect 17014 69062 17066 69114
rect 17078 69062 17130 69114
rect 17142 69062 17194 69114
rect 17206 69062 17258 69114
rect 21950 69062 22002 69114
rect 22014 69062 22066 69114
rect 22078 69062 22130 69114
rect 22142 69062 22194 69114
rect 22206 69062 22258 69114
rect 26950 69062 27002 69114
rect 27014 69062 27066 69114
rect 27078 69062 27130 69114
rect 27142 69062 27194 69114
rect 27206 69062 27258 69114
rect 31950 69062 32002 69114
rect 32014 69062 32066 69114
rect 32078 69062 32130 69114
rect 32142 69062 32194 69114
rect 32206 69062 32258 69114
rect 36950 69062 37002 69114
rect 37014 69062 37066 69114
rect 37078 69062 37130 69114
rect 37142 69062 37194 69114
rect 37206 69062 37258 69114
rect 36176 68824 36228 68876
rect 16488 68688 16540 68740
rect 35992 68731 36044 68740
rect 35992 68697 36001 68731
rect 36001 68697 36035 68731
rect 36035 68697 36044 68731
rect 35992 68688 36044 68697
rect 16672 68620 16724 68672
rect 36544 68620 36596 68672
rect 36636 68663 36688 68672
rect 36636 68629 36645 68663
rect 36645 68629 36679 68663
rect 36679 68629 36688 68663
rect 36636 68620 36688 68629
rect 37372 68620 37424 68672
rect 2610 68518 2662 68570
rect 2674 68518 2726 68570
rect 2738 68518 2790 68570
rect 2802 68518 2854 68570
rect 2866 68518 2918 68570
rect 7610 68518 7662 68570
rect 7674 68518 7726 68570
rect 7738 68518 7790 68570
rect 7802 68518 7854 68570
rect 7866 68518 7918 68570
rect 12610 68518 12662 68570
rect 12674 68518 12726 68570
rect 12738 68518 12790 68570
rect 12802 68518 12854 68570
rect 12866 68518 12918 68570
rect 17610 68518 17662 68570
rect 17674 68518 17726 68570
rect 17738 68518 17790 68570
rect 17802 68518 17854 68570
rect 17866 68518 17918 68570
rect 22610 68518 22662 68570
rect 22674 68518 22726 68570
rect 22738 68518 22790 68570
rect 22802 68518 22854 68570
rect 22866 68518 22918 68570
rect 27610 68518 27662 68570
rect 27674 68518 27726 68570
rect 27738 68518 27790 68570
rect 27802 68518 27854 68570
rect 27866 68518 27918 68570
rect 32610 68518 32662 68570
rect 32674 68518 32726 68570
rect 32738 68518 32790 68570
rect 32802 68518 32854 68570
rect 32866 68518 32918 68570
rect 37610 68518 37662 68570
rect 37674 68518 37726 68570
rect 37738 68518 37790 68570
rect 37802 68518 37854 68570
rect 37866 68518 37918 68570
rect 6828 68323 6880 68332
rect 6828 68289 6837 68323
rect 6837 68289 6871 68323
rect 6871 68289 6880 68323
rect 6828 68280 6880 68289
rect 7288 68323 7340 68332
rect 7288 68289 7297 68323
rect 7297 68289 7331 68323
rect 7331 68289 7340 68323
rect 7288 68280 7340 68289
rect 9128 68391 9180 68400
rect 9128 68357 9137 68391
rect 9137 68357 9171 68391
rect 9171 68357 9180 68391
rect 9128 68348 9180 68357
rect 18696 68348 18748 68400
rect 29092 68348 29144 68400
rect 32404 68323 32456 68332
rect 32404 68289 32413 68323
rect 32413 68289 32447 68323
rect 32447 68289 32456 68323
rect 32404 68280 32456 68289
rect 31852 68212 31904 68264
rect 34152 68212 34204 68264
rect 9036 68076 9088 68128
rect 9588 68144 9640 68196
rect 9312 68119 9364 68128
rect 9312 68085 9321 68119
rect 9321 68085 9355 68119
rect 9355 68085 9364 68119
rect 9312 68076 9364 68085
rect 1950 67974 2002 68026
rect 2014 67974 2066 68026
rect 2078 67974 2130 68026
rect 2142 67974 2194 68026
rect 2206 67974 2258 68026
rect 6950 67974 7002 68026
rect 7014 67974 7066 68026
rect 7078 67974 7130 68026
rect 7142 67974 7194 68026
rect 7206 67974 7258 68026
rect 11950 67974 12002 68026
rect 12014 67974 12066 68026
rect 12078 67974 12130 68026
rect 12142 67974 12194 68026
rect 12206 67974 12258 68026
rect 16950 67974 17002 68026
rect 17014 67974 17066 68026
rect 17078 67974 17130 68026
rect 17142 67974 17194 68026
rect 17206 67974 17258 68026
rect 21950 67974 22002 68026
rect 22014 67974 22066 68026
rect 22078 67974 22130 68026
rect 22142 67974 22194 68026
rect 22206 67974 22258 68026
rect 26950 67974 27002 68026
rect 27014 67974 27066 68026
rect 27078 67974 27130 68026
rect 27142 67974 27194 68026
rect 27206 67974 27258 68026
rect 31950 67974 32002 68026
rect 32014 67974 32066 68026
rect 32078 67974 32130 68026
rect 32142 67974 32194 68026
rect 32206 67974 32258 68026
rect 36950 67974 37002 68026
rect 37014 67974 37066 68026
rect 37078 67974 37130 68026
rect 37142 67974 37194 68026
rect 37206 67974 37258 68026
rect 2504 67804 2556 67856
rect 2320 67668 2372 67720
rect 7472 67668 7524 67720
rect 37464 67736 37516 67788
rect 29920 67668 29972 67720
rect 6368 67643 6420 67652
rect 6368 67609 6377 67643
rect 6377 67609 6411 67643
rect 6411 67609 6420 67643
rect 6368 67600 6420 67609
rect 24860 67643 24912 67652
rect 24860 67609 24869 67643
rect 24869 67609 24903 67643
rect 24903 67609 24912 67643
rect 24860 67600 24912 67609
rect 25044 67643 25096 67652
rect 25044 67609 25053 67643
rect 25053 67609 25087 67643
rect 25087 67609 25096 67643
rect 25044 67600 25096 67609
rect 34152 67643 34204 67652
rect 34152 67609 34161 67643
rect 34161 67609 34195 67643
rect 34195 67609 34204 67643
rect 34152 67600 34204 67609
rect 34520 67643 34572 67652
rect 34520 67609 34529 67643
rect 34529 67609 34563 67643
rect 34563 67609 34572 67643
rect 34520 67600 34572 67609
rect 2610 67430 2662 67482
rect 2674 67430 2726 67482
rect 2738 67430 2790 67482
rect 2802 67430 2854 67482
rect 2866 67430 2918 67482
rect 7610 67430 7662 67482
rect 7674 67430 7726 67482
rect 7738 67430 7790 67482
rect 7802 67430 7854 67482
rect 7866 67430 7918 67482
rect 12610 67430 12662 67482
rect 12674 67430 12726 67482
rect 12738 67430 12790 67482
rect 12802 67430 12854 67482
rect 12866 67430 12918 67482
rect 17610 67430 17662 67482
rect 17674 67430 17726 67482
rect 17738 67430 17790 67482
rect 17802 67430 17854 67482
rect 17866 67430 17918 67482
rect 22610 67430 22662 67482
rect 22674 67430 22726 67482
rect 22738 67430 22790 67482
rect 22802 67430 22854 67482
rect 22866 67430 22918 67482
rect 27610 67430 27662 67482
rect 27674 67430 27726 67482
rect 27738 67430 27790 67482
rect 27802 67430 27854 67482
rect 27866 67430 27918 67482
rect 32610 67430 32662 67482
rect 32674 67430 32726 67482
rect 32738 67430 32790 67482
rect 32802 67430 32854 67482
rect 32866 67430 32918 67482
rect 37610 67430 37662 67482
rect 37674 67430 37726 67482
rect 37738 67430 37790 67482
rect 37802 67430 37854 67482
rect 37866 67430 37918 67482
rect 14280 67235 14332 67244
rect 14280 67201 14289 67235
rect 14289 67201 14323 67235
rect 14323 67201 14332 67235
rect 14280 67192 14332 67201
rect 14188 67167 14240 67176
rect 14188 67133 14197 67167
rect 14197 67133 14231 67167
rect 14231 67133 14240 67167
rect 14188 67124 14240 67133
rect 15016 67167 15068 67176
rect 15016 67133 15025 67167
rect 15025 67133 15059 67167
rect 15059 67133 15068 67167
rect 15016 67124 15068 67133
rect 17316 67124 17368 67176
rect 1950 66886 2002 66938
rect 2014 66886 2066 66938
rect 2078 66886 2130 66938
rect 2142 66886 2194 66938
rect 2206 66886 2258 66938
rect 6950 66886 7002 66938
rect 7014 66886 7066 66938
rect 7078 66886 7130 66938
rect 7142 66886 7194 66938
rect 7206 66886 7258 66938
rect 11950 66886 12002 66938
rect 12014 66886 12066 66938
rect 12078 66886 12130 66938
rect 12142 66886 12194 66938
rect 12206 66886 12258 66938
rect 16950 66886 17002 66938
rect 17014 66886 17066 66938
rect 17078 66886 17130 66938
rect 17142 66886 17194 66938
rect 17206 66886 17258 66938
rect 21950 66886 22002 66938
rect 22014 66886 22066 66938
rect 22078 66886 22130 66938
rect 22142 66886 22194 66938
rect 22206 66886 22258 66938
rect 26950 66886 27002 66938
rect 27014 66886 27066 66938
rect 27078 66886 27130 66938
rect 27142 66886 27194 66938
rect 27206 66886 27258 66938
rect 31950 66886 32002 66938
rect 32014 66886 32066 66938
rect 32078 66886 32130 66938
rect 32142 66886 32194 66938
rect 32206 66886 32258 66938
rect 36950 66886 37002 66938
rect 37014 66886 37066 66938
rect 37078 66886 37130 66938
rect 37142 66886 37194 66938
rect 37206 66886 37258 66938
rect 6460 66623 6512 66632
rect 6460 66589 6469 66623
rect 6469 66589 6503 66623
rect 6503 66589 6512 66623
rect 6460 66580 6512 66589
rect 6644 66487 6696 66496
rect 6644 66453 6653 66487
rect 6653 66453 6687 66487
rect 6687 66453 6696 66487
rect 6644 66444 6696 66453
rect 2610 66342 2662 66394
rect 2674 66342 2726 66394
rect 2738 66342 2790 66394
rect 2802 66342 2854 66394
rect 2866 66342 2918 66394
rect 7610 66342 7662 66394
rect 7674 66342 7726 66394
rect 7738 66342 7790 66394
rect 7802 66342 7854 66394
rect 7866 66342 7918 66394
rect 12610 66342 12662 66394
rect 12674 66342 12726 66394
rect 12738 66342 12790 66394
rect 12802 66342 12854 66394
rect 12866 66342 12918 66394
rect 17610 66342 17662 66394
rect 17674 66342 17726 66394
rect 17738 66342 17790 66394
rect 17802 66342 17854 66394
rect 17866 66342 17918 66394
rect 22610 66342 22662 66394
rect 22674 66342 22726 66394
rect 22738 66342 22790 66394
rect 22802 66342 22854 66394
rect 22866 66342 22918 66394
rect 27610 66342 27662 66394
rect 27674 66342 27726 66394
rect 27738 66342 27790 66394
rect 27802 66342 27854 66394
rect 27866 66342 27918 66394
rect 32610 66342 32662 66394
rect 32674 66342 32726 66394
rect 32738 66342 32790 66394
rect 32802 66342 32854 66394
rect 32866 66342 32918 66394
rect 37610 66342 37662 66394
rect 37674 66342 37726 66394
rect 37738 66342 37790 66394
rect 37802 66342 37854 66394
rect 37866 66342 37918 66394
rect 3608 66104 3660 66156
rect 9128 66104 9180 66156
rect 24216 66104 24268 66156
rect 25504 65968 25556 66020
rect 1950 65798 2002 65850
rect 2014 65798 2066 65850
rect 2078 65798 2130 65850
rect 2142 65798 2194 65850
rect 2206 65798 2258 65850
rect 6950 65798 7002 65850
rect 7014 65798 7066 65850
rect 7078 65798 7130 65850
rect 7142 65798 7194 65850
rect 7206 65798 7258 65850
rect 11950 65798 12002 65850
rect 12014 65798 12066 65850
rect 12078 65798 12130 65850
rect 12142 65798 12194 65850
rect 12206 65798 12258 65850
rect 16950 65798 17002 65850
rect 17014 65798 17066 65850
rect 17078 65798 17130 65850
rect 17142 65798 17194 65850
rect 17206 65798 17258 65850
rect 21950 65798 22002 65850
rect 22014 65798 22066 65850
rect 22078 65798 22130 65850
rect 22142 65798 22194 65850
rect 22206 65798 22258 65850
rect 26950 65798 27002 65850
rect 27014 65798 27066 65850
rect 27078 65798 27130 65850
rect 27142 65798 27194 65850
rect 27206 65798 27258 65850
rect 31950 65798 32002 65850
rect 32014 65798 32066 65850
rect 32078 65798 32130 65850
rect 32142 65798 32194 65850
rect 32206 65798 32258 65850
rect 36950 65798 37002 65850
rect 37014 65798 37066 65850
rect 37078 65798 37130 65850
rect 37142 65798 37194 65850
rect 37206 65798 37258 65850
rect 6460 65739 6512 65748
rect 6460 65705 6469 65739
rect 6469 65705 6503 65739
rect 6503 65705 6512 65739
rect 6460 65696 6512 65705
rect 2610 65254 2662 65306
rect 2674 65254 2726 65306
rect 2738 65254 2790 65306
rect 2802 65254 2854 65306
rect 2866 65254 2918 65306
rect 7610 65254 7662 65306
rect 7674 65254 7726 65306
rect 7738 65254 7790 65306
rect 7802 65254 7854 65306
rect 7866 65254 7918 65306
rect 12610 65254 12662 65306
rect 12674 65254 12726 65306
rect 12738 65254 12790 65306
rect 12802 65254 12854 65306
rect 12866 65254 12918 65306
rect 17610 65254 17662 65306
rect 17674 65254 17726 65306
rect 17738 65254 17790 65306
rect 17802 65254 17854 65306
rect 17866 65254 17918 65306
rect 22610 65254 22662 65306
rect 22674 65254 22726 65306
rect 22738 65254 22790 65306
rect 22802 65254 22854 65306
rect 22866 65254 22918 65306
rect 27610 65254 27662 65306
rect 27674 65254 27726 65306
rect 27738 65254 27790 65306
rect 27802 65254 27854 65306
rect 27866 65254 27918 65306
rect 32610 65254 32662 65306
rect 32674 65254 32726 65306
rect 32738 65254 32790 65306
rect 32802 65254 32854 65306
rect 32866 65254 32918 65306
rect 37610 65254 37662 65306
rect 37674 65254 37726 65306
rect 37738 65254 37790 65306
rect 37802 65254 37854 65306
rect 37866 65254 37918 65306
rect 17408 65084 17460 65136
rect 23112 65084 23164 65136
rect 10692 64991 10744 65000
rect 10692 64957 10701 64991
rect 10701 64957 10735 64991
rect 10735 64957 10744 64991
rect 10692 64948 10744 64957
rect 10784 64991 10836 65000
rect 10784 64957 10793 64991
rect 10793 64957 10827 64991
rect 10827 64957 10836 64991
rect 10784 64948 10836 64957
rect 10968 64991 11020 65000
rect 10968 64957 10977 64991
rect 10977 64957 11011 64991
rect 11011 64957 11020 64991
rect 10968 64948 11020 64957
rect 23020 65016 23072 65068
rect 2412 64923 2464 64932
rect 2412 64889 2421 64923
rect 2421 64889 2455 64923
rect 2455 64889 2464 64923
rect 2412 64880 2464 64889
rect 22376 64880 22428 64932
rect 23296 64948 23348 65000
rect 35440 64948 35492 65000
rect 26700 64880 26752 64932
rect 1950 64710 2002 64762
rect 2014 64710 2066 64762
rect 2078 64710 2130 64762
rect 2142 64710 2194 64762
rect 2206 64710 2258 64762
rect 6950 64710 7002 64762
rect 7014 64710 7066 64762
rect 7078 64710 7130 64762
rect 7142 64710 7194 64762
rect 7206 64710 7258 64762
rect 11950 64710 12002 64762
rect 12014 64710 12066 64762
rect 12078 64710 12130 64762
rect 12142 64710 12194 64762
rect 12206 64710 12258 64762
rect 16950 64710 17002 64762
rect 17014 64710 17066 64762
rect 17078 64710 17130 64762
rect 17142 64710 17194 64762
rect 17206 64710 17258 64762
rect 21950 64710 22002 64762
rect 22014 64710 22066 64762
rect 22078 64710 22130 64762
rect 22142 64710 22194 64762
rect 22206 64710 22258 64762
rect 26950 64710 27002 64762
rect 27014 64710 27066 64762
rect 27078 64710 27130 64762
rect 27142 64710 27194 64762
rect 27206 64710 27258 64762
rect 31950 64710 32002 64762
rect 32014 64710 32066 64762
rect 32078 64710 32130 64762
rect 32142 64710 32194 64762
rect 32206 64710 32258 64762
rect 36950 64710 37002 64762
rect 37014 64710 37066 64762
rect 37078 64710 37130 64762
rect 37142 64710 37194 64762
rect 37206 64710 37258 64762
rect 11060 64447 11112 64456
rect 11060 64413 11069 64447
rect 11069 64413 11103 64447
rect 11103 64413 11112 64447
rect 11060 64404 11112 64413
rect 17500 64472 17552 64524
rect 12348 64404 12400 64456
rect 15016 64404 15068 64456
rect 16488 64379 16540 64388
rect 16488 64345 16497 64379
rect 16497 64345 16531 64379
rect 16531 64345 16540 64379
rect 16488 64336 16540 64345
rect 16672 64404 16724 64456
rect 11796 64311 11848 64320
rect 11796 64277 11805 64311
rect 11805 64277 11839 64311
rect 11839 64277 11848 64311
rect 11796 64268 11848 64277
rect 16580 64268 16632 64320
rect 16764 64311 16816 64320
rect 16764 64277 16773 64311
rect 16773 64277 16807 64311
rect 16807 64277 16816 64311
rect 16764 64268 16816 64277
rect 19892 64268 19944 64320
rect 24860 64268 24912 64320
rect 26700 64379 26752 64388
rect 26700 64345 26709 64379
rect 26709 64345 26743 64379
rect 26743 64345 26752 64379
rect 26700 64336 26752 64345
rect 27528 64268 27580 64320
rect 2610 64166 2662 64218
rect 2674 64166 2726 64218
rect 2738 64166 2790 64218
rect 2802 64166 2854 64218
rect 2866 64166 2918 64218
rect 7610 64166 7662 64218
rect 7674 64166 7726 64218
rect 7738 64166 7790 64218
rect 7802 64166 7854 64218
rect 7866 64166 7918 64218
rect 12610 64166 12662 64218
rect 12674 64166 12726 64218
rect 12738 64166 12790 64218
rect 12802 64166 12854 64218
rect 12866 64166 12918 64218
rect 17610 64166 17662 64218
rect 17674 64166 17726 64218
rect 17738 64166 17790 64218
rect 17802 64166 17854 64218
rect 17866 64166 17918 64218
rect 22610 64166 22662 64218
rect 22674 64166 22726 64218
rect 22738 64166 22790 64218
rect 22802 64166 22854 64218
rect 22866 64166 22918 64218
rect 27610 64166 27662 64218
rect 27674 64166 27726 64218
rect 27738 64166 27790 64218
rect 27802 64166 27854 64218
rect 27866 64166 27918 64218
rect 32610 64166 32662 64218
rect 32674 64166 32726 64218
rect 32738 64166 32790 64218
rect 32802 64166 32854 64218
rect 32866 64166 32918 64218
rect 37610 64166 37662 64218
rect 37674 64166 37726 64218
rect 37738 64166 37790 64218
rect 37802 64166 37854 64218
rect 37866 64166 37918 64218
rect 16580 64064 16632 64116
rect 36544 64064 36596 64116
rect 5724 63928 5776 63980
rect 14372 63928 14424 63980
rect 15660 63928 15712 63980
rect 18972 63996 19024 64048
rect 18604 63971 18656 63980
rect 18604 63937 18613 63971
rect 18613 63937 18647 63971
rect 18647 63937 18656 63971
rect 18604 63928 18656 63937
rect 18696 63928 18748 63980
rect 21824 63928 21876 63980
rect 27436 63860 27488 63912
rect 14096 63724 14148 63776
rect 15292 63767 15344 63776
rect 15292 63733 15301 63767
rect 15301 63733 15335 63767
rect 15335 63733 15344 63767
rect 15292 63724 15344 63733
rect 18512 63724 18564 63776
rect 20720 63724 20772 63776
rect 32496 63724 32548 63776
rect 1950 63622 2002 63674
rect 2014 63622 2066 63674
rect 2078 63622 2130 63674
rect 2142 63622 2194 63674
rect 2206 63622 2258 63674
rect 6950 63622 7002 63674
rect 7014 63622 7066 63674
rect 7078 63622 7130 63674
rect 7142 63622 7194 63674
rect 7206 63622 7258 63674
rect 11950 63622 12002 63674
rect 12014 63622 12066 63674
rect 12078 63622 12130 63674
rect 12142 63622 12194 63674
rect 12206 63622 12258 63674
rect 16950 63622 17002 63674
rect 17014 63622 17066 63674
rect 17078 63622 17130 63674
rect 17142 63622 17194 63674
rect 17206 63622 17258 63674
rect 21950 63622 22002 63674
rect 22014 63622 22066 63674
rect 22078 63622 22130 63674
rect 22142 63622 22194 63674
rect 22206 63622 22258 63674
rect 26950 63622 27002 63674
rect 27014 63622 27066 63674
rect 27078 63622 27130 63674
rect 27142 63622 27194 63674
rect 27206 63622 27258 63674
rect 31950 63622 32002 63674
rect 32014 63622 32066 63674
rect 32078 63622 32130 63674
rect 32142 63622 32194 63674
rect 32206 63622 32258 63674
rect 36950 63622 37002 63674
rect 37014 63622 37066 63674
rect 37078 63622 37130 63674
rect 37142 63622 37194 63674
rect 37206 63622 37258 63674
rect 4068 63520 4120 63572
rect 24860 63520 24912 63572
rect 25136 63520 25188 63572
rect 17408 63452 17460 63504
rect 3608 63316 3660 63368
rect 20352 63359 20404 63368
rect 20352 63325 20361 63359
rect 20361 63325 20395 63359
rect 20395 63325 20404 63359
rect 20352 63316 20404 63325
rect 33232 63316 33284 63368
rect 24216 63180 24268 63232
rect 2610 63078 2662 63130
rect 2674 63078 2726 63130
rect 2738 63078 2790 63130
rect 2802 63078 2854 63130
rect 2866 63078 2918 63130
rect 7610 63078 7662 63130
rect 7674 63078 7726 63130
rect 7738 63078 7790 63130
rect 7802 63078 7854 63130
rect 7866 63078 7918 63130
rect 12610 63078 12662 63130
rect 12674 63078 12726 63130
rect 12738 63078 12790 63130
rect 12802 63078 12854 63130
rect 12866 63078 12918 63130
rect 17610 63078 17662 63130
rect 17674 63078 17726 63130
rect 17738 63078 17790 63130
rect 17802 63078 17854 63130
rect 17866 63078 17918 63130
rect 22610 63078 22662 63130
rect 22674 63078 22726 63130
rect 22738 63078 22790 63130
rect 22802 63078 22854 63130
rect 22866 63078 22918 63130
rect 27610 63078 27662 63130
rect 27674 63078 27726 63130
rect 27738 63078 27790 63130
rect 27802 63078 27854 63130
rect 27866 63078 27918 63130
rect 32610 63078 32662 63130
rect 32674 63078 32726 63130
rect 32738 63078 32790 63130
rect 32802 63078 32854 63130
rect 32866 63078 32918 63130
rect 37610 63078 37662 63130
rect 37674 63078 37726 63130
rect 37738 63078 37790 63130
rect 37802 63078 37854 63130
rect 37866 63078 37918 63130
rect 24860 62840 24912 62892
rect 36084 62636 36136 62688
rect 1950 62534 2002 62586
rect 2014 62534 2066 62586
rect 2078 62534 2130 62586
rect 2142 62534 2194 62586
rect 2206 62534 2258 62586
rect 6950 62534 7002 62586
rect 7014 62534 7066 62586
rect 7078 62534 7130 62586
rect 7142 62534 7194 62586
rect 7206 62534 7258 62586
rect 11950 62534 12002 62586
rect 12014 62534 12066 62586
rect 12078 62534 12130 62586
rect 12142 62534 12194 62586
rect 12206 62534 12258 62586
rect 16950 62534 17002 62586
rect 17014 62534 17066 62586
rect 17078 62534 17130 62586
rect 17142 62534 17194 62586
rect 17206 62534 17258 62586
rect 21950 62534 22002 62586
rect 22014 62534 22066 62586
rect 22078 62534 22130 62586
rect 22142 62534 22194 62586
rect 22206 62534 22258 62586
rect 26950 62534 27002 62586
rect 27014 62534 27066 62586
rect 27078 62534 27130 62586
rect 27142 62534 27194 62586
rect 27206 62534 27258 62586
rect 31950 62534 32002 62586
rect 32014 62534 32066 62586
rect 32078 62534 32130 62586
rect 32142 62534 32194 62586
rect 32206 62534 32258 62586
rect 36950 62534 37002 62586
rect 37014 62534 37066 62586
rect 37078 62534 37130 62586
rect 37142 62534 37194 62586
rect 37206 62534 37258 62586
rect 11244 62296 11296 62348
rect 36820 62228 36872 62280
rect 39764 62228 39816 62280
rect 39948 62228 40000 62280
rect 19616 62203 19668 62212
rect 19616 62169 19625 62203
rect 19625 62169 19659 62203
rect 19659 62169 19668 62203
rect 19616 62160 19668 62169
rect 39304 62160 39356 62212
rect 39488 62203 39540 62212
rect 39488 62169 39497 62203
rect 39497 62169 39531 62203
rect 39531 62169 39540 62203
rect 39488 62160 39540 62169
rect 11336 62092 11388 62144
rect 19892 62135 19944 62144
rect 19892 62101 19901 62135
rect 19901 62101 19935 62135
rect 19935 62101 19944 62135
rect 19892 62092 19944 62101
rect 24952 62092 25004 62144
rect 40408 62135 40460 62144
rect 40408 62101 40417 62135
rect 40417 62101 40451 62135
rect 40451 62101 40460 62135
rect 40408 62092 40460 62101
rect 2610 61990 2662 62042
rect 2674 61990 2726 62042
rect 2738 61990 2790 62042
rect 2802 61990 2854 62042
rect 2866 61990 2918 62042
rect 7610 61990 7662 62042
rect 7674 61990 7726 62042
rect 7738 61990 7790 62042
rect 7802 61990 7854 62042
rect 7866 61990 7918 62042
rect 12610 61990 12662 62042
rect 12674 61990 12726 62042
rect 12738 61990 12790 62042
rect 12802 61990 12854 62042
rect 12866 61990 12918 62042
rect 17610 61990 17662 62042
rect 17674 61990 17726 62042
rect 17738 61990 17790 62042
rect 17802 61990 17854 62042
rect 17866 61990 17918 62042
rect 22610 61990 22662 62042
rect 22674 61990 22726 62042
rect 22738 61990 22790 62042
rect 22802 61990 22854 62042
rect 22866 61990 22918 62042
rect 27610 61990 27662 62042
rect 27674 61990 27726 62042
rect 27738 61990 27790 62042
rect 27802 61990 27854 62042
rect 27866 61990 27918 62042
rect 32610 61990 32662 62042
rect 32674 61990 32726 62042
rect 32738 61990 32790 62042
rect 32802 61990 32854 62042
rect 32866 61990 32918 62042
rect 37610 61990 37662 62042
rect 37674 61990 37726 62042
rect 37738 61990 37790 62042
rect 37802 61990 37854 62042
rect 37866 61990 37918 62042
rect 25228 61752 25280 61804
rect 26148 61591 26200 61600
rect 26148 61557 26157 61591
rect 26157 61557 26191 61591
rect 26191 61557 26200 61591
rect 26148 61548 26200 61557
rect 1950 61446 2002 61498
rect 2014 61446 2066 61498
rect 2078 61446 2130 61498
rect 2142 61446 2194 61498
rect 2206 61446 2258 61498
rect 6950 61446 7002 61498
rect 7014 61446 7066 61498
rect 7078 61446 7130 61498
rect 7142 61446 7194 61498
rect 7206 61446 7258 61498
rect 11950 61446 12002 61498
rect 12014 61446 12066 61498
rect 12078 61446 12130 61498
rect 12142 61446 12194 61498
rect 12206 61446 12258 61498
rect 16950 61446 17002 61498
rect 17014 61446 17066 61498
rect 17078 61446 17130 61498
rect 17142 61446 17194 61498
rect 17206 61446 17258 61498
rect 21950 61446 22002 61498
rect 22014 61446 22066 61498
rect 22078 61446 22130 61498
rect 22142 61446 22194 61498
rect 22206 61446 22258 61498
rect 26950 61446 27002 61498
rect 27014 61446 27066 61498
rect 27078 61446 27130 61498
rect 27142 61446 27194 61498
rect 27206 61446 27258 61498
rect 31950 61446 32002 61498
rect 32014 61446 32066 61498
rect 32078 61446 32130 61498
rect 32142 61446 32194 61498
rect 32206 61446 32258 61498
rect 36950 61446 37002 61498
rect 37014 61446 37066 61498
rect 37078 61446 37130 61498
rect 37142 61446 37194 61498
rect 37206 61446 37258 61498
rect 2610 60902 2662 60954
rect 2674 60902 2726 60954
rect 2738 60902 2790 60954
rect 2802 60902 2854 60954
rect 2866 60902 2918 60954
rect 7610 60902 7662 60954
rect 7674 60902 7726 60954
rect 7738 60902 7790 60954
rect 7802 60902 7854 60954
rect 7866 60902 7918 60954
rect 12610 60902 12662 60954
rect 12674 60902 12726 60954
rect 12738 60902 12790 60954
rect 12802 60902 12854 60954
rect 12866 60902 12918 60954
rect 17610 60902 17662 60954
rect 17674 60902 17726 60954
rect 17738 60902 17790 60954
rect 17802 60902 17854 60954
rect 17866 60902 17918 60954
rect 22610 60902 22662 60954
rect 22674 60902 22726 60954
rect 22738 60902 22790 60954
rect 22802 60902 22854 60954
rect 22866 60902 22918 60954
rect 27610 60902 27662 60954
rect 27674 60902 27726 60954
rect 27738 60902 27790 60954
rect 27802 60902 27854 60954
rect 27866 60902 27918 60954
rect 32610 60902 32662 60954
rect 32674 60902 32726 60954
rect 32738 60902 32790 60954
rect 32802 60902 32854 60954
rect 32866 60902 32918 60954
rect 37610 60902 37662 60954
rect 37674 60902 37726 60954
rect 37738 60902 37790 60954
rect 37802 60902 37854 60954
rect 37866 60902 37918 60954
rect 1950 60358 2002 60410
rect 2014 60358 2066 60410
rect 2078 60358 2130 60410
rect 2142 60358 2194 60410
rect 2206 60358 2258 60410
rect 6950 60358 7002 60410
rect 7014 60358 7066 60410
rect 7078 60358 7130 60410
rect 7142 60358 7194 60410
rect 7206 60358 7258 60410
rect 11950 60358 12002 60410
rect 12014 60358 12066 60410
rect 12078 60358 12130 60410
rect 12142 60358 12194 60410
rect 12206 60358 12258 60410
rect 16950 60358 17002 60410
rect 17014 60358 17066 60410
rect 17078 60358 17130 60410
rect 17142 60358 17194 60410
rect 17206 60358 17258 60410
rect 21950 60358 22002 60410
rect 22014 60358 22066 60410
rect 22078 60358 22130 60410
rect 22142 60358 22194 60410
rect 22206 60358 22258 60410
rect 26950 60358 27002 60410
rect 27014 60358 27066 60410
rect 27078 60358 27130 60410
rect 27142 60358 27194 60410
rect 27206 60358 27258 60410
rect 31950 60358 32002 60410
rect 32014 60358 32066 60410
rect 32078 60358 32130 60410
rect 32142 60358 32194 60410
rect 32206 60358 32258 60410
rect 36950 60358 37002 60410
rect 37014 60358 37066 60410
rect 37078 60358 37130 60410
rect 37142 60358 37194 60410
rect 37206 60358 37258 60410
rect 38476 60256 38528 60308
rect 24860 60095 24912 60104
rect 24860 60061 24869 60095
rect 24869 60061 24903 60095
rect 24903 60061 24912 60095
rect 24860 60052 24912 60061
rect 29644 60052 29696 60104
rect 23020 59984 23072 60036
rect 23388 59984 23440 60036
rect 37464 59984 37516 60036
rect 38200 59984 38252 60036
rect 23204 59916 23256 59968
rect 38292 59916 38344 59968
rect 2610 59814 2662 59866
rect 2674 59814 2726 59866
rect 2738 59814 2790 59866
rect 2802 59814 2854 59866
rect 2866 59814 2918 59866
rect 7610 59814 7662 59866
rect 7674 59814 7726 59866
rect 7738 59814 7790 59866
rect 7802 59814 7854 59866
rect 7866 59814 7918 59866
rect 12610 59814 12662 59866
rect 12674 59814 12726 59866
rect 12738 59814 12790 59866
rect 12802 59814 12854 59866
rect 12866 59814 12918 59866
rect 17610 59814 17662 59866
rect 17674 59814 17726 59866
rect 17738 59814 17790 59866
rect 17802 59814 17854 59866
rect 17866 59814 17918 59866
rect 22610 59814 22662 59866
rect 22674 59814 22726 59866
rect 22738 59814 22790 59866
rect 22802 59814 22854 59866
rect 22866 59814 22918 59866
rect 27610 59814 27662 59866
rect 27674 59814 27726 59866
rect 27738 59814 27790 59866
rect 27802 59814 27854 59866
rect 27866 59814 27918 59866
rect 32610 59814 32662 59866
rect 32674 59814 32726 59866
rect 32738 59814 32790 59866
rect 32802 59814 32854 59866
rect 32866 59814 32918 59866
rect 37610 59814 37662 59866
rect 37674 59814 37726 59866
rect 37738 59814 37790 59866
rect 37802 59814 37854 59866
rect 37866 59814 37918 59866
rect 1950 59270 2002 59322
rect 2014 59270 2066 59322
rect 2078 59270 2130 59322
rect 2142 59270 2194 59322
rect 2206 59270 2258 59322
rect 6950 59270 7002 59322
rect 7014 59270 7066 59322
rect 7078 59270 7130 59322
rect 7142 59270 7194 59322
rect 7206 59270 7258 59322
rect 11950 59270 12002 59322
rect 12014 59270 12066 59322
rect 12078 59270 12130 59322
rect 12142 59270 12194 59322
rect 12206 59270 12258 59322
rect 16950 59270 17002 59322
rect 17014 59270 17066 59322
rect 17078 59270 17130 59322
rect 17142 59270 17194 59322
rect 17206 59270 17258 59322
rect 21950 59270 22002 59322
rect 22014 59270 22066 59322
rect 22078 59270 22130 59322
rect 22142 59270 22194 59322
rect 22206 59270 22258 59322
rect 26950 59270 27002 59322
rect 27014 59270 27066 59322
rect 27078 59270 27130 59322
rect 27142 59270 27194 59322
rect 27206 59270 27258 59322
rect 31950 59270 32002 59322
rect 32014 59270 32066 59322
rect 32078 59270 32130 59322
rect 32142 59270 32194 59322
rect 32206 59270 32258 59322
rect 36950 59270 37002 59322
rect 37014 59270 37066 59322
rect 37078 59270 37130 59322
rect 37142 59270 37194 59322
rect 37206 59270 37258 59322
rect 7472 58964 7524 59016
rect 25228 58964 25280 59016
rect 25596 58964 25648 59016
rect 8024 58828 8076 58880
rect 2610 58726 2662 58778
rect 2674 58726 2726 58778
rect 2738 58726 2790 58778
rect 2802 58726 2854 58778
rect 2866 58726 2918 58778
rect 7610 58726 7662 58778
rect 7674 58726 7726 58778
rect 7738 58726 7790 58778
rect 7802 58726 7854 58778
rect 7866 58726 7918 58778
rect 12610 58726 12662 58778
rect 12674 58726 12726 58778
rect 12738 58726 12790 58778
rect 12802 58726 12854 58778
rect 12866 58726 12918 58778
rect 17610 58726 17662 58778
rect 17674 58726 17726 58778
rect 17738 58726 17790 58778
rect 17802 58726 17854 58778
rect 17866 58726 17918 58778
rect 22610 58726 22662 58778
rect 22674 58726 22726 58778
rect 22738 58726 22790 58778
rect 22802 58726 22854 58778
rect 22866 58726 22918 58778
rect 27610 58726 27662 58778
rect 27674 58726 27726 58778
rect 27738 58726 27790 58778
rect 27802 58726 27854 58778
rect 27866 58726 27918 58778
rect 32610 58726 32662 58778
rect 32674 58726 32726 58778
rect 32738 58726 32790 58778
rect 32802 58726 32854 58778
rect 32866 58726 32918 58778
rect 37610 58726 37662 58778
rect 37674 58726 37726 58778
rect 37738 58726 37790 58778
rect 37802 58726 37854 58778
rect 37866 58726 37918 58778
rect 38936 58488 38988 58540
rect 35440 58420 35492 58472
rect 33232 58284 33284 58336
rect 1950 58182 2002 58234
rect 2014 58182 2066 58234
rect 2078 58182 2130 58234
rect 2142 58182 2194 58234
rect 2206 58182 2258 58234
rect 6950 58182 7002 58234
rect 7014 58182 7066 58234
rect 7078 58182 7130 58234
rect 7142 58182 7194 58234
rect 7206 58182 7258 58234
rect 11950 58182 12002 58234
rect 12014 58182 12066 58234
rect 12078 58182 12130 58234
rect 12142 58182 12194 58234
rect 12206 58182 12258 58234
rect 16950 58182 17002 58234
rect 17014 58182 17066 58234
rect 17078 58182 17130 58234
rect 17142 58182 17194 58234
rect 17206 58182 17258 58234
rect 21950 58182 22002 58234
rect 22014 58182 22066 58234
rect 22078 58182 22130 58234
rect 22142 58182 22194 58234
rect 22206 58182 22258 58234
rect 26950 58182 27002 58234
rect 27014 58182 27066 58234
rect 27078 58182 27130 58234
rect 27142 58182 27194 58234
rect 27206 58182 27258 58234
rect 31950 58182 32002 58234
rect 32014 58182 32066 58234
rect 32078 58182 32130 58234
rect 32142 58182 32194 58234
rect 32206 58182 32258 58234
rect 36950 58182 37002 58234
rect 37014 58182 37066 58234
rect 37078 58182 37130 58234
rect 37142 58182 37194 58234
rect 37206 58182 37258 58234
rect 10508 57876 10560 57928
rect 10784 57876 10836 57928
rect 39212 57876 39264 57928
rect 40132 57919 40184 57928
rect 40132 57885 40141 57919
rect 40141 57885 40175 57919
rect 40175 57885 40184 57919
rect 40132 57876 40184 57885
rect 3332 57808 3384 57860
rect 29828 57808 29880 57860
rect 39028 57808 39080 57860
rect 39304 57808 39356 57860
rect 29736 57740 29788 57792
rect 36820 57740 36872 57792
rect 39672 57740 39724 57792
rect 2610 57638 2662 57690
rect 2674 57638 2726 57690
rect 2738 57638 2790 57690
rect 2802 57638 2854 57690
rect 2866 57638 2918 57690
rect 7610 57638 7662 57690
rect 7674 57638 7726 57690
rect 7738 57638 7790 57690
rect 7802 57638 7854 57690
rect 7866 57638 7918 57690
rect 12610 57638 12662 57690
rect 12674 57638 12726 57690
rect 12738 57638 12790 57690
rect 12802 57638 12854 57690
rect 12866 57638 12918 57690
rect 17610 57638 17662 57690
rect 17674 57638 17726 57690
rect 17738 57638 17790 57690
rect 17802 57638 17854 57690
rect 17866 57638 17918 57690
rect 22610 57638 22662 57690
rect 22674 57638 22726 57690
rect 22738 57638 22790 57690
rect 22802 57638 22854 57690
rect 22866 57638 22918 57690
rect 27610 57638 27662 57690
rect 27674 57638 27726 57690
rect 27738 57638 27790 57690
rect 27802 57638 27854 57690
rect 27866 57638 27918 57690
rect 32610 57638 32662 57690
rect 32674 57638 32726 57690
rect 32738 57638 32790 57690
rect 32802 57638 32854 57690
rect 32866 57638 32918 57690
rect 37610 57638 37662 57690
rect 37674 57638 37726 57690
rect 37738 57638 37790 57690
rect 37802 57638 37854 57690
rect 37866 57638 37918 57690
rect 8300 57536 8352 57588
rect 29828 57579 29880 57588
rect 29828 57545 29837 57579
rect 29837 57545 29871 57579
rect 29871 57545 29880 57579
rect 29828 57536 29880 57545
rect 5724 57511 5776 57520
rect 5724 57477 5733 57511
rect 5733 57477 5767 57511
rect 5767 57477 5776 57511
rect 5724 57468 5776 57477
rect 40132 57536 40184 57588
rect 3884 57400 3936 57452
rect 5540 57443 5592 57452
rect 5540 57409 5549 57443
rect 5549 57409 5583 57443
rect 5583 57409 5592 57443
rect 5540 57400 5592 57409
rect 23112 57400 23164 57452
rect 29828 57443 29880 57452
rect 29828 57409 29837 57443
rect 29837 57409 29871 57443
rect 29871 57409 29880 57443
rect 29828 57400 29880 57409
rect 4988 57375 5040 57384
rect 4988 57341 4997 57375
rect 4997 57341 5031 57375
rect 5031 57341 5040 57375
rect 4988 57332 5040 57341
rect 5264 57375 5316 57384
rect 5264 57341 5273 57375
rect 5273 57341 5307 57375
rect 5307 57341 5316 57375
rect 5264 57332 5316 57341
rect 5356 57375 5408 57384
rect 5356 57341 5365 57375
rect 5365 57341 5399 57375
rect 5399 57341 5408 57375
rect 5356 57332 5408 57341
rect 6092 57375 6144 57384
rect 6092 57341 6101 57375
rect 6101 57341 6135 57375
rect 6135 57341 6144 57375
rect 6092 57332 6144 57341
rect 24124 57332 24176 57384
rect 29736 57375 29788 57384
rect 29736 57341 29745 57375
rect 29745 57341 29779 57375
rect 29779 57341 29788 57375
rect 29736 57332 29788 57341
rect 25780 57196 25832 57248
rect 31668 57468 31720 57520
rect 36176 57511 36228 57520
rect 36176 57477 36185 57511
rect 36185 57477 36219 57511
rect 36219 57477 36228 57511
rect 36176 57468 36228 57477
rect 36452 57443 36504 57452
rect 36452 57409 36461 57443
rect 36461 57409 36495 57443
rect 36495 57409 36504 57443
rect 36452 57400 36504 57409
rect 39948 57400 40000 57452
rect 37280 57264 37332 57316
rect 1950 57094 2002 57146
rect 2014 57094 2066 57146
rect 2078 57094 2130 57146
rect 2142 57094 2194 57146
rect 2206 57094 2258 57146
rect 6950 57094 7002 57146
rect 7014 57094 7066 57146
rect 7078 57094 7130 57146
rect 7142 57094 7194 57146
rect 7206 57094 7258 57146
rect 11950 57094 12002 57146
rect 12014 57094 12066 57146
rect 12078 57094 12130 57146
rect 12142 57094 12194 57146
rect 12206 57094 12258 57146
rect 16950 57094 17002 57146
rect 17014 57094 17066 57146
rect 17078 57094 17130 57146
rect 17142 57094 17194 57146
rect 17206 57094 17258 57146
rect 21950 57094 22002 57146
rect 22014 57094 22066 57146
rect 22078 57094 22130 57146
rect 22142 57094 22194 57146
rect 22206 57094 22258 57146
rect 26950 57094 27002 57146
rect 27014 57094 27066 57146
rect 27078 57094 27130 57146
rect 27142 57094 27194 57146
rect 27206 57094 27258 57146
rect 31950 57094 32002 57146
rect 32014 57094 32066 57146
rect 32078 57094 32130 57146
rect 32142 57094 32194 57146
rect 32206 57094 32258 57146
rect 36950 57094 37002 57146
rect 37014 57094 37066 57146
rect 37078 57094 37130 57146
rect 37142 57094 37194 57146
rect 37206 57094 37258 57146
rect 29828 56992 29880 57044
rect 39488 56992 39540 57044
rect 5264 56856 5316 56908
rect 8392 56856 8444 56908
rect 7380 56788 7432 56840
rect 10508 56788 10560 56840
rect 2504 56720 2556 56772
rect 29828 56720 29880 56772
rect 36452 56720 36504 56772
rect 8300 56652 8352 56704
rect 30564 56652 30616 56704
rect 2610 56550 2662 56602
rect 2674 56550 2726 56602
rect 2738 56550 2790 56602
rect 2802 56550 2854 56602
rect 2866 56550 2918 56602
rect 7610 56550 7662 56602
rect 7674 56550 7726 56602
rect 7738 56550 7790 56602
rect 7802 56550 7854 56602
rect 7866 56550 7918 56602
rect 12610 56550 12662 56602
rect 12674 56550 12726 56602
rect 12738 56550 12790 56602
rect 12802 56550 12854 56602
rect 12866 56550 12918 56602
rect 17610 56550 17662 56602
rect 17674 56550 17726 56602
rect 17738 56550 17790 56602
rect 17802 56550 17854 56602
rect 17866 56550 17918 56602
rect 22610 56550 22662 56602
rect 22674 56550 22726 56602
rect 22738 56550 22790 56602
rect 22802 56550 22854 56602
rect 22866 56550 22918 56602
rect 27610 56550 27662 56602
rect 27674 56550 27726 56602
rect 27738 56550 27790 56602
rect 27802 56550 27854 56602
rect 27866 56550 27918 56602
rect 32610 56550 32662 56602
rect 32674 56550 32726 56602
rect 32738 56550 32790 56602
rect 32802 56550 32854 56602
rect 32866 56550 32918 56602
rect 37610 56550 37662 56602
rect 37674 56550 37726 56602
rect 37738 56550 37790 56602
rect 37802 56550 37854 56602
rect 37866 56550 37918 56602
rect 33416 56448 33468 56500
rect 34152 56448 34204 56500
rect 28540 56380 28592 56432
rect 29000 56423 29052 56432
rect 29000 56389 29009 56423
rect 29009 56389 29043 56423
rect 29043 56389 29052 56423
rect 29000 56380 29052 56389
rect 33692 56423 33744 56432
rect 33692 56389 33701 56423
rect 33701 56389 33735 56423
rect 33735 56389 33744 56423
rect 33692 56380 33744 56389
rect 33876 56423 33928 56432
rect 33876 56389 33885 56423
rect 33885 56389 33919 56423
rect 33919 56389 33928 56423
rect 33876 56380 33928 56389
rect 37464 56380 37516 56432
rect 38844 56380 38896 56432
rect 37280 56355 37332 56364
rect 37280 56321 37289 56355
rect 37289 56321 37323 56355
rect 37323 56321 37332 56355
rect 37280 56312 37332 56321
rect 38016 56244 38068 56296
rect 38108 56244 38160 56296
rect 28540 56151 28592 56160
rect 28540 56117 28549 56151
rect 28549 56117 28583 56151
rect 28583 56117 28592 56151
rect 28540 56108 28592 56117
rect 28632 56108 28684 56160
rect 29184 56151 29236 56160
rect 29184 56117 29193 56151
rect 29193 56117 29227 56151
rect 29227 56117 29236 56151
rect 29184 56108 29236 56117
rect 33508 56151 33560 56160
rect 33508 56117 33517 56151
rect 33517 56117 33551 56151
rect 33551 56117 33560 56151
rect 33508 56108 33560 56117
rect 33600 56108 33652 56160
rect 1950 56006 2002 56058
rect 2014 56006 2066 56058
rect 2078 56006 2130 56058
rect 2142 56006 2194 56058
rect 2206 56006 2258 56058
rect 6950 56006 7002 56058
rect 7014 56006 7066 56058
rect 7078 56006 7130 56058
rect 7142 56006 7194 56058
rect 7206 56006 7258 56058
rect 11950 56006 12002 56058
rect 12014 56006 12066 56058
rect 12078 56006 12130 56058
rect 12142 56006 12194 56058
rect 12206 56006 12258 56058
rect 16950 56006 17002 56058
rect 17014 56006 17066 56058
rect 17078 56006 17130 56058
rect 17142 56006 17194 56058
rect 17206 56006 17258 56058
rect 21950 56006 22002 56058
rect 22014 56006 22066 56058
rect 22078 56006 22130 56058
rect 22142 56006 22194 56058
rect 22206 56006 22258 56058
rect 26950 56006 27002 56058
rect 27014 56006 27066 56058
rect 27078 56006 27130 56058
rect 27142 56006 27194 56058
rect 27206 56006 27258 56058
rect 31950 56006 32002 56058
rect 32014 56006 32066 56058
rect 32078 56006 32130 56058
rect 32142 56006 32194 56058
rect 32206 56006 32258 56058
rect 36950 56006 37002 56058
rect 37014 56006 37066 56058
rect 37078 56006 37130 56058
rect 37142 56006 37194 56058
rect 37206 56006 37258 56058
rect 12348 55836 12400 55888
rect 38108 55836 38160 55888
rect 21456 55768 21508 55820
rect 21824 55768 21876 55820
rect 20536 55632 20588 55684
rect 33416 55632 33468 55684
rect 28632 55564 28684 55616
rect 29644 55607 29696 55616
rect 29644 55573 29653 55607
rect 29653 55573 29687 55607
rect 29687 55573 29696 55607
rect 29644 55564 29696 55573
rect 2610 55462 2662 55514
rect 2674 55462 2726 55514
rect 2738 55462 2790 55514
rect 2802 55462 2854 55514
rect 2866 55462 2918 55514
rect 7610 55462 7662 55514
rect 7674 55462 7726 55514
rect 7738 55462 7790 55514
rect 7802 55462 7854 55514
rect 7866 55462 7918 55514
rect 12610 55462 12662 55514
rect 12674 55462 12726 55514
rect 12738 55462 12790 55514
rect 12802 55462 12854 55514
rect 12866 55462 12918 55514
rect 17610 55462 17662 55514
rect 17674 55462 17726 55514
rect 17738 55462 17790 55514
rect 17802 55462 17854 55514
rect 17866 55462 17918 55514
rect 22610 55462 22662 55514
rect 22674 55462 22726 55514
rect 22738 55462 22790 55514
rect 22802 55462 22854 55514
rect 22866 55462 22918 55514
rect 27610 55462 27662 55514
rect 27674 55462 27726 55514
rect 27738 55462 27790 55514
rect 27802 55462 27854 55514
rect 27866 55462 27918 55514
rect 32610 55462 32662 55514
rect 32674 55462 32726 55514
rect 32738 55462 32790 55514
rect 32802 55462 32854 55514
rect 32866 55462 32918 55514
rect 37610 55462 37662 55514
rect 37674 55462 37726 55514
rect 37738 55462 37790 55514
rect 37802 55462 37854 55514
rect 37866 55462 37918 55514
rect 16856 55292 16908 55344
rect 20536 55267 20588 55276
rect 20536 55233 20545 55267
rect 20545 55233 20579 55267
rect 20579 55233 20588 55267
rect 20536 55224 20588 55233
rect 22284 55292 22336 55344
rect 27436 55360 27488 55412
rect 29920 55292 29972 55344
rect 30564 55267 30616 55276
rect 30564 55233 30573 55267
rect 30573 55233 30607 55267
rect 30607 55233 30616 55267
rect 30564 55224 30616 55233
rect 39856 55267 39908 55276
rect 39856 55233 39865 55267
rect 39865 55233 39899 55267
rect 39899 55233 39908 55267
rect 39856 55224 39908 55233
rect 39948 55267 40000 55276
rect 39948 55233 39957 55267
rect 39957 55233 39991 55267
rect 39991 55233 40000 55267
rect 39948 55224 40000 55233
rect 23020 55020 23072 55072
rect 1950 54918 2002 54970
rect 2014 54918 2066 54970
rect 2078 54918 2130 54970
rect 2142 54918 2194 54970
rect 2206 54918 2258 54970
rect 6950 54918 7002 54970
rect 7014 54918 7066 54970
rect 7078 54918 7130 54970
rect 7142 54918 7194 54970
rect 7206 54918 7258 54970
rect 11950 54918 12002 54970
rect 12014 54918 12066 54970
rect 12078 54918 12130 54970
rect 12142 54918 12194 54970
rect 12206 54918 12258 54970
rect 16950 54918 17002 54970
rect 17014 54918 17066 54970
rect 17078 54918 17130 54970
rect 17142 54918 17194 54970
rect 17206 54918 17258 54970
rect 21950 54918 22002 54970
rect 22014 54918 22066 54970
rect 22078 54918 22130 54970
rect 22142 54918 22194 54970
rect 22206 54918 22258 54970
rect 26950 54918 27002 54970
rect 27014 54918 27066 54970
rect 27078 54918 27130 54970
rect 27142 54918 27194 54970
rect 27206 54918 27258 54970
rect 31950 54918 32002 54970
rect 32014 54918 32066 54970
rect 32078 54918 32130 54970
rect 32142 54918 32194 54970
rect 32206 54918 32258 54970
rect 36950 54918 37002 54970
rect 37014 54918 37066 54970
rect 37078 54918 37130 54970
rect 37142 54918 37194 54970
rect 37206 54918 37258 54970
rect 23388 54680 23440 54732
rect 39028 54680 39080 54732
rect 22376 54476 22428 54528
rect 34980 54476 35032 54528
rect 39212 54612 39264 54664
rect 39672 54655 39724 54664
rect 39672 54621 39681 54655
rect 39681 54621 39715 54655
rect 39715 54621 39724 54655
rect 39672 54612 39724 54621
rect 39580 54519 39632 54528
rect 39580 54485 39589 54519
rect 39589 54485 39623 54519
rect 39623 54485 39632 54519
rect 39580 54476 39632 54485
rect 2610 54374 2662 54426
rect 2674 54374 2726 54426
rect 2738 54374 2790 54426
rect 2802 54374 2854 54426
rect 2866 54374 2918 54426
rect 7610 54374 7662 54426
rect 7674 54374 7726 54426
rect 7738 54374 7790 54426
rect 7802 54374 7854 54426
rect 7866 54374 7918 54426
rect 12610 54374 12662 54426
rect 12674 54374 12726 54426
rect 12738 54374 12790 54426
rect 12802 54374 12854 54426
rect 12866 54374 12918 54426
rect 17610 54374 17662 54426
rect 17674 54374 17726 54426
rect 17738 54374 17790 54426
rect 17802 54374 17854 54426
rect 17866 54374 17918 54426
rect 22610 54374 22662 54426
rect 22674 54374 22726 54426
rect 22738 54374 22790 54426
rect 22802 54374 22854 54426
rect 22866 54374 22918 54426
rect 27610 54374 27662 54426
rect 27674 54374 27726 54426
rect 27738 54374 27790 54426
rect 27802 54374 27854 54426
rect 27866 54374 27918 54426
rect 32610 54374 32662 54426
rect 32674 54374 32726 54426
rect 32738 54374 32790 54426
rect 32802 54374 32854 54426
rect 32866 54374 32918 54426
rect 37610 54374 37662 54426
rect 37674 54374 37726 54426
rect 37738 54374 37790 54426
rect 37802 54374 37854 54426
rect 37866 54374 37918 54426
rect 8392 54179 8444 54188
rect 8392 54145 8401 54179
rect 8401 54145 8435 54179
rect 8435 54145 8444 54179
rect 8392 54136 8444 54145
rect 9772 54136 9824 54188
rect 14740 54136 14792 54188
rect 23112 54204 23164 54256
rect 22376 54136 22428 54188
rect 8668 54111 8720 54120
rect 8668 54077 8677 54111
rect 8677 54077 8711 54111
rect 8711 54077 8720 54111
rect 8668 54068 8720 54077
rect 17408 54043 17460 54052
rect 17408 54009 17417 54043
rect 17417 54009 17451 54043
rect 17451 54009 17460 54043
rect 17408 54000 17460 54009
rect 13820 53932 13872 53984
rect 23388 54068 23440 54120
rect 1950 53830 2002 53882
rect 2014 53830 2066 53882
rect 2078 53830 2130 53882
rect 2142 53830 2194 53882
rect 2206 53830 2258 53882
rect 6950 53830 7002 53882
rect 7014 53830 7066 53882
rect 7078 53830 7130 53882
rect 7142 53830 7194 53882
rect 7206 53830 7258 53882
rect 11950 53830 12002 53882
rect 12014 53830 12066 53882
rect 12078 53830 12130 53882
rect 12142 53830 12194 53882
rect 12206 53830 12258 53882
rect 16950 53830 17002 53882
rect 17014 53830 17066 53882
rect 17078 53830 17130 53882
rect 17142 53830 17194 53882
rect 17206 53830 17258 53882
rect 21950 53830 22002 53882
rect 22014 53830 22066 53882
rect 22078 53830 22130 53882
rect 22142 53830 22194 53882
rect 22206 53830 22258 53882
rect 26950 53830 27002 53882
rect 27014 53830 27066 53882
rect 27078 53830 27130 53882
rect 27142 53830 27194 53882
rect 27206 53830 27258 53882
rect 31950 53830 32002 53882
rect 32014 53830 32066 53882
rect 32078 53830 32130 53882
rect 32142 53830 32194 53882
rect 32206 53830 32258 53882
rect 36950 53830 37002 53882
rect 37014 53830 37066 53882
rect 37078 53830 37130 53882
rect 37142 53830 37194 53882
rect 37206 53830 37258 53882
rect 38292 53728 38344 53780
rect 28908 53592 28960 53644
rect 13544 53567 13596 53576
rect 13544 53533 13553 53567
rect 13553 53533 13587 53567
rect 13587 53533 13596 53567
rect 13544 53524 13596 53533
rect 27436 53524 27488 53576
rect 36084 53524 36136 53576
rect 25320 53456 25372 53508
rect 31576 53456 31628 53508
rect 34520 53456 34572 53508
rect 17316 53388 17368 53440
rect 37464 53456 37516 53508
rect 2610 53286 2662 53338
rect 2674 53286 2726 53338
rect 2738 53286 2790 53338
rect 2802 53286 2854 53338
rect 2866 53286 2918 53338
rect 7610 53286 7662 53338
rect 7674 53286 7726 53338
rect 7738 53286 7790 53338
rect 7802 53286 7854 53338
rect 7866 53286 7918 53338
rect 12610 53286 12662 53338
rect 12674 53286 12726 53338
rect 12738 53286 12790 53338
rect 12802 53286 12854 53338
rect 12866 53286 12918 53338
rect 17610 53286 17662 53338
rect 17674 53286 17726 53338
rect 17738 53286 17790 53338
rect 17802 53286 17854 53338
rect 17866 53286 17918 53338
rect 22610 53286 22662 53338
rect 22674 53286 22726 53338
rect 22738 53286 22790 53338
rect 22802 53286 22854 53338
rect 22866 53286 22918 53338
rect 27610 53286 27662 53338
rect 27674 53286 27726 53338
rect 27738 53286 27790 53338
rect 27802 53286 27854 53338
rect 27866 53286 27918 53338
rect 32610 53286 32662 53338
rect 32674 53286 32726 53338
rect 32738 53286 32790 53338
rect 32802 53286 32854 53338
rect 32866 53286 32918 53338
rect 37610 53286 37662 53338
rect 37674 53286 37726 53338
rect 37738 53286 37790 53338
rect 37802 53286 37854 53338
rect 37866 53286 37918 53338
rect 22376 53184 22428 53236
rect 31576 53184 31628 53236
rect 6368 53116 6420 53168
rect 23296 52980 23348 53032
rect 24676 53023 24728 53032
rect 24676 52989 24685 53023
rect 24685 52989 24719 53023
rect 24719 52989 24728 53023
rect 24676 52980 24728 52989
rect 28908 52980 28960 53032
rect 5264 52844 5316 52896
rect 25044 52844 25096 52896
rect 1950 52742 2002 52794
rect 2014 52742 2066 52794
rect 2078 52742 2130 52794
rect 2142 52742 2194 52794
rect 2206 52742 2258 52794
rect 6950 52742 7002 52794
rect 7014 52742 7066 52794
rect 7078 52742 7130 52794
rect 7142 52742 7194 52794
rect 7206 52742 7258 52794
rect 11950 52742 12002 52794
rect 12014 52742 12066 52794
rect 12078 52742 12130 52794
rect 12142 52742 12194 52794
rect 12206 52742 12258 52794
rect 16950 52742 17002 52794
rect 17014 52742 17066 52794
rect 17078 52742 17130 52794
rect 17142 52742 17194 52794
rect 17206 52742 17258 52794
rect 21950 52742 22002 52794
rect 22014 52742 22066 52794
rect 22078 52742 22130 52794
rect 22142 52742 22194 52794
rect 22206 52742 22258 52794
rect 26950 52742 27002 52794
rect 27014 52742 27066 52794
rect 27078 52742 27130 52794
rect 27142 52742 27194 52794
rect 27206 52742 27258 52794
rect 31950 52742 32002 52794
rect 32014 52742 32066 52794
rect 32078 52742 32130 52794
rect 32142 52742 32194 52794
rect 32206 52742 32258 52794
rect 36950 52742 37002 52794
rect 37014 52742 37066 52794
rect 37078 52742 37130 52794
rect 37142 52742 37194 52794
rect 37206 52742 37258 52794
rect 4068 52640 4120 52692
rect 33140 52572 33192 52624
rect 5080 52479 5132 52488
rect 5080 52445 5089 52479
rect 5089 52445 5123 52479
rect 5123 52445 5132 52479
rect 5080 52436 5132 52445
rect 5264 52479 5316 52488
rect 5264 52445 5273 52479
rect 5273 52445 5307 52479
rect 5307 52445 5316 52479
rect 5264 52436 5316 52445
rect 25320 52504 25372 52556
rect 5632 52479 5684 52488
rect 5632 52445 5641 52479
rect 5641 52445 5675 52479
rect 5675 52445 5684 52479
rect 5632 52436 5684 52445
rect 15936 52436 15988 52488
rect 24124 52479 24176 52488
rect 24124 52445 24133 52479
rect 24133 52445 24167 52479
rect 24167 52445 24176 52479
rect 24124 52436 24176 52445
rect 25044 52436 25096 52488
rect 26056 52436 26108 52488
rect 4344 52411 4396 52420
rect 4344 52377 4353 52411
rect 4353 52377 4387 52411
rect 4387 52377 4396 52411
rect 4344 52368 4396 52377
rect 18696 52368 18748 52420
rect 28540 52368 28592 52420
rect 28816 52368 28868 52420
rect 6184 52300 6236 52352
rect 25504 52300 25556 52352
rect 36360 52436 36412 52488
rect 34152 52300 34204 52352
rect 38200 52368 38252 52420
rect 2610 52198 2662 52250
rect 2674 52198 2726 52250
rect 2738 52198 2790 52250
rect 2802 52198 2854 52250
rect 2866 52198 2918 52250
rect 7610 52198 7662 52250
rect 7674 52198 7726 52250
rect 7738 52198 7790 52250
rect 7802 52198 7854 52250
rect 7866 52198 7918 52250
rect 12610 52198 12662 52250
rect 12674 52198 12726 52250
rect 12738 52198 12790 52250
rect 12802 52198 12854 52250
rect 12866 52198 12918 52250
rect 17610 52198 17662 52250
rect 17674 52198 17726 52250
rect 17738 52198 17790 52250
rect 17802 52198 17854 52250
rect 17866 52198 17918 52250
rect 22610 52198 22662 52250
rect 22674 52198 22726 52250
rect 22738 52198 22790 52250
rect 22802 52198 22854 52250
rect 22866 52198 22918 52250
rect 27610 52198 27662 52250
rect 27674 52198 27726 52250
rect 27738 52198 27790 52250
rect 27802 52198 27854 52250
rect 27866 52198 27918 52250
rect 32610 52198 32662 52250
rect 32674 52198 32726 52250
rect 32738 52198 32790 52250
rect 32802 52198 32854 52250
rect 32866 52198 32918 52250
rect 37610 52198 37662 52250
rect 37674 52198 37726 52250
rect 37738 52198 37790 52250
rect 37802 52198 37854 52250
rect 37866 52198 37918 52250
rect 4344 52139 4396 52148
rect 4344 52105 4353 52139
rect 4353 52105 4387 52139
rect 4387 52105 4396 52139
rect 4344 52096 4396 52105
rect 11060 52096 11112 52148
rect 12348 52096 12400 52148
rect 4068 51960 4120 52012
rect 10416 52003 10468 52012
rect 10416 51969 10425 52003
rect 10425 51969 10459 52003
rect 10459 51969 10468 52003
rect 10416 51960 10468 51969
rect 13820 51960 13872 52012
rect 10232 51935 10284 51944
rect 10232 51901 10241 51935
rect 10241 51901 10275 51935
rect 10275 51901 10284 51935
rect 10232 51892 10284 51901
rect 17500 51892 17552 51944
rect 32312 51960 32364 52012
rect 27528 51892 27580 51944
rect 21364 51824 21416 51876
rect 33048 51824 33100 51876
rect 31300 51799 31352 51808
rect 31300 51765 31309 51799
rect 31309 51765 31343 51799
rect 31343 51765 31352 51799
rect 31300 51756 31352 51765
rect 33140 51756 33192 51808
rect 1950 51654 2002 51706
rect 2014 51654 2066 51706
rect 2078 51654 2130 51706
rect 2142 51654 2194 51706
rect 2206 51654 2258 51706
rect 6950 51654 7002 51706
rect 7014 51654 7066 51706
rect 7078 51654 7130 51706
rect 7142 51654 7194 51706
rect 7206 51654 7258 51706
rect 11950 51654 12002 51706
rect 12014 51654 12066 51706
rect 12078 51654 12130 51706
rect 12142 51654 12194 51706
rect 12206 51654 12258 51706
rect 16950 51654 17002 51706
rect 17014 51654 17066 51706
rect 17078 51654 17130 51706
rect 17142 51654 17194 51706
rect 17206 51654 17258 51706
rect 21950 51654 22002 51706
rect 22014 51654 22066 51706
rect 22078 51654 22130 51706
rect 22142 51654 22194 51706
rect 22206 51654 22258 51706
rect 26950 51654 27002 51706
rect 27014 51654 27066 51706
rect 27078 51654 27130 51706
rect 27142 51654 27194 51706
rect 27206 51654 27258 51706
rect 31950 51654 32002 51706
rect 32014 51654 32066 51706
rect 32078 51654 32130 51706
rect 32142 51654 32194 51706
rect 32206 51654 32258 51706
rect 36950 51654 37002 51706
rect 37014 51654 37066 51706
rect 37078 51654 37130 51706
rect 37142 51654 37194 51706
rect 37206 51654 37258 51706
rect 28816 51552 28868 51604
rect 34152 51552 34204 51604
rect 11244 51391 11296 51400
rect 11244 51357 11253 51391
rect 11253 51357 11287 51391
rect 11287 51357 11296 51391
rect 11704 51416 11756 51468
rect 11244 51348 11296 51357
rect 10784 51323 10836 51332
rect 10784 51289 10793 51323
rect 10793 51289 10827 51323
rect 10827 51289 10836 51323
rect 10784 51280 10836 51289
rect 11336 51323 11388 51332
rect 11336 51289 11345 51323
rect 11345 51289 11379 51323
rect 11379 51289 11388 51323
rect 11336 51280 11388 51289
rect 16580 51391 16632 51400
rect 16580 51357 16589 51391
rect 16589 51357 16623 51391
rect 16623 51357 16632 51391
rect 16580 51348 16632 51357
rect 18696 51416 18748 51468
rect 16856 51391 16908 51400
rect 16856 51357 16865 51391
rect 16865 51357 16899 51391
rect 16899 51357 16908 51391
rect 16856 51348 16908 51357
rect 17316 51348 17368 51400
rect 17500 51348 17552 51400
rect 17960 51348 18012 51400
rect 19616 51280 19668 51332
rect 19984 51280 20036 51332
rect 11612 51212 11664 51264
rect 34520 51280 34572 51332
rect 33140 51255 33192 51264
rect 33140 51221 33149 51255
rect 33149 51221 33183 51255
rect 33183 51221 33192 51255
rect 33140 51212 33192 51221
rect 2610 51110 2662 51162
rect 2674 51110 2726 51162
rect 2738 51110 2790 51162
rect 2802 51110 2854 51162
rect 2866 51110 2918 51162
rect 7610 51110 7662 51162
rect 7674 51110 7726 51162
rect 7738 51110 7790 51162
rect 7802 51110 7854 51162
rect 7866 51110 7918 51162
rect 12610 51110 12662 51162
rect 12674 51110 12726 51162
rect 12738 51110 12790 51162
rect 12802 51110 12854 51162
rect 12866 51110 12918 51162
rect 17610 51110 17662 51162
rect 17674 51110 17726 51162
rect 17738 51110 17790 51162
rect 17802 51110 17854 51162
rect 17866 51110 17918 51162
rect 22610 51110 22662 51162
rect 22674 51110 22726 51162
rect 22738 51110 22790 51162
rect 22802 51110 22854 51162
rect 22866 51110 22918 51162
rect 27610 51110 27662 51162
rect 27674 51110 27726 51162
rect 27738 51110 27790 51162
rect 27802 51110 27854 51162
rect 27866 51110 27918 51162
rect 32610 51110 32662 51162
rect 32674 51110 32726 51162
rect 32738 51110 32790 51162
rect 32802 51110 32854 51162
rect 32866 51110 32918 51162
rect 37610 51110 37662 51162
rect 37674 51110 37726 51162
rect 37738 51110 37790 51162
rect 37802 51110 37854 51162
rect 37866 51110 37918 51162
rect 13084 50915 13136 50924
rect 13084 50881 13093 50915
rect 13093 50881 13127 50915
rect 13127 50881 13136 50915
rect 13084 50872 13136 50881
rect 12440 50804 12492 50856
rect 29092 50804 29144 50856
rect 8300 50736 8352 50788
rect 8484 50736 8536 50788
rect 12992 50779 13044 50788
rect 12992 50745 13001 50779
rect 13001 50745 13035 50779
rect 13035 50745 13044 50779
rect 12992 50736 13044 50745
rect 22376 50668 22428 50720
rect 1950 50566 2002 50618
rect 2014 50566 2066 50618
rect 2078 50566 2130 50618
rect 2142 50566 2194 50618
rect 2206 50566 2258 50618
rect 6950 50566 7002 50618
rect 7014 50566 7066 50618
rect 7078 50566 7130 50618
rect 7142 50566 7194 50618
rect 7206 50566 7258 50618
rect 11950 50566 12002 50618
rect 12014 50566 12066 50618
rect 12078 50566 12130 50618
rect 12142 50566 12194 50618
rect 12206 50566 12258 50618
rect 16950 50566 17002 50618
rect 17014 50566 17066 50618
rect 17078 50566 17130 50618
rect 17142 50566 17194 50618
rect 17206 50566 17258 50618
rect 21950 50566 22002 50618
rect 22014 50566 22066 50618
rect 22078 50566 22130 50618
rect 22142 50566 22194 50618
rect 22206 50566 22258 50618
rect 26950 50566 27002 50618
rect 27014 50566 27066 50618
rect 27078 50566 27130 50618
rect 27142 50566 27194 50618
rect 27206 50566 27258 50618
rect 31950 50566 32002 50618
rect 32014 50566 32066 50618
rect 32078 50566 32130 50618
rect 32142 50566 32194 50618
rect 32206 50566 32258 50618
rect 36950 50566 37002 50618
rect 37014 50566 37066 50618
rect 37078 50566 37130 50618
rect 37142 50566 37194 50618
rect 37206 50566 37258 50618
rect 29552 50464 29604 50516
rect 24952 50303 25004 50312
rect 24952 50269 24961 50303
rect 24961 50269 24995 50303
rect 24995 50269 25004 50303
rect 24952 50260 25004 50269
rect 14372 50192 14424 50244
rect 14832 50192 14884 50244
rect 24860 50192 24912 50244
rect 37464 50328 37516 50380
rect 38384 50328 38436 50380
rect 34152 50235 34204 50244
rect 34152 50201 34161 50235
rect 34161 50201 34195 50235
rect 34195 50201 34204 50235
rect 34152 50192 34204 50201
rect 38660 50192 38712 50244
rect 33784 50167 33836 50176
rect 33784 50133 33793 50167
rect 33793 50133 33827 50167
rect 33827 50133 33836 50167
rect 33784 50124 33836 50133
rect 33968 50167 34020 50176
rect 33968 50133 33977 50167
rect 33977 50133 34011 50167
rect 34011 50133 34020 50167
rect 33968 50124 34020 50133
rect 36544 50124 36596 50176
rect 2610 50022 2662 50074
rect 2674 50022 2726 50074
rect 2738 50022 2790 50074
rect 2802 50022 2854 50074
rect 2866 50022 2918 50074
rect 7610 50022 7662 50074
rect 7674 50022 7726 50074
rect 7738 50022 7790 50074
rect 7802 50022 7854 50074
rect 7866 50022 7918 50074
rect 12610 50022 12662 50074
rect 12674 50022 12726 50074
rect 12738 50022 12790 50074
rect 12802 50022 12854 50074
rect 12866 50022 12918 50074
rect 17610 50022 17662 50074
rect 17674 50022 17726 50074
rect 17738 50022 17790 50074
rect 17802 50022 17854 50074
rect 17866 50022 17918 50074
rect 22610 50022 22662 50074
rect 22674 50022 22726 50074
rect 22738 50022 22790 50074
rect 22802 50022 22854 50074
rect 22866 50022 22918 50074
rect 27610 50022 27662 50074
rect 27674 50022 27726 50074
rect 27738 50022 27790 50074
rect 27802 50022 27854 50074
rect 27866 50022 27918 50074
rect 32610 50022 32662 50074
rect 32674 50022 32726 50074
rect 32738 50022 32790 50074
rect 32802 50022 32854 50074
rect 32866 50022 32918 50074
rect 37610 50022 37662 50074
rect 37674 50022 37726 50074
rect 37738 50022 37790 50074
rect 37802 50022 37854 50074
rect 37866 50022 37918 50074
rect 29368 49920 29420 49972
rect 10968 49784 11020 49836
rect 15108 49784 15160 49836
rect 29092 49827 29144 49836
rect 29092 49793 29101 49827
rect 29101 49793 29135 49827
rect 29135 49793 29144 49827
rect 29092 49784 29144 49793
rect 36544 49716 36596 49768
rect 36728 49716 36780 49768
rect 1950 49478 2002 49530
rect 2014 49478 2066 49530
rect 2078 49478 2130 49530
rect 2142 49478 2194 49530
rect 2206 49478 2258 49530
rect 6950 49478 7002 49530
rect 7014 49478 7066 49530
rect 7078 49478 7130 49530
rect 7142 49478 7194 49530
rect 7206 49478 7258 49530
rect 11950 49478 12002 49530
rect 12014 49478 12066 49530
rect 12078 49478 12130 49530
rect 12142 49478 12194 49530
rect 12206 49478 12258 49530
rect 16950 49478 17002 49530
rect 17014 49478 17066 49530
rect 17078 49478 17130 49530
rect 17142 49478 17194 49530
rect 17206 49478 17258 49530
rect 21950 49478 22002 49530
rect 22014 49478 22066 49530
rect 22078 49478 22130 49530
rect 22142 49478 22194 49530
rect 22206 49478 22258 49530
rect 26950 49478 27002 49530
rect 27014 49478 27066 49530
rect 27078 49478 27130 49530
rect 27142 49478 27194 49530
rect 27206 49478 27258 49530
rect 31950 49478 32002 49530
rect 32014 49478 32066 49530
rect 32078 49478 32130 49530
rect 32142 49478 32194 49530
rect 32206 49478 32258 49530
rect 36950 49478 37002 49530
rect 37014 49478 37066 49530
rect 37078 49478 37130 49530
rect 37142 49478 37194 49530
rect 37206 49478 37258 49530
rect 24768 49376 24820 49428
rect 33416 49376 33468 49428
rect 33600 49376 33652 49428
rect 14464 49104 14516 49156
rect 15016 49104 15068 49156
rect 9036 49036 9088 49088
rect 24400 49079 24452 49088
rect 24400 49045 24409 49079
rect 24409 49045 24443 49079
rect 24443 49045 24452 49079
rect 24400 49036 24452 49045
rect 26516 49104 26568 49156
rect 33324 49147 33376 49156
rect 33324 49113 33333 49147
rect 33333 49113 33367 49147
rect 33367 49113 33376 49147
rect 33324 49104 33376 49113
rect 31760 49036 31812 49088
rect 33140 49079 33192 49088
rect 33140 49045 33167 49079
rect 33167 49045 33192 49079
rect 33140 49036 33192 49045
rect 2610 48934 2662 48986
rect 2674 48934 2726 48986
rect 2738 48934 2790 48986
rect 2802 48934 2854 48986
rect 2866 48934 2918 48986
rect 7610 48934 7662 48986
rect 7674 48934 7726 48986
rect 7738 48934 7790 48986
rect 7802 48934 7854 48986
rect 7866 48934 7918 48986
rect 12610 48934 12662 48986
rect 12674 48934 12726 48986
rect 12738 48934 12790 48986
rect 12802 48934 12854 48986
rect 12866 48934 12918 48986
rect 17610 48934 17662 48986
rect 17674 48934 17726 48986
rect 17738 48934 17790 48986
rect 17802 48934 17854 48986
rect 17866 48934 17918 48986
rect 22610 48934 22662 48986
rect 22674 48934 22726 48986
rect 22738 48934 22790 48986
rect 22802 48934 22854 48986
rect 22866 48934 22918 48986
rect 27610 48934 27662 48986
rect 27674 48934 27726 48986
rect 27738 48934 27790 48986
rect 27802 48934 27854 48986
rect 27866 48934 27918 48986
rect 32610 48934 32662 48986
rect 32674 48934 32726 48986
rect 32738 48934 32790 48986
rect 32802 48934 32854 48986
rect 32866 48934 32918 48986
rect 37610 48934 37662 48986
rect 37674 48934 37726 48986
rect 37738 48934 37790 48986
rect 37802 48934 37854 48986
rect 37866 48934 37918 48986
rect 9404 48696 9456 48748
rect 12440 48696 12492 48748
rect 21640 48739 21692 48748
rect 21640 48705 21649 48739
rect 21649 48705 21683 48739
rect 21683 48705 21692 48739
rect 21640 48696 21692 48705
rect 4988 48492 5040 48544
rect 20996 48492 21048 48544
rect 1950 48390 2002 48442
rect 2014 48390 2066 48442
rect 2078 48390 2130 48442
rect 2142 48390 2194 48442
rect 2206 48390 2258 48442
rect 6950 48390 7002 48442
rect 7014 48390 7066 48442
rect 7078 48390 7130 48442
rect 7142 48390 7194 48442
rect 7206 48390 7258 48442
rect 11950 48390 12002 48442
rect 12014 48390 12066 48442
rect 12078 48390 12130 48442
rect 12142 48390 12194 48442
rect 12206 48390 12258 48442
rect 16950 48390 17002 48442
rect 17014 48390 17066 48442
rect 17078 48390 17130 48442
rect 17142 48390 17194 48442
rect 17206 48390 17258 48442
rect 21950 48390 22002 48442
rect 22014 48390 22066 48442
rect 22078 48390 22130 48442
rect 22142 48390 22194 48442
rect 22206 48390 22258 48442
rect 26950 48390 27002 48442
rect 27014 48390 27066 48442
rect 27078 48390 27130 48442
rect 27142 48390 27194 48442
rect 27206 48390 27258 48442
rect 31950 48390 32002 48442
rect 32014 48390 32066 48442
rect 32078 48390 32130 48442
rect 32142 48390 32194 48442
rect 32206 48390 32258 48442
rect 36950 48390 37002 48442
rect 37014 48390 37066 48442
rect 37078 48390 37130 48442
rect 37142 48390 37194 48442
rect 37206 48390 37258 48442
rect 26516 48288 26568 48340
rect 33416 48288 33468 48340
rect 3424 48152 3476 48204
rect 4068 48152 4120 48204
rect 25780 48220 25832 48272
rect 33600 48152 33652 48204
rect 30380 48127 30432 48136
rect 30380 48093 30389 48127
rect 30389 48093 30423 48127
rect 30423 48093 30432 48127
rect 30380 48084 30432 48093
rect 33876 48127 33928 48136
rect 33876 48093 33885 48127
rect 33885 48093 33919 48127
rect 33919 48093 33928 48127
rect 33876 48084 33928 48093
rect 15936 48016 15988 48068
rect 29736 48059 29788 48068
rect 29736 48025 29745 48059
rect 29745 48025 29779 48059
rect 29779 48025 29788 48059
rect 29736 48016 29788 48025
rect 6092 47948 6144 48000
rect 6828 47948 6880 48000
rect 2610 47846 2662 47898
rect 2674 47846 2726 47898
rect 2738 47846 2790 47898
rect 2802 47846 2854 47898
rect 2866 47846 2918 47898
rect 7610 47846 7662 47898
rect 7674 47846 7726 47898
rect 7738 47846 7790 47898
rect 7802 47846 7854 47898
rect 7866 47846 7918 47898
rect 12610 47846 12662 47898
rect 12674 47846 12726 47898
rect 12738 47846 12790 47898
rect 12802 47846 12854 47898
rect 12866 47846 12918 47898
rect 17610 47846 17662 47898
rect 17674 47846 17726 47898
rect 17738 47846 17790 47898
rect 17802 47846 17854 47898
rect 17866 47846 17918 47898
rect 22610 47846 22662 47898
rect 22674 47846 22726 47898
rect 22738 47846 22790 47898
rect 22802 47846 22854 47898
rect 22866 47846 22918 47898
rect 27610 47846 27662 47898
rect 27674 47846 27726 47898
rect 27738 47846 27790 47898
rect 27802 47846 27854 47898
rect 27866 47846 27918 47898
rect 32610 47846 32662 47898
rect 32674 47846 32726 47898
rect 32738 47846 32790 47898
rect 32802 47846 32854 47898
rect 32866 47846 32918 47898
rect 37610 47846 37662 47898
rect 37674 47846 37726 47898
rect 37738 47846 37790 47898
rect 37802 47846 37854 47898
rect 37866 47846 37918 47898
rect 30380 47608 30432 47660
rect 40224 47608 40276 47660
rect 13820 47540 13872 47592
rect 21456 47540 21508 47592
rect 35164 47447 35216 47456
rect 35164 47413 35173 47447
rect 35173 47413 35207 47447
rect 35207 47413 35216 47447
rect 35164 47404 35216 47413
rect 1950 47302 2002 47354
rect 2014 47302 2066 47354
rect 2078 47302 2130 47354
rect 2142 47302 2194 47354
rect 2206 47302 2258 47354
rect 6950 47302 7002 47354
rect 7014 47302 7066 47354
rect 7078 47302 7130 47354
rect 7142 47302 7194 47354
rect 7206 47302 7258 47354
rect 11950 47302 12002 47354
rect 12014 47302 12066 47354
rect 12078 47302 12130 47354
rect 12142 47302 12194 47354
rect 12206 47302 12258 47354
rect 16950 47302 17002 47354
rect 17014 47302 17066 47354
rect 17078 47302 17130 47354
rect 17142 47302 17194 47354
rect 17206 47302 17258 47354
rect 21950 47302 22002 47354
rect 22014 47302 22066 47354
rect 22078 47302 22130 47354
rect 22142 47302 22194 47354
rect 22206 47302 22258 47354
rect 26950 47302 27002 47354
rect 27014 47302 27066 47354
rect 27078 47302 27130 47354
rect 27142 47302 27194 47354
rect 27206 47302 27258 47354
rect 31950 47302 32002 47354
rect 32014 47302 32066 47354
rect 32078 47302 32130 47354
rect 32142 47302 32194 47354
rect 32206 47302 32258 47354
rect 36950 47302 37002 47354
rect 37014 47302 37066 47354
rect 37078 47302 37130 47354
rect 37142 47302 37194 47354
rect 37206 47302 37258 47354
rect 38108 47200 38160 47252
rect 33048 47132 33100 47184
rect 13820 47064 13872 47116
rect 25412 47064 25464 47116
rect 25780 47064 25832 47116
rect 1676 47039 1728 47048
rect 1676 47005 1685 47039
rect 1685 47005 1719 47039
rect 1719 47005 1728 47039
rect 1676 46996 1728 47005
rect 10324 46996 10376 47048
rect 30380 46996 30432 47048
rect 30472 46996 30524 47048
rect 38200 46996 38252 47048
rect 19892 46928 19944 46980
rect 1860 46903 1912 46912
rect 1860 46869 1869 46903
rect 1869 46869 1903 46903
rect 1903 46869 1912 46903
rect 1860 46860 1912 46869
rect 2610 46758 2662 46810
rect 2674 46758 2726 46810
rect 2738 46758 2790 46810
rect 2802 46758 2854 46810
rect 2866 46758 2918 46810
rect 7610 46758 7662 46810
rect 7674 46758 7726 46810
rect 7738 46758 7790 46810
rect 7802 46758 7854 46810
rect 7866 46758 7918 46810
rect 12610 46758 12662 46810
rect 12674 46758 12726 46810
rect 12738 46758 12790 46810
rect 12802 46758 12854 46810
rect 12866 46758 12918 46810
rect 17610 46758 17662 46810
rect 17674 46758 17726 46810
rect 17738 46758 17790 46810
rect 17802 46758 17854 46810
rect 17866 46758 17918 46810
rect 22610 46758 22662 46810
rect 22674 46758 22726 46810
rect 22738 46758 22790 46810
rect 22802 46758 22854 46810
rect 22866 46758 22918 46810
rect 27610 46758 27662 46810
rect 27674 46758 27726 46810
rect 27738 46758 27790 46810
rect 27802 46758 27854 46810
rect 27866 46758 27918 46810
rect 32610 46758 32662 46810
rect 32674 46758 32726 46810
rect 32738 46758 32790 46810
rect 32802 46758 32854 46810
rect 32866 46758 32918 46810
rect 37610 46758 37662 46810
rect 37674 46758 37726 46810
rect 37738 46758 37790 46810
rect 37802 46758 37854 46810
rect 37866 46758 37918 46810
rect 28816 46563 28868 46572
rect 28816 46529 28825 46563
rect 28825 46529 28859 46563
rect 28859 46529 28868 46563
rect 28816 46520 28868 46529
rect 28908 46316 28960 46368
rect 1950 46214 2002 46266
rect 2014 46214 2066 46266
rect 2078 46214 2130 46266
rect 2142 46214 2194 46266
rect 2206 46214 2258 46266
rect 6950 46214 7002 46266
rect 7014 46214 7066 46266
rect 7078 46214 7130 46266
rect 7142 46214 7194 46266
rect 7206 46214 7258 46266
rect 11950 46214 12002 46266
rect 12014 46214 12066 46266
rect 12078 46214 12130 46266
rect 12142 46214 12194 46266
rect 12206 46214 12258 46266
rect 16950 46214 17002 46266
rect 17014 46214 17066 46266
rect 17078 46214 17130 46266
rect 17142 46214 17194 46266
rect 17206 46214 17258 46266
rect 21950 46214 22002 46266
rect 22014 46214 22066 46266
rect 22078 46214 22130 46266
rect 22142 46214 22194 46266
rect 22206 46214 22258 46266
rect 26950 46214 27002 46266
rect 27014 46214 27066 46266
rect 27078 46214 27130 46266
rect 27142 46214 27194 46266
rect 27206 46214 27258 46266
rect 31950 46214 32002 46266
rect 32014 46214 32066 46266
rect 32078 46214 32130 46266
rect 32142 46214 32194 46266
rect 32206 46214 32258 46266
rect 36950 46214 37002 46266
rect 37014 46214 37066 46266
rect 37078 46214 37130 46266
rect 37142 46214 37194 46266
rect 37206 46214 37258 46266
rect 34612 46112 34664 46164
rect 9588 45908 9640 45960
rect 14556 45883 14608 45892
rect 14556 45849 14565 45883
rect 14565 45849 14599 45883
rect 14599 45849 14608 45883
rect 14556 45840 14608 45849
rect 15384 45840 15436 45892
rect 29736 45908 29788 45960
rect 23020 45840 23072 45892
rect 26516 45883 26568 45892
rect 26516 45849 26525 45883
rect 26525 45849 26559 45883
rect 26559 45849 26568 45883
rect 26516 45840 26568 45849
rect 28908 45883 28960 45892
rect 28908 45849 28917 45883
rect 28917 45849 28951 45883
rect 28951 45849 28960 45883
rect 28908 45840 28960 45849
rect 18696 45815 18748 45824
rect 18696 45781 18705 45815
rect 18705 45781 18739 45815
rect 18739 45781 18748 45815
rect 18696 45772 18748 45781
rect 25964 45772 26016 45824
rect 2610 45670 2662 45722
rect 2674 45670 2726 45722
rect 2738 45670 2790 45722
rect 2802 45670 2854 45722
rect 2866 45670 2918 45722
rect 7610 45670 7662 45722
rect 7674 45670 7726 45722
rect 7738 45670 7790 45722
rect 7802 45670 7854 45722
rect 7866 45670 7918 45722
rect 12610 45670 12662 45722
rect 12674 45670 12726 45722
rect 12738 45670 12790 45722
rect 12802 45670 12854 45722
rect 12866 45670 12918 45722
rect 17610 45670 17662 45722
rect 17674 45670 17726 45722
rect 17738 45670 17790 45722
rect 17802 45670 17854 45722
rect 17866 45670 17918 45722
rect 22610 45670 22662 45722
rect 22674 45670 22726 45722
rect 22738 45670 22790 45722
rect 22802 45670 22854 45722
rect 22866 45670 22918 45722
rect 27610 45670 27662 45722
rect 27674 45670 27726 45722
rect 27738 45670 27790 45722
rect 27802 45670 27854 45722
rect 27866 45670 27918 45722
rect 32610 45670 32662 45722
rect 32674 45670 32726 45722
rect 32738 45670 32790 45722
rect 32802 45670 32854 45722
rect 32866 45670 32918 45722
rect 37610 45670 37662 45722
rect 37674 45670 37726 45722
rect 37738 45670 37790 45722
rect 37802 45670 37854 45722
rect 37866 45670 37918 45722
rect 8300 45568 8352 45620
rect 9588 45568 9640 45620
rect 3056 45500 3108 45552
rect 14832 45500 14884 45552
rect 1400 45407 1452 45416
rect 1400 45373 1409 45407
rect 1409 45373 1443 45407
rect 1443 45373 1452 45407
rect 1400 45364 1452 45373
rect 8300 45432 8352 45484
rect 16856 45432 16908 45484
rect 3148 45407 3200 45416
rect 3148 45373 3157 45407
rect 3157 45373 3191 45407
rect 3191 45373 3200 45407
rect 3148 45364 3200 45373
rect 14280 45364 14332 45416
rect 35164 45296 35216 45348
rect 1950 45126 2002 45178
rect 2014 45126 2066 45178
rect 2078 45126 2130 45178
rect 2142 45126 2194 45178
rect 2206 45126 2258 45178
rect 6950 45126 7002 45178
rect 7014 45126 7066 45178
rect 7078 45126 7130 45178
rect 7142 45126 7194 45178
rect 7206 45126 7258 45178
rect 11950 45126 12002 45178
rect 12014 45126 12066 45178
rect 12078 45126 12130 45178
rect 12142 45126 12194 45178
rect 12206 45126 12258 45178
rect 16950 45126 17002 45178
rect 17014 45126 17066 45178
rect 17078 45126 17130 45178
rect 17142 45126 17194 45178
rect 17206 45126 17258 45178
rect 21950 45126 22002 45178
rect 22014 45126 22066 45178
rect 22078 45126 22130 45178
rect 22142 45126 22194 45178
rect 22206 45126 22258 45178
rect 26950 45126 27002 45178
rect 27014 45126 27066 45178
rect 27078 45126 27130 45178
rect 27142 45126 27194 45178
rect 27206 45126 27258 45178
rect 31950 45126 32002 45178
rect 32014 45126 32066 45178
rect 32078 45126 32130 45178
rect 32142 45126 32194 45178
rect 32206 45126 32258 45178
rect 36950 45126 37002 45178
rect 37014 45126 37066 45178
rect 37078 45126 37130 45178
rect 37142 45126 37194 45178
rect 37206 45126 37258 45178
rect 1400 45024 1452 45076
rect 10416 45024 10468 45076
rect 5356 44956 5408 45008
rect 19432 44956 19484 45008
rect 3056 44888 3108 44940
rect 2504 44752 2556 44804
rect 5540 44888 5592 44940
rect 10416 44888 10468 44940
rect 20904 44888 20956 44940
rect 5264 44820 5316 44872
rect 5724 44820 5776 44872
rect 19432 44820 19484 44872
rect 35992 44888 36044 44940
rect 30564 44820 30616 44872
rect 5448 44752 5500 44804
rect 8484 44752 8536 44804
rect 5540 44684 5592 44736
rect 22284 44752 22336 44804
rect 22468 44752 22520 44804
rect 22376 44727 22428 44736
rect 22376 44693 22385 44727
rect 22385 44693 22419 44727
rect 22419 44693 22428 44727
rect 22376 44684 22428 44693
rect 2610 44582 2662 44634
rect 2674 44582 2726 44634
rect 2738 44582 2790 44634
rect 2802 44582 2854 44634
rect 2866 44582 2918 44634
rect 7610 44582 7662 44634
rect 7674 44582 7726 44634
rect 7738 44582 7790 44634
rect 7802 44582 7854 44634
rect 7866 44582 7918 44634
rect 12610 44582 12662 44634
rect 12674 44582 12726 44634
rect 12738 44582 12790 44634
rect 12802 44582 12854 44634
rect 12866 44582 12918 44634
rect 17610 44582 17662 44634
rect 17674 44582 17726 44634
rect 17738 44582 17790 44634
rect 17802 44582 17854 44634
rect 17866 44582 17918 44634
rect 22610 44582 22662 44634
rect 22674 44582 22726 44634
rect 22738 44582 22790 44634
rect 22802 44582 22854 44634
rect 22866 44582 22918 44634
rect 27610 44582 27662 44634
rect 27674 44582 27726 44634
rect 27738 44582 27790 44634
rect 27802 44582 27854 44634
rect 27866 44582 27918 44634
rect 32610 44582 32662 44634
rect 32674 44582 32726 44634
rect 32738 44582 32790 44634
rect 32802 44582 32854 44634
rect 32866 44582 32918 44634
rect 37610 44582 37662 44634
rect 37674 44582 37726 44634
rect 37738 44582 37790 44634
rect 37802 44582 37854 44634
rect 37866 44582 37918 44634
rect 14280 44140 14332 44192
rect 14648 44140 14700 44192
rect 16856 44140 16908 44192
rect 17316 44140 17368 44192
rect 1950 44038 2002 44090
rect 2014 44038 2066 44090
rect 2078 44038 2130 44090
rect 2142 44038 2194 44090
rect 2206 44038 2258 44090
rect 6950 44038 7002 44090
rect 7014 44038 7066 44090
rect 7078 44038 7130 44090
rect 7142 44038 7194 44090
rect 7206 44038 7258 44090
rect 11950 44038 12002 44090
rect 12014 44038 12066 44090
rect 12078 44038 12130 44090
rect 12142 44038 12194 44090
rect 12206 44038 12258 44090
rect 16950 44038 17002 44090
rect 17014 44038 17066 44090
rect 17078 44038 17130 44090
rect 17142 44038 17194 44090
rect 17206 44038 17258 44090
rect 21950 44038 22002 44090
rect 22014 44038 22066 44090
rect 22078 44038 22130 44090
rect 22142 44038 22194 44090
rect 22206 44038 22258 44090
rect 26950 44038 27002 44090
rect 27014 44038 27066 44090
rect 27078 44038 27130 44090
rect 27142 44038 27194 44090
rect 27206 44038 27258 44090
rect 31950 44038 32002 44090
rect 32014 44038 32066 44090
rect 32078 44038 32130 44090
rect 32142 44038 32194 44090
rect 32206 44038 32258 44090
rect 36950 44038 37002 44090
rect 37014 44038 37066 44090
rect 37078 44038 37130 44090
rect 37142 44038 37194 44090
rect 37206 44038 37258 44090
rect 24860 43843 24912 43852
rect 24860 43809 24869 43843
rect 24869 43809 24903 43843
rect 24903 43809 24912 43843
rect 24860 43800 24912 43809
rect 25504 43843 25556 43852
rect 25504 43809 25513 43843
rect 25513 43809 25547 43843
rect 25547 43809 25556 43843
rect 25504 43800 25556 43809
rect 28264 43732 28316 43784
rect 29092 43664 29144 43716
rect 29276 43664 29328 43716
rect 4804 43596 4856 43648
rect 2610 43494 2662 43546
rect 2674 43494 2726 43546
rect 2738 43494 2790 43546
rect 2802 43494 2854 43546
rect 2866 43494 2918 43546
rect 7610 43494 7662 43546
rect 7674 43494 7726 43546
rect 7738 43494 7790 43546
rect 7802 43494 7854 43546
rect 7866 43494 7918 43546
rect 12610 43494 12662 43546
rect 12674 43494 12726 43546
rect 12738 43494 12790 43546
rect 12802 43494 12854 43546
rect 12866 43494 12918 43546
rect 17610 43494 17662 43546
rect 17674 43494 17726 43546
rect 17738 43494 17790 43546
rect 17802 43494 17854 43546
rect 17866 43494 17918 43546
rect 22610 43494 22662 43546
rect 22674 43494 22726 43546
rect 22738 43494 22790 43546
rect 22802 43494 22854 43546
rect 22866 43494 22918 43546
rect 27610 43494 27662 43546
rect 27674 43494 27726 43546
rect 27738 43494 27790 43546
rect 27802 43494 27854 43546
rect 27866 43494 27918 43546
rect 32610 43494 32662 43546
rect 32674 43494 32726 43546
rect 32738 43494 32790 43546
rect 32802 43494 32854 43546
rect 32866 43494 32918 43546
rect 37610 43494 37662 43546
rect 37674 43494 37726 43546
rect 37738 43494 37790 43546
rect 37802 43494 37854 43546
rect 37866 43494 37918 43546
rect 1950 42950 2002 43002
rect 2014 42950 2066 43002
rect 2078 42950 2130 43002
rect 2142 42950 2194 43002
rect 2206 42950 2258 43002
rect 6950 42950 7002 43002
rect 7014 42950 7066 43002
rect 7078 42950 7130 43002
rect 7142 42950 7194 43002
rect 7206 42950 7258 43002
rect 11950 42950 12002 43002
rect 12014 42950 12066 43002
rect 12078 42950 12130 43002
rect 12142 42950 12194 43002
rect 12206 42950 12258 43002
rect 16950 42950 17002 43002
rect 17014 42950 17066 43002
rect 17078 42950 17130 43002
rect 17142 42950 17194 43002
rect 17206 42950 17258 43002
rect 21950 42950 22002 43002
rect 22014 42950 22066 43002
rect 22078 42950 22130 43002
rect 22142 42950 22194 43002
rect 22206 42950 22258 43002
rect 26950 42950 27002 43002
rect 27014 42950 27066 43002
rect 27078 42950 27130 43002
rect 27142 42950 27194 43002
rect 27206 42950 27258 43002
rect 31950 42950 32002 43002
rect 32014 42950 32066 43002
rect 32078 42950 32130 43002
rect 32142 42950 32194 43002
rect 32206 42950 32258 43002
rect 36950 42950 37002 43002
rect 37014 42950 37066 43002
rect 37078 42950 37130 43002
rect 37142 42950 37194 43002
rect 37206 42950 37258 43002
rect 2610 42406 2662 42458
rect 2674 42406 2726 42458
rect 2738 42406 2790 42458
rect 2802 42406 2854 42458
rect 2866 42406 2918 42458
rect 7610 42406 7662 42458
rect 7674 42406 7726 42458
rect 7738 42406 7790 42458
rect 7802 42406 7854 42458
rect 7866 42406 7918 42458
rect 12610 42406 12662 42458
rect 12674 42406 12726 42458
rect 12738 42406 12790 42458
rect 12802 42406 12854 42458
rect 12866 42406 12918 42458
rect 17610 42406 17662 42458
rect 17674 42406 17726 42458
rect 17738 42406 17790 42458
rect 17802 42406 17854 42458
rect 17866 42406 17918 42458
rect 22610 42406 22662 42458
rect 22674 42406 22726 42458
rect 22738 42406 22790 42458
rect 22802 42406 22854 42458
rect 22866 42406 22918 42458
rect 27610 42406 27662 42458
rect 27674 42406 27726 42458
rect 27738 42406 27790 42458
rect 27802 42406 27854 42458
rect 27866 42406 27918 42458
rect 32610 42406 32662 42458
rect 32674 42406 32726 42458
rect 32738 42406 32790 42458
rect 32802 42406 32854 42458
rect 32866 42406 32918 42458
rect 37610 42406 37662 42458
rect 37674 42406 37726 42458
rect 37738 42406 37790 42458
rect 37802 42406 37854 42458
rect 37866 42406 37918 42458
rect 1950 41862 2002 41914
rect 2014 41862 2066 41914
rect 2078 41862 2130 41914
rect 2142 41862 2194 41914
rect 2206 41862 2258 41914
rect 6950 41862 7002 41914
rect 7014 41862 7066 41914
rect 7078 41862 7130 41914
rect 7142 41862 7194 41914
rect 7206 41862 7258 41914
rect 11950 41862 12002 41914
rect 12014 41862 12066 41914
rect 12078 41862 12130 41914
rect 12142 41862 12194 41914
rect 12206 41862 12258 41914
rect 16950 41862 17002 41914
rect 17014 41862 17066 41914
rect 17078 41862 17130 41914
rect 17142 41862 17194 41914
rect 17206 41862 17258 41914
rect 21950 41862 22002 41914
rect 22014 41862 22066 41914
rect 22078 41862 22130 41914
rect 22142 41862 22194 41914
rect 22206 41862 22258 41914
rect 26950 41862 27002 41914
rect 27014 41862 27066 41914
rect 27078 41862 27130 41914
rect 27142 41862 27194 41914
rect 27206 41862 27258 41914
rect 31950 41862 32002 41914
rect 32014 41862 32066 41914
rect 32078 41862 32130 41914
rect 32142 41862 32194 41914
rect 32206 41862 32258 41914
rect 36950 41862 37002 41914
rect 37014 41862 37066 41914
rect 37078 41862 37130 41914
rect 37142 41862 37194 41914
rect 37206 41862 37258 41914
rect 13544 41760 13596 41812
rect 26056 41692 26108 41744
rect 30748 41692 30800 41744
rect 28908 41624 28960 41676
rect 13820 41556 13872 41608
rect 14280 41556 14332 41608
rect 14924 41556 14976 41608
rect 15384 41599 15436 41608
rect 15384 41565 15393 41599
rect 15393 41565 15427 41599
rect 15427 41565 15436 41599
rect 15384 41556 15436 41565
rect 25044 41531 25096 41540
rect 25044 41497 25053 41531
rect 25053 41497 25087 41531
rect 25087 41497 25096 41531
rect 25044 41488 25096 41497
rect 26332 41488 26384 41540
rect 5264 41420 5316 41472
rect 15568 41420 15620 41472
rect 19984 41420 20036 41472
rect 30472 41624 30524 41676
rect 26700 41488 26752 41540
rect 27988 41488 28040 41540
rect 28908 41488 28960 41540
rect 36820 41556 36872 41608
rect 37280 41488 37332 41540
rect 30748 41420 30800 41472
rect 2610 41318 2662 41370
rect 2674 41318 2726 41370
rect 2738 41318 2790 41370
rect 2802 41318 2854 41370
rect 2866 41318 2918 41370
rect 7610 41318 7662 41370
rect 7674 41318 7726 41370
rect 7738 41318 7790 41370
rect 7802 41318 7854 41370
rect 7866 41318 7918 41370
rect 12610 41318 12662 41370
rect 12674 41318 12726 41370
rect 12738 41318 12790 41370
rect 12802 41318 12854 41370
rect 12866 41318 12918 41370
rect 17610 41318 17662 41370
rect 17674 41318 17726 41370
rect 17738 41318 17790 41370
rect 17802 41318 17854 41370
rect 17866 41318 17918 41370
rect 22610 41318 22662 41370
rect 22674 41318 22726 41370
rect 22738 41318 22790 41370
rect 22802 41318 22854 41370
rect 22866 41318 22918 41370
rect 27610 41318 27662 41370
rect 27674 41318 27726 41370
rect 27738 41318 27790 41370
rect 27802 41318 27854 41370
rect 27866 41318 27918 41370
rect 32610 41318 32662 41370
rect 32674 41318 32726 41370
rect 32738 41318 32790 41370
rect 32802 41318 32854 41370
rect 32866 41318 32918 41370
rect 37610 41318 37662 41370
rect 37674 41318 37726 41370
rect 37738 41318 37790 41370
rect 37802 41318 37854 41370
rect 37866 41318 37918 41370
rect 16120 41216 16172 41268
rect 16672 41216 16724 41268
rect 22376 41148 22428 41200
rect 7564 41080 7616 41132
rect 7380 41012 7432 41064
rect 8300 41080 8352 41132
rect 25596 41123 25648 41132
rect 25596 41089 25605 41123
rect 25605 41089 25639 41123
rect 25639 41089 25648 41123
rect 25596 41080 25648 41089
rect 8208 41012 8260 41064
rect 14188 41012 14240 41064
rect 33876 41012 33928 41064
rect 7472 40876 7524 40928
rect 1950 40774 2002 40826
rect 2014 40774 2066 40826
rect 2078 40774 2130 40826
rect 2142 40774 2194 40826
rect 2206 40774 2258 40826
rect 6950 40774 7002 40826
rect 7014 40774 7066 40826
rect 7078 40774 7130 40826
rect 7142 40774 7194 40826
rect 7206 40774 7258 40826
rect 11950 40774 12002 40826
rect 12014 40774 12066 40826
rect 12078 40774 12130 40826
rect 12142 40774 12194 40826
rect 12206 40774 12258 40826
rect 16950 40774 17002 40826
rect 17014 40774 17066 40826
rect 17078 40774 17130 40826
rect 17142 40774 17194 40826
rect 17206 40774 17258 40826
rect 21950 40774 22002 40826
rect 22014 40774 22066 40826
rect 22078 40774 22130 40826
rect 22142 40774 22194 40826
rect 22206 40774 22258 40826
rect 26950 40774 27002 40826
rect 27014 40774 27066 40826
rect 27078 40774 27130 40826
rect 27142 40774 27194 40826
rect 27206 40774 27258 40826
rect 31950 40774 32002 40826
rect 32014 40774 32066 40826
rect 32078 40774 32130 40826
rect 32142 40774 32194 40826
rect 32206 40774 32258 40826
rect 36950 40774 37002 40826
rect 37014 40774 37066 40826
rect 37078 40774 37130 40826
rect 37142 40774 37194 40826
rect 37206 40774 37258 40826
rect 10600 40672 10652 40724
rect 10784 40672 10836 40724
rect 7380 40604 7432 40656
rect 31300 40604 31352 40656
rect 3608 40579 3660 40588
rect 3608 40545 3617 40579
rect 3617 40545 3651 40579
rect 3651 40545 3660 40579
rect 3608 40536 3660 40545
rect 16764 40468 16816 40520
rect 17500 40468 17552 40520
rect 15844 40400 15896 40452
rect 16120 40400 16172 40452
rect 2610 40230 2662 40282
rect 2674 40230 2726 40282
rect 2738 40230 2790 40282
rect 2802 40230 2854 40282
rect 2866 40230 2918 40282
rect 7610 40230 7662 40282
rect 7674 40230 7726 40282
rect 7738 40230 7790 40282
rect 7802 40230 7854 40282
rect 7866 40230 7918 40282
rect 12610 40230 12662 40282
rect 12674 40230 12726 40282
rect 12738 40230 12790 40282
rect 12802 40230 12854 40282
rect 12866 40230 12918 40282
rect 17610 40230 17662 40282
rect 17674 40230 17726 40282
rect 17738 40230 17790 40282
rect 17802 40230 17854 40282
rect 17866 40230 17918 40282
rect 22610 40230 22662 40282
rect 22674 40230 22726 40282
rect 22738 40230 22790 40282
rect 22802 40230 22854 40282
rect 22866 40230 22918 40282
rect 27610 40230 27662 40282
rect 27674 40230 27726 40282
rect 27738 40230 27790 40282
rect 27802 40230 27854 40282
rect 27866 40230 27918 40282
rect 32610 40230 32662 40282
rect 32674 40230 32726 40282
rect 32738 40230 32790 40282
rect 32802 40230 32854 40282
rect 32866 40230 32918 40282
rect 37610 40230 37662 40282
rect 37674 40230 37726 40282
rect 37738 40230 37790 40282
rect 37802 40230 37854 40282
rect 37866 40230 37918 40282
rect 1950 39686 2002 39738
rect 2014 39686 2066 39738
rect 2078 39686 2130 39738
rect 2142 39686 2194 39738
rect 2206 39686 2258 39738
rect 6950 39686 7002 39738
rect 7014 39686 7066 39738
rect 7078 39686 7130 39738
rect 7142 39686 7194 39738
rect 7206 39686 7258 39738
rect 11950 39686 12002 39738
rect 12014 39686 12066 39738
rect 12078 39686 12130 39738
rect 12142 39686 12194 39738
rect 12206 39686 12258 39738
rect 16950 39686 17002 39738
rect 17014 39686 17066 39738
rect 17078 39686 17130 39738
rect 17142 39686 17194 39738
rect 17206 39686 17258 39738
rect 21950 39686 22002 39738
rect 22014 39686 22066 39738
rect 22078 39686 22130 39738
rect 22142 39686 22194 39738
rect 22206 39686 22258 39738
rect 26950 39686 27002 39738
rect 27014 39686 27066 39738
rect 27078 39686 27130 39738
rect 27142 39686 27194 39738
rect 27206 39686 27258 39738
rect 31950 39686 32002 39738
rect 32014 39686 32066 39738
rect 32078 39686 32130 39738
rect 32142 39686 32194 39738
rect 32206 39686 32258 39738
rect 36950 39686 37002 39738
rect 37014 39686 37066 39738
rect 37078 39686 37130 39738
rect 37142 39686 37194 39738
rect 37206 39686 37258 39738
rect 22008 39448 22060 39500
rect 25228 39448 25280 39500
rect 14188 39380 14240 39432
rect 23756 39380 23808 39432
rect 26056 39380 26108 39432
rect 29736 39380 29788 39432
rect 8116 39312 8168 39364
rect 22192 39312 22244 39364
rect 30840 39287 30892 39296
rect 30840 39253 30849 39287
rect 30849 39253 30883 39287
rect 30883 39253 30892 39287
rect 30840 39244 30892 39253
rect 2610 39142 2662 39194
rect 2674 39142 2726 39194
rect 2738 39142 2790 39194
rect 2802 39142 2854 39194
rect 2866 39142 2918 39194
rect 7610 39142 7662 39194
rect 7674 39142 7726 39194
rect 7738 39142 7790 39194
rect 7802 39142 7854 39194
rect 7866 39142 7918 39194
rect 12610 39142 12662 39194
rect 12674 39142 12726 39194
rect 12738 39142 12790 39194
rect 12802 39142 12854 39194
rect 12866 39142 12918 39194
rect 17610 39142 17662 39194
rect 17674 39142 17726 39194
rect 17738 39142 17790 39194
rect 17802 39142 17854 39194
rect 17866 39142 17918 39194
rect 22610 39142 22662 39194
rect 22674 39142 22726 39194
rect 22738 39142 22790 39194
rect 22802 39142 22854 39194
rect 22866 39142 22918 39194
rect 27610 39142 27662 39194
rect 27674 39142 27726 39194
rect 27738 39142 27790 39194
rect 27802 39142 27854 39194
rect 27866 39142 27918 39194
rect 32610 39142 32662 39194
rect 32674 39142 32726 39194
rect 32738 39142 32790 39194
rect 32802 39142 32854 39194
rect 32866 39142 32918 39194
rect 37610 39142 37662 39194
rect 37674 39142 37726 39194
rect 37738 39142 37790 39194
rect 37802 39142 37854 39194
rect 37866 39142 37918 39194
rect 14188 39083 14240 39092
rect 14188 39049 14197 39083
rect 14197 39049 14231 39083
rect 14231 39049 14240 39083
rect 14188 39040 14240 39049
rect 22192 39040 22244 39092
rect 22008 38972 22060 39024
rect 18880 38904 18932 38956
rect 20904 38947 20956 38956
rect 20904 38913 20913 38947
rect 20913 38913 20947 38947
rect 20947 38913 20956 38947
rect 20904 38904 20956 38913
rect 21364 38947 21416 38956
rect 21364 38913 21373 38947
rect 21373 38913 21407 38947
rect 21407 38913 21416 38947
rect 21364 38904 21416 38913
rect 8392 38836 8444 38888
rect 9588 38836 9640 38888
rect 23204 38904 23256 38956
rect 24124 38904 24176 38956
rect 12992 38768 13044 38820
rect 21732 38700 21784 38752
rect 25228 38700 25280 38752
rect 26056 38700 26108 38752
rect 1950 38598 2002 38650
rect 2014 38598 2066 38650
rect 2078 38598 2130 38650
rect 2142 38598 2194 38650
rect 2206 38598 2258 38650
rect 6950 38598 7002 38650
rect 7014 38598 7066 38650
rect 7078 38598 7130 38650
rect 7142 38598 7194 38650
rect 7206 38598 7258 38650
rect 11950 38598 12002 38650
rect 12014 38598 12066 38650
rect 12078 38598 12130 38650
rect 12142 38598 12194 38650
rect 12206 38598 12258 38650
rect 16950 38598 17002 38650
rect 17014 38598 17066 38650
rect 17078 38598 17130 38650
rect 17142 38598 17194 38650
rect 17206 38598 17258 38650
rect 21950 38598 22002 38650
rect 22014 38598 22066 38650
rect 22078 38598 22130 38650
rect 22142 38598 22194 38650
rect 22206 38598 22258 38650
rect 26950 38598 27002 38650
rect 27014 38598 27066 38650
rect 27078 38598 27130 38650
rect 27142 38598 27194 38650
rect 27206 38598 27258 38650
rect 31950 38598 32002 38650
rect 32014 38598 32066 38650
rect 32078 38598 32130 38650
rect 32142 38598 32194 38650
rect 32206 38598 32258 38650
rect 36950 38598 37002 38650
rect 37014 38598 37066 38650
rect 37078 38598 37130 38650
rect 37142 38598 37194 38650
rect 37206 38598 37258 38650
rect 25596 38496 25648 38548
rect 26792 38496 26844 38548
rect 9220 38360 9272 38412
rect 6368 38335 6420 38344
rect 6368 38301 6377 38335
rect 6377 38301 6411 38335
rect 6411 38301 6420 38335
rect 6368 38292 6420 38301
rect 2610 38054 2662 38106
rect 2674 38054 2726 38106
rect 2738 38054 2790 38106
rect 2802 38054 2854 38106
rect 2866 38054 2918 38106
rect 7610 38054 7662 38106
rect 7674 38054 7726 38106
rect 7738 38054 7790 38106
rect 7802 38054 7854 38106
rect 7866 38054 7918 38106
rect 12610 38054 12662 38106
rect 12674 38054 12726 38106
rect 12738 38054 12790 38106
rect 12802 38054 12854 38106
rect 12866 38054 12918 38106
rect 17610 38054 17662 38106
rect 17674 38054 17726 38106
rect 17738 38054 17790 38106
rect 17802 38054 17854 38106
rect 17866 38054 17918 38106
rect 22610 38054 22662 38106
rect 22674 38054 22726 38106
rect 22738 38054 22790 38106
rect 22802 38054 22854 38106
rect 22866 38054 22918 38106
rect 27610 38054 27662 38106
rect 27674 38054 27726 38106
rect 27738 38054 27790 38106
rect 27802 38054 27854 38106
rect 27866 38054 27918 38106
rect 32610 38054 32662 38106
rect 32674 38054 32726 38106
rect 32738 38054 32790 38106
rect 32802 38054 32854 38106
rect 32866 38054 32918 38106
rect 37610 38054 37662 38106
rect 37674 38054 37726 38106
rect 37738 38054 37790 38106
rect 37802 38054 37854 38106
rect 37866 38054 37918 38106
rect 5724 37952 5776 38004
rect 25596 37884 25648 37936
rect 24952 37816 25004 37868
rect 31576 37884 31628 37936
rect 31852 37884 31904 37936
rect 29000 37791 29052 37800
rect 18972 37680 19024 37732
rect 29000 37757 29009 37791
rect 29009 37757 29043 37791
rect 29043 37757 29052 37791
rect 29000 37748 29052 37757
rect 32404 37816 32456 37868
rect 31852 37748 31904 37800
rect 37280 37612 37332 37664
rect 1950 37510 2002 37562
rect 2014 37510 2066 37562
rect 2078 37510 2130 37562
rect 2142 37510 2194 37562
rect 2206 37510 2258 37562
rect 6950 37510 7002 37562
rect 7014 37510 7066 37562
rect 7078 37510 7130 37562
rect 7142 37510 7194 37562
rect 7206 37510 7258 37562
rect 11950 37510 12002 37562
rect 12014 37510 12066 37562
rect 12078 37510 12130 37562
rect 12142 37510 12194 37562
rect 12206 37510 12258 37562
rect 16950 37510 17002 37562
rect 17014 37510 17066 37562
rect 17078 37510 17130 37562
rect 17142 37510 17194 37562
rect 17206 37510 17258 37562
rect 21950 37510 22002 37562
rect 22014 37510 22066 37562
rect 22078 37510 22130 37562
rect 22142 37510 22194 37562
rect 22206 37510 22258 37562
rect 26950 37510 27002 37562
rect 27014 37510 27066 37562
rect 27078 37510 27130 37562
rect 27142 37510 27194 37562
rect 27206 37510 27258 37562
rect 31950 37510 32002 37562
rect 32014 37510 32066 37562
rect 32078 37510 32130 37562
rect 32142 37510 32194 37562
rect 32206 37510 32258 37562
rect 36950 37510 37002 37562
rect 37014 37510 37066 37562
rect 37078 37510 37130 37562
rect 37142 37510 37194 37562
rect 37206 37510 37258 37562
rect 29000 37408 29052 37460
rect 40040 37408 40092 37460
rect 14280 37204 14332 37256
rect 27988 37136 28040 37188
rect 2610 36966 2662 37018
rect 2674 36966 2726 37018
rect 2738 36966 2790 37018
rect 2802 36966 2854 37018
rect 2866 36966 2918 37018
rect 7610 36966 7662 37018
rect 7674 36966 7726 37018
rect 7738 36966 7790 37018
rect 7802 36966 7854 37018
rect 7866 36966 7918 37018
rect 12610 36966 12662 37018
rect 12674 36966 12726 37018
rect 12738 36966 12790 37018
rect 12802 36966 12854 37018
rect 12866 36966 12918 37018
rect 17610 36966 17662 37018
rect 17674 36966 17726 37018
rect 17738 36966 17790 37018
rect 17802 36966 17854 37018
rect 17866 36966 17918 37018
rect 22610 36966 22662 37018
rect 22674 36966 22726 37018
rect 22738 36966 22790 37018
rect 22802 36966 22854 37018
rect 22866 36966 22918 37018
rect 27610 36966 27662 37018
rect 27674 36966 27726 37018
rect 27738 36966 27790 37018
rect 27802 36966 27854 37018
rect 27866 36966 27918 37018
rect 32610 36966 32662 37018
rect 32674 36966 32726 37018
rect 32738 36966 32790 37018
rect 32802 36966 32854 37018
rect 32866 36966 32918 37018
rect 37610 36966 37662 37018
rect 37674 36966 37726 37018
rect 37738 36966 37790 37018
rect 37802 36966 37854 37018
rect 37866 36966 37918 37018
rect 8300 36864 8352 36916
rect 8392 36796 8444 36848
rect 9220 36728 9272 36780
rect 27436 36864 27488 36916
rect 26792 36728 26844 36780
rect 31484 36660 31536 36712
rect 31576 36592 31628 36644
rect 1950 36422 2002 36474
rect 2014 36422 2066 36474
rect 2078 36422 2130 36474
rect 2142 36422 2194 36474
rect 2206 36422 2258 36474
rect 6950 36422 7002 36474
rect 7014 36422 7066 36474
rect 7078 36422 7130 36474
rect 7142 36422 7194 36474
rect 7206 36422 7258 36474
rect 11950 36422 12002 36474
rect 12014 36422 12066 36474
rect 12078 36422 12130 36474
rect 12142 36422 12194 36474
rect 12206 36422 12258 36474
rect 16950 36422 17002 36474
rect 17014 36422 17066 36474
rect 17078 36422 17130 36474
rect 17142 36422 17194 36474
rect 17206 36422 17258 36474
rect 21950 36422 22002 36474
rect 22014 36422 22066 36474
rect 22078 36422 22130 36474
rect 22142 36422 22194 36474
rect 22206 36422 22258 36474
rect 26950 36422 27002 36474
rect 27014 36422 27066 36474
rect 27078 36422 27130 36474
rect 27142 36422 27194 36474
rect 27206 36422 27258 36474
rect 31950 36422 32002 36474
rect 32014 36422 32066 36474
rect 32078 36422 32130 36474
rect 32142 36422 32194 36474
rect 32206 36422 32258 36474
rect 36950 36422 37002 36474
rect 37014 36422 37066 36474
rect 37078 36422 37130 36474
rect 37142 36422 37194 36474
rect 37206 36422 37258 36474
rect 9404 36320 9456 36372
rect 30656 36252 30708 36304
rect 32220 36252 32272 36304
rect 8484 36116 8536 36168
rect 18972 36184 19024 36236
rect 31852 36116 31904 36168
rect 32036 36159 32088 36168
rect 32036 36125 32045 36159
rect 32045 36125 32079 36159
rect 32079 36125 32088 36159
rect 32036 36116 32088 36125
rect 18604 35980 18656 36032
rect 32404 36184 32456 36236
rect 33048 36184 33100 36236
rect 40224 36227 40276 36236
rect 40224 36193 40233 36227
rect 40233 36193 40267 36227
rect 40267 36193 40276 36227
rect 40224 36184 40276 36193
rect 40500 36159 40552 36168
rect 40500 36125 40509 36159
rect 40509 36125 40543 36159
rect 40543 36125 40552 36159
rect 40500 36116 40552 36125
rect 32404 36091 32456 36100
rect 32404 36057 32413 36091
rect 32413 36057 32447 36091
rect 32447 36057 32456 36091
rect 32404 36048 32456 36057
rect 32220 36023 32272 36032
rect 32220 35989 32229 36023
rect 32229 35989 32263 36023
rect 32263 35989 32272 36023
rect 32220 35980 32272 35989
rect 32956 35980 33008 36032
rect 2610 35878 2662 35930
rect 2674 35878 2726 35930
rect 2738 35878 2790 35930
rect 2802 35878 2854 35930
rect 2866 35878 2918 35930
rect 7610 35878 7662 35930
rect 7674 35878 7726 35930
rect 7738 35878 7790 35930
rect 7802 35878 7854 35930
rect 7866 35878 7918 35930
rect 12610 35878 12662 35930
rect 12674 35878 12726 35930
rect 12738 35878 12790 35930
rect 12802 35878 12854 35930
rect 12866 35878 12918 35930
rect 17610 35878 17662 35930
rect 17674 35878 17726 35930
rect 17738 35878 17790 35930
rect 17802 35878 17854 35930
rect 17866 35878 17918 35930
rect 22610 35878 22662 35930
rect 22674 35878 22726 35930
rect 22738 35878 22790 35930
rect 22802 35878 22854 35930
rect 22866 35878 22918 35930
rect 27610 35878 27662 35930
rect 27674 35878 27726 35930
rect 27738 35878 27790 35930
rect 27802 35878 27854 35930
rect 27866 35878 27918 35930
rect 32610 35878 32662 35930
rect 32674 35878 32726 35930
rect 32738 35878 32790 35930
rect 32802 35878 32854 35930
rect 32866 35878 32918 35930
rect 37610 35878 37662 35930
rect 37674 35878 37726 35930
rect 37738 35878 37790 35930
rect 37802 35878 37854 35930
rect 37866 35878 37918 35930
rect 34980 35683 35032 35692
rect 34980 35649 34987 35683
rect 34987 35649 35021 35683
rect 35021 35649 35032 35683
rect 34980 35640 35032 35649
rect 20352 35504 20404 35556
rect 15936 35436 15988 35488
rect 35440 35615 35492 35624
rect 35440 35581 35449 35615
rect 35449 35581 35483 35615
rect 35483 35581 35492 35615
rect 35440 35572 35492 35581
rect 35348 35479 35400 35488
rect 35348 35445 35357 35479
rect 35357 35445 35391 35479
rect 35391 35445 35400 35479
rect 35348 35436 35400 35445
rect 39028 35436 39080 35488
rect 1950 35334 2002 35386
rect 2014 35334 2066 35386
rect 2078 35334 2130 35386
rect 2142 35334 2194 35386
rect 2206 35334 2258 35386
rect 6950 35334 7002 35386
rect 7014 35334 7066 35386
rect 7078 35334 7130 35386
rect 7142 35334 7194 35386
rect 7206 35334 7258 35386
rect 11950 35334 12002 35386
rect 12014 35334 12066 35386
rect 12078 35334 12130 35386
rect 12142 35334 12194 35386
rect 12206 35334 12258 35386
rect 16950 35334 17002 35386
rect 17014 35334 17066 35386
rect 17078 35334 17130 35386
rect 17142 35334 17194 35386
rect 17206 35334 17258 35386
rect 21950 35334 22002 35386
rect 22014 35334 22066 35386
rect 22078 35334 22130 35386
rect 22142 35334 22194 35386
rect 22206 35334 22258 35386
rect 26950 35334 27002 35386
rect 27014 35334 27066 35386
rect 27078 35334 27130 35386
rect 27142 35334 27194 35386
rect 27206 35334 27258 35386
rect 31950 35334 32002 35386
rect 32014 35334 32066 35386
rect 32078 35334 32130 35386
rect 32142 35334 32194 35386
rect 32206 35334 32258 35386
rect 36950 35334 37002 35386
rect 37014 35334 37066 35386
rect 37078 35334 37130 35386
rect 37142 35334 37194 35386
rect 37206 35334 37258 35386
rect 29828 35164 29880 35216
rect 36728 35164 36780 35216
rect 2610 34790 2662 34842
rect 2674 34790 2726 34842
rect 2738 34790 2790 34842
rect 2802 34790 2854 34842
rect 2866 34790 2918 34842
rect 7610 34790 7662 34842
rect 7674 34790 7726 34842
rect 7738 34790 7790 34842
rect 7802 34790 7854 34842
rect 7866 34790 7918 34842
rect 12610 34790 12662 34842
rect 12674 34790 12726 34842
rect 12738 34790 12790 34842
rect 12802 34790 12854 34842
rect 12866 34790 12918 34842
rect 17610 34790 17662 34842
rect 17674 34790 17726 34842
rect 17738 34790 17790 34842
rect 17802 34790 17854 34842
rect 17866 34790 17918 34842
rect 22610 34790 22662 34842
rect 22674 34790 22726 34842
rect 22738 34790 22790 34842
rect 22802 34790 22854 34842
rect 22866 34790 22918 34842
rect 27610 34790 27662 34842
rect 27674 34790 27726 34842
rect 27738 34790 27790 34842
rect 27802 34790 27854 34842
rect 27866 34790 27918 34842
rect 32610 34790 32662 34842
rect 32674 34790 32726 34842
rect 32738 34790 32790 34842
rect 32802 34790 32854 34842
rect 32866 34790 32918 34842
rect 37610 34790 37662 34842
rect 37674 34790 37726 34842
rect 37738 34790 37790 34842
rect 37802 34790 37854 34842
rect 37866 34790 37918 34842
rect 17408 34620 17460 34672
rect 15476 34552 15528 34604
rect 15936 34552 15988 34604
rect 35440 34552 35492 34604
rect 8668 34484 8720 34536
rect 1950 34246 2002 34298
rect 2014 34246 2066 34298
rect 2078 34246 2130 34298
rect 2142 34246 2194 34298
rect 2206 34246 2258 34298
rect 6950 34246 7002 34298
rect 7014 34246 7066 34298
rect 7078 34246 7130 34298
rect 7142 34246 7194 34298
rect 7206 34246 7258 34298
rect 11950 34246 12002 34298
rect 12014 34246 12066 34298
rect 12078 34246 12130 34298
rect 12142 34246 12194 34298
rect 12206 34246 12258 34298
rect 16950 34246 17002 34298
rect 17014 34246 17066 34298
rect 17078 34246 17130 34298
rect 17142 34246 17194 34298
rect 17206 34246 17258 34298
rect 21950 34246 22002 34298
rect 22014 34246 22066 34298
rect 22078 34246 22130 34298
rect 22142 34246 22194 34298
rect 22206 34246 22258 34298
rect 26950 34246 27002 34298
rect 27014 34246 27066 34298
rect 27078 34246 27130 34298
rect 27142 34246 27194 34298
rect 27206 34246 27258 34298
rect 31950 34246 32002 34298
rect 32014 34246 32066 34298
rect 32078 34246 32130 34298
rect 32142 34246 32194 34298
rect 32206 34246 32258 34298
rect 36950 34246 37002 34298
rect 37014 34246 37066 34298
rect 37078 34246 37130 34298
rect 37142 34246 37194 34298
rect 37206 34246 37258 34298
rect 18880 34144 18932 34196
rect 25136 34144 25188 34196
rect 10692 34076 10744 34128
rect 19616 33983 19668 33992
rect 19616 33949 19625 33983
rect 19625 33949 19659 33983
rect 19659 33949 19668 33983
rect 19616 33940 19668 33949
rect 23296 34008 23348 34060
rect 25136 34051 25188 34060
rect 25136 34017 25145 34051
rect 25145 34017 25179 34051
rect 25179 34017 25188 34051
rect 25136 34008 25188 34017
rect 14832 33872 14884 33924
rect 15108 33872 15160 33924
rect 21088 33847 21140 33856
rect 21088 33813 21097 33847
rect 21097 33813 21131 33847
rect 21131 33813 21140 33847
rect 21088 33804 21140 33813
rect 24584 33847 24636 33856
rect 24584 33813 24593 33847
rect 24593 33813 24627 33847
rect 24627 33813 24636 33847
rect 24584 33804 24636 33813
rect 2610 33702 2662 33754
rect 2674 33702 2726 33754
rect 2738 33702 2790 33754
rect 2802 33702 2854 33754
rect 2866 33702 2918 33754
rect 7610 33702 7662 33754
rect 7674 33702 7726 33754
rect 7738 33702 7790 33754
rect 7802 33702 7854 33754
rect 7866 33702 7918 33754
rect 12610 33702 12662 33754
rect 12674 33702 12726 33754
rect 12738 33702 12790 33754
rect 12802 33702 12854 33754
rect 12866 33702 12918 33754
rect 17610 33702 17662 33754
rect 17674 33702 17726 33754
rect 17738 33702 17790 33754
rect 17802 33702 17854 33754
rect 17866 33702 17918 33754
rect 22610 33702 22662 33754
rect 22674 33702 22726 33754
rect 22738 33702 22790 33754
rect 22802 33702 22854 33754
rect 22866 33702 22918 33754
rect 27610 33702 27662 33754
rect 27674 33702 27726 33754
rect 27738 33702 27790 33754
rect 27802 33702 27854 33754
rect 27866 33702 27918 33754
rect 32610 33702 32662 33754
rect 32674 33702 32726 33754
rect 32738 33702 32790 33754
rect 32802 33702 32854 33754
rect 32866 33702 32918 33754
rect 37610 33702 37662 33754
rect 37674 33702 37726 33754
rect 37738 33702 37790 33754
rect 37802 33702 37854 33754
rect 37866 33702 37918 33754
rect 9220 33600 9272 33652
rect 10508 33600 10560 33652
rect 14372 33600 14424 33652
rect 24584 33600 24636 33652
rect 14924 33464 14976 33516
rect 31760 33464 31812 33516
rect 10416 33260 10468 33312
rect 10692 33260 10744 33312
rect 18604 33260 18656 33312
rect 18880 33260 18932 33312
rect 24676 33260 24728 33312
rect 1950 33158 2002 33210
rect 2014 33158 2066 33210
rect 2078 33158 2130 33210
rect 2142 33158 2194 33210
rect 2206 33158 2258 33210
rect 6950 33158 7002 33210
rect 7014 33158 7066 33210
rect 7078 33158 7130 33210
rect 7142 33158 7194 33210
rect 7206 33158 7258 33210
rect 11950 33158 12002 33210
rect 12014 33158 12066 33210
rect 12078 33158 12130 33210
rect 12142 33158 12194 33210
rect 12206 33158 12258 33210
rect 16950 33158 17002 33210
rect 17014 33158 17066 33210
rect 17078 33158 17130 33210
rect 17142 33158 17194 33210
rect 17206 33158 17258 33210
rect 21950 33158 22002 33210
rect 22014 33158 22066 33210
rect 22078 33158 22130 33210
rect 22142 33158 22194 33210
rect 22206 33158 22258 33210
rect 26950 33158 27002 33210
rect 27014 33158 27066 33210
rect 27078 33158 27130 33210
rect 27142 33158 27194 33210
rect 27206 33158 27258 33210
rect 31950 33158 32002 33210
rect 32014 33158 32066 33210
rect 32078 33158 32130 33210
rect 32142 33158 32194 33210
rect 32206 33158 32258 33210
rect 36950 33158 37002 33210
rect 37014 33158 37066 33210
rect 37078 33158 37130 33210
rect 37142 33158 37194 33210
rect 37206 33158 37258 33210
rect 15384 32716 15436 32768
rect 16488 32716 16540 32768
rect 31484 32716 31536 32768
rect 38108 32716 38160 32768
rect 38568 32716 38620 32768
rect 2610 32614 2662 32666
rect 2674 32614 2726 32666
rect 2738 32614 2790 32666
rect 2802 32614 2854 32666
rect 2866 32614 2918 32666
rect 7610 32614 7662 32666
rect 7674 32614 7726 32666
rect 7738 32614 7790 32666
rect 7802 32614 7854 32666
rect 7866 32614 7918 32666
rect 12610 32614 12662 32666
rect 12674 32614 12726 32666
rect 12738 32614 12790 32666
rect 12802 32614 12854 32666
rect 12866 32614 12918 32666
rect 17610 32614 17662 32666
rect 17674 32614 17726 32666
rect 17738 32614 17790 32666
rect 17802 32614 17854 32666
rect 17866 32614 17918 32666
rect 22610 32614 22662 32666
rect 22674 32614 22726 32666
rect 22738 32614 22790 32666
rect 22802 32614 22854 32666
rect 22866 32614 22918 32666
rect 27610 32614 27662 32666
rect 27674 32614 27726 32666
rect 27738 32614 27790 32666
rect 27802 32614 27854 32666
rect 27866 32614 27918 32666
rect 32610 32614 32662 32666
rect 32674 32614 32726 32666
rect 32738 32614 32790 32666
rect 32802 32614 32854 32666
rect 32866 32614 32918 32666
rect 37610 32614 37662 32666
rect 37674 32614 37726 32666
rect 37738 32614 37790 32666
rect 37802 32614 37854 32666
rect 37866 32614 37918 32666
rect 6368 32512 6420 32564
rect 40132 32512 40184 32564
rect 13084 32444 13136 32496
rect 6828 32376 6880 32428
rect 28264 32444 28316 32496
rect 28908 32376 28960 32428
rect 31484 32419 31536 32428
rect 31484 32385 31493 32419
rect 31493 32385 31527 32419
rect 31527 32385 31536 32419
rect 31484 32376 31536 32385
rect 36820 32376 36872 32428
rect 38660 32376 38712 32428
rect 18052 32351 18104 32360
rect 18052 32317 18061 32351
rect 18061 32317 18095 32351
rect 18095 32317 18104 32351
rect 18052 32308 18104 32317
rect 19156 32308 19208 32360
rect 35440 32308 35492 32360
rect 38292 32308 38344 32360
rect 38568 32308 38620 32360
rect 25228 32240 25280 32292
rect 35348 32172 35400 32224
rect 1950 32070 2002 32122
rect 2014 32070 2066 32122
rect 2078 32070 2130 32122
rect 2142 32070 2194 32122
rect 2206 32070 2258 32122
rect 6950 32070 7002 32122
rect 7014 32070 7066 32122
rect 7078 32070 7130 32122
rect 7142 32070 7194 32122
rect 7206 32070 7258 32122
rect 11950 32070 12002 32122
rect 12014 32070 12066 32122
rect 12078 32070 12130 32122
rect 12142 32070 12194 32122
rect 12206 32070 12258 32122
rect 16950 32070 17002 32122
rect 17014 32070 17066 32122
rect 17078 32070 17130 32122
rect 17142 32070 17194 32122
rect 17206 32070 17258 32122
rect 21950 32070 22002 32122
rect 22014 32070 22066 32122
rect 22078 32070 22130 32122
rect 22142 32070 22194 32122
rect 22206 32070 22258 32122
rect 26950 32070 27002 32122
rect 27014 32070 27066 32122
rect 27078 32070 27130 32122
rect 27142 32070 27194 32122
rect 27206 32070 27258 32122
rect 31950 32070 32002 32122
rect 32014 32070 32066 32122
rect 32078 32070 32130 32122
rect 32142 32070 32194 32122
rect 32206 32070 32258 32122
rect 36950 32070 37002 32122
rect 37014 32070 37066 32122
rect 37078 32070 37130 32122
rect 37142 32070 37194 32122
rect 37206 32070 37258 32122
rect 24216 31968 24268 32020
rect 39488 31968 39540 32020
rect 39672 31968 39724 32020
rect 40132 31968 40184 32020
rect 6184 31900 6236 31952
rect 28724 31900 28776 31952
rect 25412 31875 25464 31884
rect 25412 31841 25421 31875
rect 25421 31841 25455 31875
rect 25455 31841 25464 31875
rect 25412 31832 25464 31841
rect 35440 31832 35492 31884
rect 20904 31764 20956 31816
rect 21364 31764 21416 31816
rect 25228 31807 25280 31816
rect 25228 31773 25237 31807
rect 25237 31773 25271 31807
rect 25271 31773 25280 31807
rect 25228 31764 25280 31773
rect 29828 31764 29880 31816
rect 7380 31696 7432 31748
rect 29460 31696 29512 31748
rect 34888 31764 34940 31816
rect 36452 31832 36504 31884
rect 36544 31807 36596 31816
rect 36544 31773 36553 31807
rect 36553 31773 36587 31807
rect 36587 31773 36596 31807
rect 36544 31764 36596 31773
rect 39764 31764 39816 31816
rect 2610 31526 2662 31578
rect 2674 31526 2726 31578
rect 2738 31526 2790 31578
rect 2802 31526 2854 31578
rect 2866 31526 2918 31578
rect 7610 31526 7662 31578
rect 7674 31526 7726 31578
rect 7738 31526 7790 31578
rect 7802 31526 7854 31578
rect 7866 31526 7918 31578
rect 12610 31526 12662 31578
rect 12674 31526 12726 31578
rect 12738 31526 12790 31578
rect 12802 31526 12854 31578
rect 12866 31526 12918 31578
rect 17610 31526 17662 31578
rect 17674 31526 17726 31578
rect 17738 31526 17790 31578
rect 17802 31526 17854 31578
rect 17866 31526 17918 31578
rect 22610 31526 22662 31578
rect 22674 31526 22726 31578
rect 22738 31526 22790 31578
rect 22802 31526 22854 31578
rect 22866 31526 22918 31578
rect 27610 31526 27662 31578
rect 27674 31526 27726 31578
rect 27738 31526 27790 31578
rect 27802 31526 27854 31578
rect 27866 31526 27918 31578
rect 32610 31526 32662 31578
rect 32674 31526 32726 31578
rect 32738 31526 32790 31578
rect 32802 31526 32854 31578
rect 32866 31526 32918 31578
rect 37610 31526 37662 31578
rect 37674 31526 37726 31578
rect 37738 31526 37790 31578
rect 37802 31526 37854 31578
rect 37866 31526 37918 31578
rect 14648 31424 14700 31476
rect 17408 31424 17460 31476
rect 19616 31356 19668 31408
rect 7380 31331 7432 31340
rect 7380 31297 7389 31331
rect 7389 31297 7423 31331
rect 7423 31297 7432 31331
rect 7380 31288 7432 31297
rect 8208 31288 8260 31340
rect 18144 31220 18196 31272
rect 2412 31152 2464 31204
rect 20904 31263 20956 31272
rect 20904 31229 20913 31263
rect 20913 31229 20947 31263
rect 20947 31229 20956 31263
rect 20904 31220 20956 31229
rect 31576 31424 31628 31476
rect 33600 31356 33652 31408
rect 31852 31220 31904 31272
rect 33232 31152 33284 31204
rect 16580 31084 16632 31136
rect 29460 31084 29512 31136
rect 33508 31084 33560 31136
rect 1950 30982 2002 31034
rect 2014 30982 2066 31034
rect 2078 30982 2130 31034
rect 2142 30982 2194 31034
rect 2206 30982 2258 31034
rect 6950 30982 7002 31034
rect 7014 30982 7066 31034
rect 7078 30982 7130 31034
rect 7142 30982 7194 31034
rect 7206 30982 7258 31034
rect 11950 30982 12002 31034
rect 12014 30982 12066 31034
rect 12078 30982 12130 31034
rect 12142 30982 12194 31034
rect 12206 30982 12258 31034
rect 16950 30982 17002 31034
rect 17014 30982 17066 31034
rect 17078 30982 17130 31034
rect 17142 30982 17194 31034
rect 17206 30982 17258 31034
rect 21950 30982 22002 31034
rect 22014 30982 22066 31034
rect 22078 30982 22130 31034
rect 22142 30982 22194 31034
rect 22206 30982 22258 31034
rect 26950 30982 27002 31034
rect 27014 30982 27066 31034
rect 27078 30982 27130 31034
rect 27142 30982 27194 31034
rect 27206 30982 27258 31034
rect 31950 30982 32002 31034
rect 32014 30982 32066 31034
rect 32078 30982 32130 31034
rect 32142 30982 32194 31034
rect 32206 30982 32258 31034
rect 36950 30982 37002 31034
rect 37014 30982 37066 31034
rect 37078 30982 37130 31034
rect 37142 30982 37194 31034
rect 37206 30982 37258 31034
rect 9036 30855 9088 30864
rect 9036 30821 9045 30855
rect 9045 30821 9079 30855
rect 9079 30821 9088 30855
rect 9036 30812 9088 30821
rect 14096 30880 14148 30932
rect 14556 30812 14608 30864
rect 21180 30812 21232 30864
rect 9496 30744 9548 30796
rect 11612 30744 11664 30796
rect 6460 30608 6512 30660
rect 5632 30540 5684 30592
rect 6276 30540 6328 30592
rect 33232 30676 33284 30728
rect 34152 30676 34204 30728
rect 11336 30608 11388 30660
rect 40040 30651 40092 30660
rect 40040 30617 40049 30651
rect 40049 30617 40083 30651
rect 40083 30617 40092 30651
rect 40040 30608 40092 30617
rect 2610 30438 2662 30490
rect 2674 30438 2726 30490
rect 2738 30438 2790 30490
rect 2802 30438 2854 30490
rect 2866 30438 2918 30490
rect 7610 30438 7662 30490
rect 7674 30438 7726 30490
rect 7738 30438 7790 30490
rect 7802 30438 7854 30490
rect 7866 30438 7918 30490
rect 12610 30438 12662 30490
rect 12674 30438 12726 30490
rect 12738 30438 12790 30490
rect 12802 30438 12854 30490
rect 12866 30438 12918 30490
rect 17610 30438 17662 30490
rect 17674 30438 17726 30490
rect 17738 30438 17790 30490
rect 17802 30438 17854 30490
rect 17866 30438 17918 30490
rect 22610 30438 22662 30490
rect 22674 30438 22726 30490
rect 22738 30438 22790 30490
rect 22802 30438 22854 30490
rect 22866 30438 22918 30490
rect 27610 30438 27662 30490
rect 27674 30438 27726 30490
rect 27738 30438 27790 30490
rect 27802 30438 27854 30490
rect 27866 30438 27918 30490
rect 32610 30438 32662 30490
rect 32674 30438 32726 30490
rect 32738 30438 32790 30490
rect 32802 30438 32854 30490
rect 32866 30438 32918 30490
rect 37610 30438 37662 30490
rect 37674 30438 37726 30490
rect 37738 30438 37790 30490
rect 37802 30438 37854 30490
rect 37866 30438 37918 30490
rect 3056 30336 3108 30388
rect 11336 30336 11388 30388
rect 11520 30268 11572 30320
rect 22468 30268 22520 30320
rect 23020 30268 23072 30320
rect 32404 30268 32456 30320
rect 11704 30243 11756 30252
rect 11704 30209 11713 30243
rect 11713 30209 11747 30243
rect 11747 30209 11756 30243
rect 11704 30200 11756 30209
rect 5080 30132 5132 30184
rect 18880 30200 18932 30252
rect 18604 30132 18656 30184
rect 18788 30132 18840 30184
rect 28632 30064 28684 30116
rect 16856 29996 16908 30048
rect 18420 30039 18472 30048
rect 18420 30005 18429 30039
rect 18429 30005 18463 30039
rect 18463 30005 18472 30039
rect 18420 29996 18472 30005
rect 29000 29996 29052 30048
rect 29276 29996 29328 30048
rect 1950 29894 2002 29946
rect 2014 29894 2066 29946
rect 2078 29894 2130 29946
rect 2142 29894 2194 29946
rect 2206 29894 2258 29946
rect 6950 29894 7002 29946
rect 7014 29894 7066 29946
rect 7078 29894 7130 29946
rect 7142 29894 7194 29946
rect 7206 29894 7258 29946
rect 11950 29894 12002 29946
rect 12014 29894 12066 29946
rect 12078 29894 12130 29946
rect 12142 29894 12194 29946
rect 12206 29894 12258 29946
rect 16950 29894 17002 29946
rect 17014 29894 17066 29946
rect 17078 29894 17130 29946
rect 17142 29894 17194 29946
rect 17206 29894 17258 29946
rect 21950 29894 22002 29946
rect 22014 29894 22066 29946
rect 22078 29894 22130 29946
rect 22142 29894 22194 29946
rect 22206 29894 22258 29946
rect 26950 29894 27002 29946
rect 27014 29894 27066 29946
rect 27078 29894 27130 29946
rect 27142 29894 27194 29946
rect 27206 29894 27258 29946
rect 31950 29894 32002 29946
rect 32014 29894 32066 29946
rect 32078 29894 32130 29946
rect 32142 29894 32194 29946
rect 32206 29894 32258 29946
rect 36950 29894 37002 29946
rect 37014 29894 37066 29946
rect 37078 29894 37130 29946
rect 37142 29894 37194 29946
rect 37206 29894 37258 29946
rect 3976 29792 4028 29844
rect 8484 29792 8536 29844
rect 17408 29792 17460 29844
rect 18420 29792 18472 29844
rect 31024 29792 31076 29844
rect 3884 29656 3936 29708
rect 11612 29656 11664 29708
rect 6184 29588 6236 29640
rect 8300 29631 8352 29640
rect 8300 29597 8309 29631
rect 8309 29597 8343 29631
rect 8343 29597 8352 29631
rect 14188 29656 14240 29708
rect 14280 29656 14332 29708
rect 8300 29588 8352 29597
rect 13912 29588 13964 29640
rect 6092 29520 6144 29572
rect 15292 29588 15344 29640
rect 6460 29452 6512 29504
rect 8484 29452 8536 29504
rect 2610 29350 2662 29402
rect 2674 29350 2726 29402
rect 2738 29350 2790 29402
rect 2802 29350 2854 29402
rect 2866 29350 2918 29402
rect 7610 29350 7662 29402
rect 7674 29350 7726 29402
rect 7738 29350 7790 29402
rect 7802 29350 7854 29402
rect 7866 29350 7918 29402
rect 12610 29350 12662 29402
rect 12674 29350 12726 29402
rect 12738 29350 12790 29402
rect 12802 29350 12854 29402
rect 12866 29350 12918 29402
rect 17610 29350 17662 29402
rect 17674 29350 17726 29402
rect 17738 29350 17790 29402
rect 17802 29350 17854 29402
rect 17866 29350 17918 29402
rect 22610 29350 22662 29402
rect 22674 29350 22726 29402
rect 22738 29350 22790 29402
rect 22802 29350 22854 29402
rect 22866 29350 22918 29402
rect 27610 29350 27662 29402
rect 27674 29350 27726 29402
rect 27738 29350 27790 29402
rect 27802 29350 27854 29402
rect 27866 29350 27918 29402
rect 32610 29350 32662 29402
rect 32674 29350 32726 29402
rect 32738 29350 32790 29402
rect 32802 29350 32854 29402
rect 32866 29350 32918 29402
rect 37610 29350 37662 29402
rect 37674 29350 37726 29402
rect 37738 29350 37790 29402
rect 37802 29350 37854 29402
rect 37866 29350 37918 29402
rect 15384 29248 15436 29300
rect 14464 29180 14516 29232
rect 33692 29248 33744 29300
rect 3884 29155 3936 29164
rect 3884 29121 3893 29155
rect 3893 29121 3927 29155
rect 3927 29121 3936 29155
rect 3884 29112 3936 29121
rect 5264 29112 5316 29164
rect 7380 29112 7432 29164
rect 12440 29112 12492 29164
rect 16856 29112 16908 29164
rect 17960 29180 18012 29232
rect 18420 29180 18472 29232
rect 18512 29223 18564 29232
rect 18512 29189 18521 29223
rect 18521 29189 18555 29223
rect 18555 29189 18564 29223
rect 18512 29180 18564 29189
rect 20720 29180 20772 29232
rect 23020 29112 23072 29164
rect 40224 29112 40276 29164
rect 4804 29044 4856 29096
rect 6460 29087 6512 29096
rect 6460 29053 6469 29087
rect 6469 29053 6503 29087
rect 6503 29053 6512 29087
rect 6460 29044 6512 29053
rect 18144 29044 18196 29096
rect 19524 28976 19576 29028
rect 26792 29044 26844 29096
rect 1950 28806 2002 28858
rect 2014 28806 2066 28858
rect 2078 28806 2130 28858
rect 2142 28806 2194 28858
rect 2206 28806 2258 28858
rect 6950 28806 7002 28858
rect 7014 28806 7066 28858
rect 7078 28806 7130 28858
rect 7142 28806 7194 28858
rect 7206 28806 7258 28858
rect 11950 28806 12002 28858
rect 12014 28806 12066 28858
rect 12078 28806 12130 28858
rect 12142 28806 12194 28858
rect 12206 28806 12258 28858
rect 16950 28806 17002 28858
rect 17014 28806 17066 28858
rect 17078 28806 17130 28858
rect 17142 28806 17194 28858
rect 17206 28806 17258 28858
rect 21950 28806 22002 28858
rect 22014 28806 22066 28858
rect 22078 28806 22130 28858
rect 22142 28806 22194 28858
rect 22206 28806 22258 28858
rect 26950 28806 27002 28858
rect 27014 28806 27066 28858
rect 27078 28806 27130 28858
rect 27142 28806 27194 28858
rect 27206 28806 27258 28858
rect 31950 28806 32002 28858
rect 32014 28806 32066 28858
rect 32078 28806 32130 28858
rect 32142 28806 32194 28858
rect 32206 28806 32258 28858
rect 36950 28806 37002 28858
rect 37014 28806 37066 28858
rect 37078 28806 37130 28858
rect 37142 28806 37194 28858
rect 37206 28806 37258 28858
rect 17960 28636 18012 28688
rect 19156 28636 19208 28688
rect 19984 28568 20036 28620
rect 8300 28500 8352 28552
rect 11520 28500 11572 28552
rect 11704 28432 11756 28484
rect 19800 28543 19852 28552
rect 19800 28509 19809 28543
rect 19809 28509 19843 28543
rect 19843 28509 19852 28543
rect 19800 28500 19852 28509
rect 30564 28679 30616 28688
rect 30564 28645 30573 28679
rect 30573 28645 30607 28679
rect 30607 28645 30616 28679
rect 30564 28636 30616 28645
rect 29460 28568 29512 28620
rect 33600 28568 33652 28620
rect 8208 28364 8260 28416
rect 8300 28364 8352 28416
rect 17960 28364 18012 28416
rect 19340 28407 19392 28416
rect 19340 28373 19349 28407
rect 19349 28373 19383 28407
rect 19383 28373 19392 28407
rect 19340 28364 19392 28373
rect 22008 28432 22060 28484
rect 31576 28500 31628 28552
rect 31852 28432 31904 28484
rect 19800 28364 19852 28416
rect 20444 28364 20496 28416
rect 2610 28262 2662 28314
rect 2674 28262 2726 28314
rect 2738 28262 2790 28314
rect 2802 28262 2854 28314
rect 2866 28262 2918 28314
rect 7610 28262 7662 28314
rect 7674 28262 7726 28314
rect 7738 28262 7790 28314
rect 7802 28262 7854 28314
rect 7866 28262 7918 28314
rect 12610 28262 12662 28314
rect 12674 28262 12726 28314
rect 12738 28262 12790 28314
rect 12802 28262 12854 28314
rect 12866 28262 12918 28314
rect 17610 28262 17662 28314
rect 17674 28262 17726 28314
rect 17738 28262 17790 28314
rect 17802 28262 17854 28314
rect 17866 28262 17918 28314
rect 22610 28262 22662 28314
rect 22674 28262 22726 28314
rect 22738 28262 22790 28314
rect 22802 28262 22854 28314
rect 22866 28262 22918 28314
rect 27610 28262 27662 28314
rect 27674 28262 27726 28314
rect 27738 28262 27790 28314
rect 27802 28262 27854 28314
rect 27866 28262 27918 28314
rect 32610 28262 32662 28314
rect 32674 28262 32726 28314
rect 32738 28262 32790 28314
rect 32802 28262 32854 28314
rect 32866 28262 32918 28314
rect 37610 28262 37662 28314
rect 37674 28262 37726 28314
rect 37738 28262 37790 28314
rect 37802 28262 37854 28314
rect 37866 28262 37918 28314
rect 29092 28160 29144 28212
rect 29552 28203 29604 28212
rect 29552 28169 29561 28203
rect 29561 28169 29595 28203
rect 29595 28169 29604 28203
rect 29552 28160 29604 28169
rect 31852 28160 31904 28212
rect 32404 28160 32456 28212
rect 17500 28092 17552 28144
rect 29276 28092 29328 28144
rect 20444 28024 20496 28076
rect 22008 28067 22060 28076
rect 22008 28033 22017 28067
rect 22017 28033 22051 28067
rect 22051 28033 22060 28067
rect 22008 28024 22060 28033
rect 9864 27888 9916 27940
rect 10600 27888 10652 27940
rect 29092 28024 29144 28076
rect 38568 27888 38620 27940
rect 29092 27820 29144 27872
rect 1950 27718 2002 27770
rect 2014 27718 2066 27770
rect 2078 27718 2130 27770
rect 2142 27718 2194 27770
rect 2206 27718 2258 27770
rect 6950 27718 7002 27770
rect 7014 27718 7066 27770
rect 7078 27718 7130 27770
rect 7142 27718 7194 27770
rect 7206 27718 7258 27770
rect 11950 27718 12002 27770
rect 12014 27718 12066 27770
rect 12078 27718 12130 27770
rect 12142 27718 12194 27770
rect 12206 27718 12258 27770
rect 16950 27718 17002 27770
rect 17014 27718 17066 27770
rect 17078 27718 17130 27770
rect 17142 27718 17194 27770
rect 17206 27718 17258 27770
rect 21950 27718 22002 27770
rect 22014 27718 22066 27770
rect 22078 27718 22130 27770
rect 22142 27718 22194 27770
rect 22206 27718 22258 27770
rect 26950 27718 27002 27770
rect 27014 27718 27066 27770
rect 27078 27718 27130 27770
rect 27142 27718 27194 27770
rect 27206 27718 27258 27770
rect 31950 27718 32002 27770
rect 32014 27718 32066 27770
rect 32078 27718 32130 27770
rect 32142 27718 32194 27770
rect 32206 27718 32258 27770
rect 36950 27718 37002 27770
rect 37014 27718 37066 27770
rect 37078 27718 37130 27770
rect 37142 27718 37194 27770
rect 37206 27718 37258 27770
rect 22468 27616 22520 27668
rect 19984 27548 20036 27600
rect 29000 27548 29052 27600
rect 31668 27548 31720 27600
rect 12348 27480 12400 27532
rect 18144 27412 18196 27464
rect 19984 27455 20036 27464
rect 19984 27421 19993 27455
rect 19993 27421 20027 27455
rect 20027 27421 20036 27455
rect 19984 27412 20036 27421
rect 20444 27523 20496 27532
rect 20444 27489 20453 27523
rect 20453 27489 20487 27523
rect 20487 27489 20496 27523
rect 20444 27480 20496 27489
rect 15844 27387 15896 27396
rect 15844 27353 15853 27387
rect 15853 27353 15887 27387
rect 15887 27353 15896 27387
rect 15844 27344 15896 27353
rect 32496 27344 32548 27396
rect 38016 27276 38068 27328
rect 2610 27174 2662 27226
rect 2674 27174 2726 27226
rect 2738 27174 2790 27226
rect 2802 27174 2854 27226
rect 2866 27174 2918 27226
rect 7610 27174 7662 27226
rect 7674 27174 7726 27226
rect 7738 27174 7790 27226
rect 7802 27174 7854 27226
rect 7866 27174 7918 27226
rect 12610 27174 12662 27226
rect 12674 27174 12726 27226
rect 12738 27174 12790 27226
rect 12802 27174 12854 27226
rect 12866 27174 12918 27226
rect 17610 27174 17662 27226
rect 17674 27174 17726 27226
rect 17738 27174 17790 27226
rect 17802 27174 17854 27226
rect 17866 27174 17918 27226
rect 22610 27174 22662 27226
rect 22674 27174 22726 27226
rect 22738 27174 22790 27226
rect 22802 27174 22854 27226
rect 22866 27174 22918 27226
rect 27610 27174 27662 27226
rect 27674 27174 27726 27226
rect 27738 27174 27790 27226
rect 27802 27174 27854 27226
rect 27866 27174 27918 27226
rect 32610 27174 32662 27226
rect 32674 27174 32726 27226
rect 32738 27174 32790 27226
rect 32802 27174 32854 27226
rect 32866 27174 32918 27226
rect 37610 27174 37662 27226
rect 37674 27174 37726 27226
rect 37738 27174 37790 27226
rect 37802 27174 37854 27226
rect 37866 27174 37918 27226
rect 8392 27072 8444 27124
rect 14280 27072 14332 27124
rect 19984 27072 20036 27124
rect 18052 27004 18104 27056
rect 8668 26936 8720 26988
rect 9220 26775 9272 26784
rect 9220 26741 9229 26775
rect 9229 26741 9263 26775
rect 9263 26741 9272 26775
rect 9220 26732 9272 26741
rect 1950 26630 2002 26682
rect 2014 26630 2066 26682
rect 2078 26630 2130 26682
rect 2142 26630 2194 26682
rect 2206 26630 2258 26682
rect 6950 26630 7002 26682
rect 7014 26630 7066 26682
rect 7078 26630 7130 26682
rect 7142 26630 7194 26682
rect 7206 26630 7258 26682
rect 11950 26630 12002 26682
rect 12014 26630 12066 26682
rect 12078 26630 12130 26682
rect 12142 26630 12194 26682
rect 12206 26630 12258 26682
rect 16950 26630 17002 26682
rect 17014 26630 17066 26682
rect 17078 26630 17130 26682
rect 17142 26630 17194 26682
rect 17206 26630 17258 26682
rect 21950 26630 22002 26682
rect 22014 26630 22066 26682
rect 22078 26630 22130 26682
rect 22142 26630 22194 26682
rect 22206 26630 22258 26682
rect 26950 26630 27002 26682
rect 27014 26630 27066 26682
rect 27078 26630 27130 26682
rect 27142 26630 27194 26682
rect 27206 26630 27258 26682
rect 31950 26630 32002 26682
rect 32014 26630 32066 26682
rect 32078 26630 32130 26682
rect 32142 26630 32194 26682
rect 32206 26630 32258 26682
rect 36950 26630 37002 26682
rect 37014 26630 37066 26682
rect 37078 26630 37130 26682
rect 37142 26630 37194 26682
rect 37206 26630 37258 26682
rect 2610 26086 2662 26138
rect 2674 26086 2726 26138
rect 2738 26086 2790 26138
rect 2802 26086 2854 26138
rect 2866 26086 2918 26138
rect 7610 26086 7662 26138
rect 7674 26086 7726 26138
rect 7738 26086 7790 26138
rect 7802 26086 7854 26138
rect 7866 26086 7918 26138
rect 12610 26086 12662 26138
rect 12674 26086 12726 26138
rect 12738 26086 12790 26138
rect 12802 26086 12854 26138
rect 12866 26086 12918 26138
rect 17610 26086 17662 26138
rect 17674 26086 17726 26138
rect 17738 26086 17790 26138
rect 17802 26086 17854 26138
rect 17866 26086 17918 26138
rect 22610 26086 22662 26138
rect 22674 26086 22726 26138
rect 22738 26086 22790 26138
rect 22802 26086 22854 26138
rect 22866 26086 22918 26138
rect 27610 26086 27662 26138
rect 27674 26086 27726 26138
rect 27738 26086 27790 26138
rect 27802 26086 27854 26138
rect 27866 26086 27918 26138
rect 32610 26086 32662 26138
rect 32674 26086 32726 26138
rect 32738 26086 32790 26138
rect 32802 26086 32854 26138
rect 32866 26086 32918 26138
rect 37610 26086 37662 26138
rect 37674 26086 37726 26138
rect 37738 26086 37790 26138
rect 37802 26086 37854 26138
rect 37866 26086 37918 26138
rect 36636 25984 36688 26036
rect 31852 25916 31904 25968
rect 32956 25848 33008 25900
rect 33048 25780 33100 25832
rect 32312 25712 32364 25764
rect 1950 25542 2002 25594
rect 2014 25542 2066 25594
rect 2078 25542 2130 25594
rect 2142 25542 2194 25594
rect 2206 25542 2258 25594
rect 6950 25542 7002 25594
rect 7014 25542 7066 25594
rect 7078 25542 7130 25594
rect 7142 25542 7194 25594
rect 7206 25542 7258 25594
rect 11950 25542 12002 25594
rect 12014 25542 12066 25594
rect 12078 25542 12130 25594
rect 12142 25542 12194 25594
rect 12206 25542 12258 25594
rect 16950 25542 17002 25594
rect 17014 25542 17066 25594
rect 17078 25542 17130 25594
rect 17142 25542 17194 25594
rect 17206 25542 17258 25594
rect 21950 25542 22002 25594
rect 22014 25542 22066 25594
rect 22078 25542 22130 25594
rect 22142 25542 22194 25594
rect 22206 25542 22258 25594
rect 26950 25542 27002 25594
rect 27014 25542 27066 25594
rect 27078 25542 27130 25594
rect 27142 25542 27194 25594
rect 27206 25542 27258 25594
rect 31950 25542 32002 25594
rect 32014 25542 32066 25594
rect 32078 25542 32130 25594
rect 32142 25542 32194 25594
rect 32206 25542 32258 25594
rect 36950 25542 37002 25594
rect 37014 25542 37066 25594
rect 37078 25542 37130 25594
rect 37142 25542 37194 25594
rect 37206 25542 37258 25594
rect 9588 25440 9640 25492
rect 11612 25304 11664 25356
rect 14096 25304 14148 25356
rect 14832 25304 14884 25356
rect 15844 25304 15896 25356
rect 26148 25168 26200 25220
rect 29368 25236 29420 25288
rect 29092 25211 29144 25220
rect 29092 25177 29101 25211
rect 29101 25177 29135 25211
rect 29135 25177 29144 25211
rect 29092 25168 29144 25177
rect 29000 25143 29052 25152
rect 29000 25109 29009 25143
rect 29009 25109 29043 25143
rect 29043 25109 29052 25143
rect 29000 25100 29052 25109
rect 29276 25100 29328 25152
rect 2610 24998 2662 25050
rect 2674 24998 2726 25050
rect 2738 24998 2790 25050
rect 2802 24998 2854 25050
rect 2866 24998 2918 25050
rect 7610 24998 7662 25050
rect 7674 24998 7726 25050
rect 7738 24998 7790 25050
rect 7802 24998 7854 25050
rect 7866 24998 7918 25050
rect 12610 24998 12662 25050
rect 12674 24998 12726 25050
rect 12738 24998 12790 25050
rect 12802 24998 12854 25050
rect 12866 24998 12918 25050
rect 17610 24998 17662 25050
rect 17674 24998 17726 25050
rect 17738 24998 17790 25050
rect 17802 24998 17854 25050
rect 17866 24998 17918 25050
rect 22610 24998 22662 25050
rect 22674 24998 22726 25050
rect 22738 24998 22790 25050
rect 22802 24998 22854 25050
rect 22866 24998 22918 25050
rect 27610 24998 27662 25050
rect 27674 24998 27726 25050
rect 27738 24998 27790 25050
rect 27802 24998 27854 25050
rect 27866 24998 27918 25050
rect 32610 24998 32662 25050
rect 32674 24998 32726 25050
rect 32738 24998 32790 25050
rect 32802 24998 32854 25050
rect 32866 24998 32918 25050
rect 37610 24998 37662 25050
rect 37674 24998 37726 25050
rect 37738 24998 37790 25050
rect 37802 24998 37854 25050
rect 37866 24998 37918 25050
rect 24216 24828 24268 24880
rect 5724 24760 5776 24812
rect 6736 24760 6788 24812
rect 18144 24760 18196 24812
rect 23480 24803 23532 24812
rect 23480 24769 23489 24803
rect 23489 24769 23523 24803
rect 23523 24769 23532 24803
rect 23480 24760 23532 24769
rect 23020 24692 23072 24744
rect 6736 24556 6788 24608
rect 31208 24692 31260 24744
rect 1950 24454 2002 24506
rect 2014 24454 2066 24506
rect 2078 24454 2130 24506
rect 2142 24454 2194 24506
rect 2206 24454 2258 24506
rect 6950 24454 7002 24506
rect 7014 24454 7066 24506
rect 7078 24454 7130 24506
rect 7142 24454 7194 24506
rect 7206 24454 7258 24506
rect 11950 24454 12002 24506
rect 12014 24454 12066 24506
rect 12078 24454 12130 24506
rect 12142 24454 12194 24506
rect 12206 24454 12258 24506
rect 16950 24454 17002 24506
rect 17014 24454 17066 24506
rect 17078 24454 17130 24506
rect 17142 24454 17194 24506
rect 17206 24454 17258 24506
rect 21950 24454 22002 24506
rect 22014 24454 22066 24506
rect 22078 24454 22130 24506
rect 22142 24454 22194 24506
rect 22206 24454 22258 24506
rect 26950 24454 27002 24506
rect 27014 24454 27066 24506
rect 27078 24454 27130 24506
rect 27142 24454 27194 24506
rect 27206 24454 27258 24506
rect 31950 24454 32002 24506
rect 32014 24454 32066 24506
rect 32078 24454 32130 24506
rect 32142 24454 32194 24506
rect 32206 24454 32258 24506
rect 36950 24454 37002 24506
rect 37014 24454 37066 24506
rect 37078 24454 37130 24506
rect 37142 24454 37194 24506
rect 37206 24454 37258 24506
rect 15568 24352 15620 24404
rect 24216 24352 24268 24404
rect 27344 24284 27396 24336
rect 24124 24216 24176 24268
rect 3424 24148 3476 24200
rect 14280 24080 14332 24132
rect 14556 24080 14608 24132
rect 34888 24191 34940 24200
rect 34888 24157 34897 24191
rect 34897 24157 34931 24191
rect 34931 24157 34940 24191
rect 34888 24148 34940 24157
rect 2610 23910 2662 23962
rect 2674 23910 2726 23962
rect 2738 23910 2790 23962
rect 2802 23910 2854 23962
rect 2866 23910 2918 23962
rect 7610 23910 7662 23962
rect 7674 23910 7726 23962
rect 7738 23910 7790 23962
rect 7802 23910 7854 23962
rect 7866 23910 7918 23962
rect 12610 23910 12662 23962
rect 12674 23910 12726 23962
rect 12738 23910 12790 23962
rect 12802 23910 12854 23962
rect 12866 23910 12918 23962
rect 17610 23910 17662 23962
rect 17674 23910 17726 23962
rect 17738 23910 17790 23962
rect 17802 23910 17854 23962
rect 17866 23910 17918 23962
rect 22610 23910 22662 23962
rect 22674 23910 22726 23962
rect 22738 23910 22790 23962
rect 22802 23910 22854 23962
rect 22866 23910 22918 23962
rect 27610 23910 27662 23962
rect 27674 23910 27726 23962
rect 27738 23910 27790 23962
rect 27802 23910 27854 23962
rect 27866 23910 27918 23962
rect 32610 23910 32662 23962
rect 32674 23910 32726 23962
rect 32738 23910 32790 23962
rect 32802 23910 32854 23962
rect 32866 23910 32918 23962
rect 37610 23910 37662 23962
rect 37674 23910 37726 23962
rect 37738 23910 37790 23962
rect 37802 23910 37854 23962
rect 37866 23910 37918 23962
rect 9680 23740 9732 23792
rect 33232 23740 33284 23792
rect 21732 23672 21784 23724
rect 2320 23536 2372 23588
rect 21824 23468 21876 23520
rect 33416 23511 33468 23520
rect 33416 23477 33425 23511
rect 33425 23477 33459 23511
rect 33459 23477 33468 23511
rect 33416 23468 33468 23477
rect 1950 23366 2002 23418
rect 2014 23366 2066 23418
rect 2078 23366 2130 23418
rect 2142 23366 2194 23418
rect 2206 23366 2258 23418
rect 6950 23366 7002 23418
rect 7014 23366 7066 23418
rect 7078 23366 7130 23418
rect 7142 23366 7194 23418
rect 7206 23366 7258 23418
rect 11950 23366 12002 23418
rect 12014 23366 12066 23418
rect 12078 23366 12130 23418
rect 12142 23366 12194 23418
rect 12206 23366 12258 23418
rect 16950 23366 17002 23418
rect 17014 23366 17066 23418
rect 17078 23366 17130 23418
rect 17142 23366 17194 23418
rect 17206 23366 17258 23418
rect 21950 23366 22002 23418
rect 22014 23366 22066 23418
rect 22078 23366 22130 23418
rect 22142 23366 22194 23418
rect 22206 23366 22258 23418
rect 26950 23366 27002 23418
rect 27014 23366 27066 23418
rect 27078 23366 27130 23418
rect 27142 23366 27194 23418
rect 27206 23366 27258 23418
rect 31950 23366 32002 23418
rect 32014 23366 32066 23418
rect 32078 23366 32130 23418
rect 32142 23366 32194 23418
rect 32206 23366 32258 23418
rect 36950 23366 37002 23418
rect 37014 23366 37066 23418
rect 37078 23366 37130 23418
rect 37142 23366 37194 23418
rect 37206 23366 37258 23418
rect 19616 23196 19668 23248
rect 10324 23060 10376 23112
rect 14188 23060 14240 23112
rect 16488 23103 16540 23112
rect 16488 23069 16497 23103
rect 16497 23069 16531 23103
rect 16531 23069 16540 23103
rect 16488 23060 16540 23069
rect 3240 22992 3292 23044
rect 25044 22992 25096 23044
rect 5632 22924 5684 22976
rect 9864 22924 9916 22976
rect 38660 22924 38712 22976
rect 2610 22822 2662 22874
rect 2674 22822 2726 22874
rect 2738 22822 2790 22874
rect 2802 22822 2854 22874
rect 2866 22822 2918 22874
rect 7610 22822 7662 22874
rect 7674 22822 7726 22874
rect 7738 22822 7790 22874
rect 7802 22822 7854 22874
rect 7866 22822 7918 22874
rect 12610 22822 12662 22874
rect 12674 22822 12726 22874
rect 12738 22822 12790 22874
rect 12802 22822 12854 22874
rect 12866 22822 12918 22874
rect 17610 22822 17662 22874
rect 17674 22822 17726 22874
rect 17738 22822 17790 22874
rect 17802 22822 17854 22874
rect 17866 22822 17918 22874
rect 22610 22822 22662 22874
rect 22674 22822 22726 22874
rect 22738 22822 22790 22874
rect 22802 22822 22854 22874
rect 22866 22822 22918 22874
rect 27610 22822 27662 22874
rect 27674 22822 27726 22874
rect 27738 22822 27790 22874
rect 27802 22822 27854 22874
rect 27866 22822 27918 22874
rect 32610 22822 32662 22874
rect 32674 22822 32726 22874
rect 32738 22822 32790 22874
rect 32802 22822 32854 22874
rect 32866 22822 32918 22874
rect 37610 22822 37662 22874
rect 37674 22822 37726 22874
rect 37738 22822 37790 22874
rect 37802 22822 37854 22874
rect 37866 22822 37918 22874
rect 3240 22763 3292 22772
rect 3240 22729 3249 22763
rect 3249 22729 3283 22763
rect 3283 22729 3292 22763
rect 3240 22720 3292 22729
rect 6828 22720 6880 22772
rect 6920 22720 6972 22772
rect 19340 22720 19392 22772
rect 7288 22652 7340 22704
rect 24584 22695 24636 22704
rect 24584 22661 24593 22695
rect 24593 22661 24627 22695
rect 24627 22661 24636 22695
rect 24584 22652 24636 22661
rect 3240 22627 3292 22636
rect 3240 22593 3249 22627
rect 3249 22593 3283 22627
rect 3283 22593 3292 22627
rect 3240 22584 3292 22593
rect 3516 22627 3568 22636
rect 3516 22593 3525 22627
rect 3525 22593 3559 22627
rect 3559 22593 3568 22627
rect 3516 22584 3568 22593
rect 5632 22516 5684 22568
rect 6184 22448 6236 22500
rect 8300 22584 8352 22636
rect 8668 22516 8720 22568
rect 36176 22448 36228 22500
rect 24676 22380 24728 22432
rect 1950 22278 2002 22330
rect 2014 22278 2066 22330
rect 2078 22278 2130 22330
rect 2142 22278 2194 22330
rect 2206 22278 2258 22330
rect 6950 22278 7002 22330
rect 7014 22278 7066 22330
rect 7078 22278 7130 22330
rect 7142 22278 7194 22330
rect 7206 22278 7258 22330
rect 11950 22278 12002 22330
rect 12014 22278 12066 22330
rect 12078 22278 12130 22330
rect 12142 22278 12194 22330
rect 12206 22278 12258 22330
rect 16950 22278 17002 22330
rect 17014 22278 17066 22330
rect 17078 22278 17130 22330
rect 17142 22278 17194 22330
rect 17206 22278 17258 22330
rect 21950 22278 22002 22330
rect 22014 22278 22066 22330
rect 22078 22278 22130 22330
rect 22142 22278 22194 22330
rect 22206 22278 22258 22330
rect 26950 22278 27002 22330
rect 27014 22278 27066 22330
rect 27078 22278 27130 22330
rect 27142 22278 27194 22330
rect 27206 22278 27258 22330
rect 31950 22278 32002 22330
rect 32014 22278 32066 22330
rect 32078 22278 32130 22330
rect 32142 22278 32194 22330
rect 32206 22278 32258 22330
rect 36950 22278 37002 22330
rect 37014 22278 37066 22330
rect 37078 22278 37130 22330
rect 37142 22278 37194 22330
rect 37206 22278 37258 22330
rect 6920 22176 6972 22228
rect 7288 22176 7340 22228
rect 9588 22176 9640 22228
rect 11612 22176 11664 22228
rect 3516 22040 3568 22092
rect 7288 22040 7340 22092
rect 8392 22040 8444 22092
rect 11060 21947 11112 21956
rect 11060 21913 11069 21947
rect 11069 21913 11103 21947
rect 11103 21913 11112 21947
rect 11060 21904 11112 21913
rect 23388 21904 23440 21956
rect 24676 21947 24728 21956
rect 24676 21913 24685 21947
rect 24685 21913 24719 21947
rect 24719 21913 24728 21947
rect 24676 21904 24728 21913
rect 2610 21734 2662 21786
rect 2674 21734 2726 21786
rect 2738 21734 2790 21786
rect 2802 21734 2854 21786
rect 2866 21734 2918 21786
rect 7610 21734 7662 21786
rect 7674 21734 7726 21786
rect 7738 21734 7790 21786
rect 7802 21734 7854 21786
rect 7866 21734 7918 21786
rect 12610 21734 12662 21786
rect 12674 21734 12726 21786
rect 12738 21734 12790 21786
rect 12802 21734 12854 21786
rect 12866 21734 12918 21786
rect 17610 21734 17662 21786
rect 17674 21734 17726 21786
rect 17738 21734 17790 21786
rect 17802 21734 17854 21786
rect 17866 21734 17918 21786
rect 22610 21734 22662 21786
rect 22674 21734 22726 21786
rect 22738 21734 22790 21786
rect 22802 21734 22854 21786
rect 22866 21734 22918 21786
rect 27610 21734 27662 21786
rect 27674 21734 27726 21786
rect 27738 21734 27790 21786
rect 27802 21734 27854 21786
rect 27866 21734 27918 21786
rect 32610 21734 32662 21786
rect 32674 21734 32726 21786
rect 32738 21734 32790 21786
rect 32802 21734 32854 21786
rect 32866 21734 32918 21786
rect 37610 21734 37662 21786
rect 37674 21734 37726 21786
rect 37738 21734 37790 21786
rect 37802 21734 37854 21786
rect 37866 21734 37918 21786
rect 22376 21564 22428 21616
rect 27528 21564 27580 21616
rect 31116 21564 31168 21616
rect 31668 21564 31720 21616
rect 22560 21539 22612 21548
rect 22560 21505 22569 21539
rect 22569 21505 22603 21539
rect 22603 21505 22612 21539
rect 22560 21496 22612 21505
rect 37372 21496 37424 21548
rect 6920 21292 6972 21344
rect 22560 21292 22612 21344
rect 23388 21292 23440 21344
rect 29000 21428 29052 21480
rect 31760 21360 31812 21412
rect 32404 21292 32456 21344
rect 36636 21428 36688 21480
rect 1950 21190 2002 21242
rect 2014 21190 2066 21242
rect 2078 21190 2130 21242
rect 2142 21190 2194 21242
rect 2206 21190 2258 21242
rect 6950 21190 7002 21242
rect 7014 21190 7066 21242
rect 7078 21190 7130 21242
rect 7142 21190 7194 21242
rect 7206 21190 7258 21242
rect 11950 21190 12002 21242
rect 12014 21190 12066 21242
rect 12078 21190 12130 21242
rect 12142 21190 12194 21242
rect 12206 21190 12258 21242
rect 16950 21190 17002 21242
rect 17014 21190 17066 21242
rect 17078 21190 17130 21242
rect 17142 21190 17194 21242
rect 17206 21190 17258 21242
rect 21950 21190 22002 21242
rect 22014 21190 22066 21242
rect 22078 21190 22130 21242
rect 22142 21190 22194 21242
rect 22206 21190 22258 21242
rect 26950 21190 27002 21242
rect 27014 21190 27066 21242
rect 27078 21190 27130 21242
rect 27142 21190 27194 21242
rect 27206 21190 27258 21242
rect 31950 21190 32002 21242
rect 32014 21190 32066 21242
rect 32078 21190 32130 21242
rect 32142 21190 32194 21242
rect 32206 21190 32258 21242
rect 36950 21190 37002 21242
rect 37014 21190 37066 21242
rect 37078 21190 37130 21242
rect 37142 21190 37194 21242
rect 37206 21190 37258 21242
rect 2610 20646 2662 20698
rect 2674 20646 2726 20698
rect 2738 20646 2790 20698
rect 2802 20646 2854 20698
rect 2866 20646 2918 20698
rect 7610 20646 7662 20698
rect 7674 20646 7726 20698
rect 7738 20646 7790 20698
rect 7802 20646 7854 20698
rect 7866 20646 7918 20698
rect 12610 20646 12662 20698
rect 12674 20646 12726 20698
rect 12738 20646 12790 20698
rect 12802 20646 12854 20698
rect 12866 20646 12918 20698
rect 17610 20646 17662 20698
rect 17674 20646 17726 20698
rect 17738 20646 17790 20698
rect 17802 20646 17854 20698
rect 17866 20646 17918 20698
rect 22610 20646 22662 20698
rect 22674 20646 22726 20698
rect 22738 20646 22790 20698
rect 22802 20646 22854 20698
rect 22866 20646 22918 20698
rect 27610 20646 27662 20698
rect 27674 20646 27726 20698
rect 27738 20646 27790 20698
rect 27802 20646 27854 20698
rect 27866 20646 27918 20698
rect 32610 20646 32662 20698
rect 32674 20646 32726 20698
rect 32738 20646 32790 20698
rect 32802 20646 32854 20698
rect 32866 20646 32918 20698
rect 37610 20646 37662 20698
rect 37674 20646 37726 20698
rect 37738 20646 37790 20698
rect 37802 20646 37854 20698
rect 37866 20646 37918 20698
rect 3424 20476 3476 20528
rect 40408 20476 40460 20528
rect 6644 20340 6696 20392
rect 39580 20204 39632 20256
rect 1950 20102 2002 20154
rect 2014 20102 2066 20154
rect 2078 20102 2130 20154
rect 2142 20102 2194 20154
rect 2206 20102 2258 20154
rect 6950 20102 7002 20154
rect 7014 20102 7066 20154
rect 7078 20102 7130 20154
rect 7142 20102 7194 20154
rect 7206 20102 7258 20154
rect 11950 20102 12002 20154
rect 12014 20102 12066 20154
rect 12078 20102 12130 20154
rect 12142 20102 12194 20154
rect 12206 20102 12258 20154
rect 16950 20102 17002 20154
rect 17014 20102 17066 20154
rect 17078 20102 17130 20154
rect 17142 20102 17194 20154
rect 17206 20102 17258 20154
rect 21950 20102 22002 20154
rect 22014 20102 22066 20154
rect 22078 20102 22130 20154
rect 22142 20102 22194 20154
rect 22206 20102 22258 20154
rect 26950 20102 27002 20154
rect 27014 20102 27066 20154
rect 27078 20102 27130 20154
rect 27142 20102 27194 20154
rect 27206 20102 27258 20154
rect 31950 20102 32002 20154
rect 32014 20102 32066 20154
rect 32078 20102 32130 20154
rect 32142 20102 32194 20154
rect 32206 20102 32258 20154
rect 36950 20102 37002 20154
rect 37014 20102 37066 20154
rect 37078 20102 37130 20154
rect 37142 20102 37194 20154
rect 37206 20102 37258 20154
rect 23020 20000 23072 20052
rect 19432 19864 19484 19916
rect 20996 19907 21048 19916
rect 20996 19873 21005 19907
rect 21005 19873 21039 19907
rect 21039 19873 21048 19907
rect 20996 19864 21048 19873
rect 23388 19864 23440 19916
rect 8208 19796 8260 19848
rect 24400 19796 24452 19848
rect 2610 19558 2662 19610
rect 2674 19558 2726 19610
rect 2738 19558 2790 19610
rect 2802 19558 2854 19610
rect 2866 19558 2918 19610
rect 7610 19558 7662 19610
rect 7674 19558 7726 19610
rect 7738 19558 7790 19610
rect 7802 19558 7854 19610
rect 7866 19558 7918 19610
rect 12610 19558 12662 19610
rect 12674 19558 12726 19610
rect 12738 19558 12790 19610
rect 12802 19558 12854 19610
rect 12866 19558 12918 19610
rect 17610 19558 17662 19610
rect 17674 19558 17726 19610
rect 17738 19558 17790 19610
rect 17802 19558 17854 19610
rect 17866 19558 17918 19610
rect 22610 19558 22662 19610
rect 22674 19558 22726 19610
rect 22738 19558 22790 19610
rect 22802 19558 22854 19610
rect 22866 19558 22918 19610
rect 27610 19558 27662 19610
rect 27674 19558 27726 19610
rect 27738 19558 27790 19610
rect 27802 19558 27854 19610
rect 27866 19558 27918 19610
rect 32610 19558 32662 19610
rect 32674 19558 32726 19610
rect 32738 19558 32790 19610
rect 32802 19558 32854 19610
rect 32866 19558 32918 19610
rect 37610 19558 37662 19610
rect 37674 19558 37726 19610
rect 37738 19558 37790 19610
rect 37802 19558 37854 19610
rect 37866 19558 37918 19610
rect 6644 19456 6696 19508
rect 9588 19456 9640 19508
rect 30840 19388 30892 19440
rect 6644 19363 6696 19372
rect 6644 19329 6653 19363
rect 6653 19329 6687 19363
rect 6687 19329 6696 19363
rect 6644 19320 6696 19329
rect 8668 19363 8720 19372
rect 8668 19329 8677 19363
rect 8677 19329 8711 19363
rect 8711 19329 8720 19363
rect 8668 19320 8720 19329
rect 1860 19252 1912 19304
rect 1950 19014 2002 19066
rect 2014 19014 2066 19066
rect 2078 19014 2130 19066
rect 2142 19014 2194 19066
rect 2206 19014 2258 19066
rect 6950 19014 7002 19066
rect 7014 19014 7066 19066
rect 7078 19014 7130 19066
rect 7142 19014 7194 19066
rect 7206 19014 7258 19066
rect 11950 19014 12002 19066
rect 12014 19014 12066 19066
rect 12078 19014 12130 19066
rect 12142 19014 12194 19066
rect 12206 19014 12258 19066
rect 16950 19014 17002 19066
rect 17014 19014 17066 19066
rect 17078 19014 17130 19066
rect 17142 19014 17194 19066
rect 17206 19014 17258 19066
rect 21950 19014 22002 19066
rect 22014 19014 22066 19066
rect 22078 19014 22130 19066
rect 22142 19014 22194 19066
rect 22206 19014 22258 19066
rect 26950 19014 27002 19066
rect 27014 19014 27066 19066
rect 27078 19014 27130 19066
rect 27142 19014 27194 19066
rect 27206 19014 27258 19066
rect 31950 19014 32002 19066
rect 32014 19014 32066 19066
rect 32078 19014 32130 19066
rect 32142 19014 32194 19066
rect 32206 19014 32258 19066
rect 36950 19014 37002 19066
rect 37014 19014 37066 19066
rect 37078 19014 37130 19066
rect 37142 19014 37194 19066
rect 37206 19014 37258 19066
rect 9588 18819 9640 18828
rect 9588 18785 9597 18819
rect 9597 18785 9631 18819
rect 9631 18785 9640 18819
rect 9588 18776 9640 18785
rect 25964 18776 26016 18828
rect 9864 18683 9916 18692
rect 9864 18649 9873 18683
rect 9873 18649 9907 18683
rect 9907 18649 9916 18683
rect 9864 18640 9916 18649
rect 3608 18615 3660 18624
rect 3608 18581 3617 18615
rect 3617 18581 3651 18615
rect 3651 18581 3660 18615
rect 3608 18572 3660 18581
rect 17316 18640 17368 18692
rect 39856 18640 39908 18692
rect 2610 18470 2662 18522
rect 2674 18470 2726 18522
rect 2738 18470 2790 18522
rect 2802 18470 2854 18522
rect 2866 18470 2918 18522
rect 7610 18470 7662 18522
rect 7674 18470 7726 18522
rect 7738 18470 7790 18522
rect 7802 18470 7854 18522
rect 7866 18470 7918 18522
rect 12610 18470 12662 18522
rect 12674 18470 12726 18522
rect 12738 18470 12790 18522
rect 12802 18470 12854 18522
rect 12866 18470 12918 18522
rect 17610 18470 17662 18522
rect 17674 18470 17726 18522
rect 17738 18470 17790 18522
rect 17802 18470 17854 18522
rect 17866 18470 17918 18522
rect 22610 18470 22662 18522
rect 22674 18470 22726 18522
rect 22738 18470 22790 18522
rect 22802 18470 22854 18522
rect 22866 18470 22918 18522
rect 27610 18470 27662 18522
rect 27674 18470 27726 18522
rect 27738 18470 27790 18522
rect 27802 18470 27854 18522
rect 27866 18470 27918 18522
rect 32610 18470 32662 18522
rect 32674 18470 32726 18522
rect 32738 18470 32790 18522
rect 32802 18470 32854 18522
rect 32866 18470 32918 18522
rect 37610 18470 37662 18522
rect 37674 18470 37726 18522
rect 37738 18470 37790 18522
rect 37802 18470 37854 18522
rect 37866 18470 37918 18522
rect 3608 18368 3660 18420
rect 9864 18368 9916 18420
rect 36636 18411 36688 18420
rect 36636 18377 36645 18411
rect 36645 18377 36679 18411
rect 36679 18377 36688 18411
rect 36636 18368 36688 18377
rect 33416 18300 33468 18352
rect 24124 18164 24176 18216
rect 9220 18096 9272 18148
rect 26792 18096 26844 18148
rect 26976 18096 27028 18148
rect 1676 18028 1728 18080
rect 24124 18028 24176 18080
rect 1950 17926 2002 17978
rect 2014 17926 2066 17978
rect 2078 17926 2130 17978
rect 2142 17926 2194 17978
rect 2206 17926 2258 17978
rect 6950 17926 7002 17978
rect 7014 17926 7066 17978
rect 7078 17926 7130 17978
rect 7142 17926 7194 17978
rect 7206 17926 7258 17978
rect 11950 17926 12002 17978
rect 12014 17926 12066 17978
rect 12078 17926 12130 17978
rect 12142 17926 12194 17978
rect 12206 17926 12258 17978
rect 16950 17926 17002 17978
rect 17014 17926 17066 17978
rect 17078 17926 17130 17978
rect 17142 17926 17194 17978
rect 17206 17926 17258 17978
rect 21950 17926 22002 17978
rect 22014 17926 22066 17978
rect 22078 17926 22130 17978
rect 22142 17926 22194 17978
rect 22206 17926 22258 17978
rect 26950 17926 27002 17978
rect 27014 17926 27066 17978
rect 27078 17926 27130 17978
rect 27142 17926 27194 17978
rect 27206 17926 27258 17978
rect 31950 17926 32002 17978
rect 32014 17926 32066 17978
rect 32078 17926 32130 17978
rect 32142 17926 32194 17978
rect 32206 17926 32258 17978
rect 36950 17926 37002 17978
rect 37014 17926 37066 17978
rect 37078 17926 37130 17978
rect 37142 17926 37194 17978
rect 37206 17926 37258 17978
rect 20812 17824 20864 17876
rect 21180 17824 21232 17876
rect 36452 17824 36504 17876
rect 3884 17620 3936 17672
rect 3332 17552 3384 17604
rect 8668 17552 8720 17604
rect 9128 17552 9180 17604
rect 2964 17484 3016 17536
rect 7472 17484 7524 17536
rect 18512 17552 18564 17604
rect 38200 17552 38252 17604
rect 36544 17484 36596 17536
rect 2610 17382 2662 17434
rect 2674 17382 2726 17434
rect 2738 17382 2790 17434
rect 2802 17382 2854 17434
rect 2866 17382 2918 17434
rect 7610 17382 7662 17434
rect 7674 17382 7726 17434
rect 7738 17382 7790 17434
rect 7802 17382 7854 17434
rect 7866 17382 7918 17434
rect 12610 17382 12662 17434
rect 12674 17382 12726 17434
rect 12738 17382 12790 17434
rect 12802 17382 12854 17434
rect 12866 17382 12918 17434
rect 17610 17382 17662 17434
rect 17674 17382 17726 17434
rect 17738 17382 17790 17434
rect 17802 17382 17854 17434
rect 17866 17382 17918 17434
rect 22610 17382 22662 17434
rect 22674 17382 22726 17434
rect 22738 17382 22790 17434
rect 22802 17382 22854 17434
rect 22866 17382 22918 17434
rect 27610 17382 27662 17434
rect 27674 17382 27726 17434
rect 27738 17382 27790 17434
rect 27802 17382 27854 17434
rect 27866 17382 27918 17434
rect 32610 17382 32662 17434
rect 32674 17382 32726 17434
rect 32738 17382 32790 17434
rect 32802 17382 32854 17434
rect 32866 17382 32918 17434
rect 37610 17382 37662 17434
rect 37674 17382 37726 17434
rect 37738 17382 37790 17434
rect 37802 17382 37854 17434
rect 37866 17382 37918 17434
rect 3332 17323 3384 17332
rect 3332 17289 3341 17323
rect 3341 17289 3375 17323
rect 3375 17289 3384 17323
rect 3332 17280 3384 17289
rect 2964 17212 3016 17264
rect 3884 17212 3936 17264
rect 6460 17212 6512 17264
rect 6184 17144 6236 17196
rect 5724 17076 5776 17128
rect 18420 17280 18472 17332
rect 18604 17280 18656 17332
rect 18788 17323 18840 17332
rect 18788 17289 18797 17323
rect 18797 17289 18831 17323
rect 18831 17289 18840 17323
rect 18788 17280 18840 17289
rect 33968 17280 34020 17332
rect 18512 17255 18564 17264
rect 18512 17221 18521 17255
rect 18521 17221 18555 17255
rect 18555 17221 18564 17255
rect 18512 17212 18564 17221
rect 18880 17255 18932 17264
rect 18880 17221 18889 17255
rect 18889 17221 18923 17255
rect 18923 17221 18932 17255
rect 18880 17212 18932 17221
rect 20444 17212 20496 17264
rect 28724 17255 28776 17264
rect 28724 17221 28733 17255
rect 28733 17221 28767 17255
rect 28767 17221 28776 17255
rect 28724 17212 28776 17221
rect 28908 17255 28960 17264
rect 28908 17221 28917 17255
rect 28917 17221 28951 17255
rect 28951 17221 28960 17255
rect 28908 17212 28960 17221
rect 29000 17212 29052 17264
rect 19524 17187 19576 17196
rect 19524 17153 19533 17187
rect 19533 17153 19567 17187
rect 19567 17153 19576 17187
rect 19524 17144 19576 17153
rect 29092 17144 29144 17196
rect 21732 17076 21784 17128
rect 15660 17008 15712 17060
rect 1676 16940 1728 16992
rect 3884 16983 3936 16992
rect 3884 16949 3893 16983
rect 3893 16949 3927 16983
rect 3927 16949 3936 16983
rect 3884 16940 3936 16949
rect 4528 16983 4580 16992
rect 4528 16949 4537 16983
rect 4537 16949 4571 16983
rect 4571 16949 4580 16983
rect 4528 16940 4580 16949
rect 17316 16940 17368 16992
rect 28540 16983 28592 16992
rect 28540 16949 28549 16983
rect 28549 16949 28583 16983
rect 28583 16949 28592 16983
rect 28540 16940 28592 16949
rect 1950 16838 2002 16890
rect 2014 16838 2066 16890
rect 2078 16838 2130 16890
rect 2142 16838 2194 16890
rect 2206 16838 2258 16890
rect 6950 16838 7002 16890
rect 7014 16838 7066 16890
rect 7078 16838 7130 16890
rect 7142 16838 7194 16890
rect 7206 16838 7258 16890
rect 11950 16838 12002 16890
rect 12014 16838 12066 16890
rect 12078 16838 12130 16890
rect 12142 16838 12194 16890
rect 12206 16838 12258 16890
rect 16950 16838 17002 16890
rect 17014 16838 17066 16890
rect 17078 16838 17130 16890
rect 17142 16838 17194 16890
rect 17206 16838 17258 16890
rect 21950 16838 22002 16890
rect 22014 16838 22066 16890
rect 22078 16838 22130 16890
rect 22142 16838 22194 16890
rect 22206 16838 22258 16890
rect 26950 16838 27002 16890
rect 27014 16838 27066 16890
rect 27078 16838 27130 16890
rect 27142 16838 27194 16890
rect 27206 16838 27258 16890
rect 31950 16838 32002 16890
rect 32014 16838 32066 16890
rect 32078 16838 32130 16890
rect 32142 16838 32194 16890
rect 32206 16838 32258 16890
rect 36950 16838 37002 16890
rect 37014 16838 37066 16890
rect 37078 16838 37130 16890
rect 37142 16838 37194 16890
rect 37206 16838 37258 16890
rect 4528 16736 4580 16788
rect 28540 16736 28592 16788
rect 14280 16643 14332 16652
rect 14280 16609 14289 16643
rect 14289 16609 14323 16643
rect 14323 16609 14332 16643
rect 14280 16600 14332 16609
rect 21180 16600 21232 16652
rect 23388 16600 23440 16652
rect 30840 16643 30892 16652
rect 30840 16609 30849 16643
rect 30849 16609 30883 16643
rect 30883 16609 30892 16643
rect 30840 16600 30892 16609
rect 31116 16643 31168 16652
rect 31116 16609 31125 16643
rect 31125 16609 31159 16643
rect 31159 16609 31168 16643
rect 31116 16600 31168 16609
rect 14740 16575 14792 16584
rect 14740 16541 14749 16575
rect 14749 16541 14783 16575
rect 14783 16541 14792 16575
rect 14740 16532 14792 16541
rect 15016 16575 15068 16584
rect 15016 16541 15025 16575
rect 15025 16541 15059 16575
rect 15059 16541 15068 16575
rect 15016 16532 15068 16541
rect 15476 16532 15528 16584
rect 34980 16532 35032 16584
rect 18696 16464 18748 16516
rect 39764 16396 39816 16448
rect 2610 16294 2662 16346
rect 2674 16294 2726 16346
rect 2738 16294 2790 16346
rect 2802 16294 2854 16346
rect 2866 16294 2918 16346
rect 7610 16294 7662 16346
rect 7674 16294 7726 16346
rect 7738 16294 7790 16346
rect 7802 16294 7854 16346
rect 7866 16294 7918 16346
rect 12610 16294 12662 16346
rect 12674 16294 12726 16346
rect 12738 16294 12790 16346
rect 12802 16294 12854 16346
rect 12866 16294 12918 16346
rect 17610 16294 17662 16346
rect 17674 16294 17726 16346
rect 17738 16294 17790 16346
rect 17802 16294 17854 16346
rect 17866 16294 17918 16346
rect 22610 16294 22662 16346
rect 22674 16294 22726 16346
rect 22738 16294 22790 16346
rect 22802 16294 22854 16346
rect 22866 16294 22918 16346
rect 27610 16294 27662 16346
rect 27674 16294 27726 16346
rect 27738 16294 27790 16346
rect 27802 16294 27854 16346
rect 27866 16294 27918 16346
rect 32610 16294 32662 16346
rect 32674 16294 32726 16346
rect 32738 16294 32790 16346
rect 32802 16294 32854 16346
rect 32866 16294 32918 16346
rect 37610 16294 37662 16346
rect 37674 16294 37726 16346
rect 37738 16294 37790 16346
rect 37802 16294 37854 16346
rect 37866 16294 37918 16346
rect 15016 16192 15068 16244
rect 20904 16192 20956 16244
rect 22744 15852 22796 15904
rect 23296 15852 23348 15904
rect 38200 15852 38252 15904
rect 1950 15750 2002 15802
rect 2014 15750 2066 15802
rect 2078 15750 2130 15802
rect 2142 15750 2194 15802
rect 2206 15750 2258 15802
rect 6950 15750 7002 15802
rect 7014 15750 7066 15802
rect 7078 15750 7130 15802
rect 7142 15750 7194 15802
rect 7206 15750 7258 15802
rect 11950 15750 12002 15802
rect 12014 15750 12066 15802
rect 12078 15750 12130 15802
rect 12142 15750 12194 15802
rect 12206 15750 12258 15802
rect 16950 15750 17002 15802
rect 17014 15750 17066 15802
rect 17078 15750 17130 15802
rect 17142 15750 17194 15802
rect 17206 15750 17258 15802
rect 21950 15750 22002 15802
rect 22014 15750 22066 15802
rect 22078 15750 22130 15802
rect 22142 15750 22194 15802
rect 22206 15750 22258 15802
rect 26950 15750 27002 15802
rect 27014 15750 27066 15802
rect 27078 15750 27130 15802
rect 27142 15750 27194 15802
rect 27206 15750 27258 15802
rect 31950 15750 32002 15802
rect 32014 15750 32066 15802
rect 32078 15750 32130 15802
rect 32142 15750 32194 15802
rect 32206 15750 32258 15802
rect 36950 15750 37002 15802
rect 37014 15750 37066 15802
rect 37078 15750 37130 15802
rect 37142 15750 37194 15802
rect 37206 15750 37258 15802
rect 14096 15487 14148 15496
rect 14096 15453 14105 15487
rect 14105 15453 14139 15487
rect 14139 15453 14148 15487
rect 14096 15444 14148 15453
rect 14372 15487 14424 15496
rect 14372 15453 14381 15487
rect 14381 15453 14415 15487
rect 14415 15453 14424 15487
rect 14372 15444 14424 15453
rect 22744 15376 22796 15428
rect 14188 15351 14240 15360
rect 14188 15317 14197 15351
rect 14197 15317 14231 15351
rect 14231 15317 14240 15351
rect 14188 15308 14240 15317
rect 33232 15308 33284 15360
rect 2610 15206 2662 15258
rect 2674 15206 2726 15258
rect 2738 15206 2790 15258
rect 2802 15206 2854 15258
rect 2866 15206 2918 15258
rect 7610 15206 7662 15258
rect 7674 15206 7726 15258
rect 7738 15206 7790 15258
rect 7802 15206 7854 15258
rect 7866 15206 7918 15258
rect 12610 15206 12662 15258
rect 12674 15206 12726 15258
rect 12738 15206 12790 15258
rect 12802 15206 12854 15258
rect 12866 15206 12918 15258
rect 17610 15206 17662 15258
rect 17674 15206 17726 15258
rect 17738 15206 17790 15258
rect 17802 15206 17854 15258
rect 17866 15206 17918 15258
rect 22610 15206 22662 15258
rect 22674 15206 22726 15258
rect 22738 15206 22790 15258
rect 22802 15206 22854 15258
rect 22866 15206 22918 15258
rect 27610 15206 27662 15258
rect 27674 15206 27726 15258
rect 27738 15206 27790 15258
rect 27802 15206 27854 15258
rect 27866 15206 27918 15258
rect 32610 15206 32662 15258
rect 32674 15206 32726 15258
rect 32738 15206 32790 15258
rect 32802 15206 32854 15258
rect 32866 15206 32918 15258
rect 37610 15206 37662 15258
rect 37674 15206 37726 15258
rect 37738 15206 37790 15258
rect 37802 15206 37854 15258
rect 37866 15206 37918 15258
rect 31208 15036 31260 15088
rect 32404 15036 32456 15088
rect 38016 15011 38068 15020
rect 38016 14977 38025 15011
rect 38025 14977 38059 15011
rect 38059 14977 38068 15011
rect 38016 14968 38068 14977
rect 38200 15011 38252 15020
rect 38200 14977 38209 15011
rect 38209 14977 38243 15011
rect 38243 14977 38252 15011
rect 38200 14968 38252 14977
rect 33324 14832 33376 14884
rect 24768 14764 24820 14816
rect 1950 14662 2002 14714
rect 2014 14662 2066 14714
rect 2078 14662 2130 14714
rect 2142 14662 2194 14714
rect 2206 14662 2258 14714
rect 6950 14662 7002 14714
rect 7014 14662 7066 14714
rect 7078 14662 7130 14714
rect 7142 14662 7194 14714
rect 7206 14662 7258 14714
rect 11950 14662 12002 14714
rect 12014 14662 12066 14714
rect 12078 14662 12130 14714
rect 12142 14662 12194 14714
rect 12206 14662 12258 14714
rect 16950 14662 17002 14714
rect 17014 14662 17066 14714
rect 17078 14662 17130 14714
rect 17142 14662 17194 14714
rect 17206 14662 17258 14714
rect 21950 14662 22002 14714
rect 22014 14662 22066 14714
rect 22078 14662 22130 14714
rect 22142 14662 22194 14714
rect 22206 14662 22258 14714
rect 26950 14662 27002 14714
rect 27014 14662 27066 14714
rect 27078 14662 27130 14714
rect 27142 14662 27194 14714
rect 27206 14662 27258 14714
rect 31950 14662 32002 14714
rect 32014 14662 32066 14714
rect 32078 14662 32130 14714
rect 32142 14662 32194 14714
rect 32206 14662 32258 14714
rect 36950 14662 37002 14714
rect 37014 14662 37066 14714
rect 37078 14662 37130 14714
rect 37142 14662 37194 14714
rect 37206 14662 37258 14714
rect 31024 14356 31076 14408
rect 38936 14399 38988 14408
rect 38936 14365 38945 14399
rect 38945 14365 38979 14399
rect 38979 14365 38988 14399
rect 38936 14356 38988 14365
rect 18604 14288 18656 14340
rect 2610 14118 2662 14170
rect 2674 14118 2726 14170
rect 2738 14118 2790 14170
rect 2802 14118 2854 14170
rect 2866 14118 2918 14170
rect 7610 14118 7662 14170
rect 7674 14118 7726 14170
rect 7738 14118 7790 14170
rect 7802 14118 7854 14170
rect 7866 14118 7918 14170
rect 12610 14118 12662 14170
rect 12674 14118 12726 14170
rect 12738 14118 12790 14170
rect 12802 14118 12854 14170
rect 12866 14118 12918 14170
rect 17610 14118 17662 14170
rect 17674 14118 17726 14170
rect 17738 14118 17790 14170
rect 17802 14118 17854 14170
rect 17866 14118 17918 14170
rect 22610 14118 22662 14170
rect 22674 14118 22726 14170
rect 22738 14118 22790 14170
rect 22802 14118 22854 14170
rect 22866 14118 22918 14170
rect 27610 14118 27662 14170
rect 27674 14118 27726 14170
rect 27738 14118 27790 14170
rect 27802 14118 27854 14170
rect 27866 14118 27918 14170
rect 32610 14118 32662 14170
rect 32674 14118 32726 14170
rect 32738 14118 32790 14170
rect 32802 14118 32854 14170
rect 32866 14118 32918 14170
rect 37610 14118 37662 14170
rect 37674 14118 37726 14170
rect 37738 14118 37790 14170
rect 37802 14118 37854 14170
rect 37866 14118 37918 14170
rect 9772 14016 9824 14068
rect 8024 13948 8076 14000
rect 18604 13948 18656 14000
rect 29736 13880 29788 13932
rect 9588 13812 9640 13864
rect 13636 13676 13688 13728
rect 1950 13574 2002 13626
rect 2014 13574 2066 13626
rect 2078 13574 2130 13626
rect 2142 13574 2194 13626
rect 2206 13574 2258 13626
rect 6950 13574 7002 13626
rect 7014 13574 7066 13626
rect 7078 13574 7130 13626
rect 7142 13574 7194 13626
rect 7206 13574 7258 13626
rect 11950 13574 12002 13626
rect 12014 13574 12066 13626
rect 12078 13574 12130 13626
rect 12142 13574 12194 13626
rect 12206 13574 12258 13626
rect 16950 13574 17002 13626
rect 17014 13574 17066 13626
rect 17078 13574 17130 13626
rect 17142 13574 17194 13626
rect 17206 13574 17258 13626
rect 21950 13574 22002 13626
rect 22014 13574 22066 13626
rect 22078 13574 22130 13626
rect 22142 13574 22194 13626
rect 22206 13574 22258 13626
rect 26950 13574 27002 13626
rect 27014 13574 27066 13626
rect 27078 13574 27130 13626
rect 27142 13574 27194 13626
rect 27206 13574 27258 13626
rect 31950 13574 32002 13626
rect 32014 13574 32066 13626
rect 32078 13574 32130 13626
rect 32142 13574 32194 13626
rect 32206 13574 32258 13626
rect 36950 13574 37002 13626
rect 37014 13574 37066 13626
rect 37078 13574 37130 13626
rect 37142 13574 37194 13626
rect 37206 13574 37258 13626
rect 27528 13472 27580 13524
rect 34888 13336 34940 13388
rect 15844 13268 15896 13320
rect 16488 13268 16540 13320
rect 39672 13336 39724 13388
rect 36452 13200 36504 13252
rect 2610 13030 2662 13082
rect 2674 13030 2726 13082
rect 2738 13030 2790 13082
rect 2802 13030 2854 13082
rect 2866 13030 2918 13082
rect 7610 13030 7662 13082
rect 7674 13030 7726 13082
rect 7738 13030 7790 13082
rect 7802 13030 7854 13082
rect 7866 13030 7918 13082
rect 12610 13030 12662 13082
rect 12674 13030 12726 13082
rect 12738 13030 12790 13082
rect 12802 13030 12854 13082
rect 12866 13030 12918 13082
rect 17610 13030 17662 13082
rect 17674 13030 17726 13082
rect 17738 13030 17790 13082
rect 17802 13030 17854 13082
rect 17866 13030 17918 13082
rect 22610 13030 22662 13082
rect 22674 13030 22726 13082
rect 22738 13030 22790 13082
rect 22802 13030 22854 13082
rect 22866 13030 22918 13082
rect 27610 13030 27662 13082
rect 27674 13030 27726 13082
rect 27738 13030 27790 13082
rect 27802 13030 27854 13082
rect 27866 13030 27918 13082
rect 32610 13030 32662 13082
rect 32674 13030 32726 13082
rect 32738 13030 32790 13082
rect 32802 13030 32854 13082
rect 32866 13030 32918 13082
rect 37610 13030 37662 13082
rect 37674 13030 37726 13082
rect 37738 13030 37790 13082
rect 37802 13030 37854 13082
rect 37866 13030 37918 13082
rect 1950 12486 2002 12538
rect 2014 12486 2066 12538
rect 2078 12486 2130 12538
rect 2142 12486 2194 12538
rect 2206 12486 2258 12538
rect 6950 12486 7002 12538
rect 7014 12486 7066 12538
rect 7078 12486 7130 12538
rect 7142 12486 7194 12538
rect 7206 12486 7258 12538
rect 11950 12486 12002 12538
rect 12014 12486 12066 12538
rect 12078 12486 12130 12538
rect 12142 12486 12194 12538
rect 12206 12486 12258 12538
rect 16950 12486 17002 12538
rect 17014 12486 17066 12538
rect 17078 12486 17130 12538
rect 17142 12486 17194 12538
rect 17206 12486 17258 12538
rect 21950 12486 22002 12538
rect 22014 12486 22066 12538
rect 22078 12486 22130 12538
rect 22142 12486 22194 12538
rect 22206 12486 22258 12538
rect 26950 12486 27002 12538
rect 27014 12486 27066 12538
rect 27078 12486 27130 12538
rect 27142 12486 27194 12538
rect 27206 12486 27258 12538
rect 31950 12486 32002 12538
rect 32014 12486 32066 12538
rect 32078 12486 32130 12538
rect 32142 12486 32194 12538
rect 32206 12486 32258 12538
rect 36950 12486 37002 12538
rect 37014 12486 37066 12538
rect 37078 12486 37130 12538
rect 37142 12486 37194 12538
rect 37206 12486 37258 12538
rect 18052 12180 18104 12232
rect 18604 12180 18656 12232
rect 18788 12180 18840 12232
rect 4712 12087 4764 12096
rect 4712 12053 4721 12087
rect 4721 12053 4755 12087
rect 4755 12053 4764 12087
rect 4712 12044 4764 12053
rect 23756 12223 23808 12232
rect 23756 12189 23765 12223
rect 23765 12189 23799 12223
rect 23799 12189 23808 12223
rect 23756 12180 23808 12189
rect 38476 12112 38528 12164
rect 25780 12044 25832 12096
rect 2610 11942 2662 11994
rect 2674 11942 2726 11994
rect 2738 11942 2790 11994
rect 2802 11942 2854 11994
rect 2866 11942 2918 11994
rect 7610 11942 7662 11994
rect 7674 11942 7726 11994
rect 7738 11942 7790 11994
rect 7802 11942 7854 11994
rect 7866 11942 7918 11994
rect 12610 11942 12662 11994
rect 12674 11942 12726 11994
rect 12738 11942 12790 11994
rect 12802 11942 12854 11994
rect 12866 11942 12918 11994
rect 17610 11942 17662 11994
rect 17674 11942 17726 11994
rect 17738 11942 17790 11994
rect 17802 11942 17854 11994
rect 17866 11942 17918 11994
rect 22610 11942 22662 11994
rect 22674 11942 22726 11994
rect 22738 11942 22790 11994
rect 22802 11942 22854 11994
rect 22866 11942 22918 11994
rect 27610 11942 27662 11994
rect 27674 11942 27726 11994
rect 27738 11942 27790 11994
rect 27802 11942 27854 11994
rect 27866 11942 27918 11994
rect 32610 11942 32662 11994
rect 32674 11942 32726 11994
rect 32738 11942 32790 11994
rect 32802 11942 32854 11994
rect 32866 11942 32918 11994
rect 37610 11942 37662 11994
rect 37674 11942 37726 11994
rect 37738 11942 37790 11994
rect 37802 11942 37854 11994
rect 37866 11942 37918 11994
rect 1950 11398 2002 11450
rect 2014 11398 2066 11450
rect 2078 11398 2130 11450
rect 2142 11398 2194 11450
rect 2206 11398 2258 11450
rect 6950 11398 7002 11450
rect 7014 11398 7066 11450
rect 7078 11398 7130 11450
rect 7142 11398 7194 11450
rect 7206 11398 7258 11450
rect 11950 11398 12002 11450
rect 12014 11398 12066 11450
rect 12078 11398 12130 11450
rect 12142 11398 12194 11450
rect 12206 11398 12258 11450
rect 16950 11398 17002 11450
rect 17014 11398 17066 11450
rect 17078 11398 17130 11450
rect 17142 11398 17194 11450
rect 17206 11398 17258 11450
rect 21950 11398 22002 11450
rect 22014 11398 22066 11450
rect 22078 11398 22130 11450
rect 22142 11398 22194 11450
rect 22206 11398 22258 11450
rect 26950 11398 27002 11450
rect 27014 11398 27066 11450
rect 27078 11398 27130 11450
rect 27142 11398 27194 11450
rect 27206 11398 27258 11450
rect 31950 11398 32002 11450
rect 32014 11398 32066 11450
rect 32078 11398 32130 11450
rect 32142 11398 32194 11450
rect 32206 11398 32258 11450
rect 36950 11398 37002 11450
rect 37014 11398 37066 11450
rect 37078 11398 37130 11450
rect 37142 11398 37194 11450
rect 37206 11398 37258 11450
rect 29644 11228 29696 11280
rect 30840 11160 30892 11212
rect 33048 11160 33100 11212
rect 6552 11024 6604 11076
rect 2610 10854 2662 10906
rect 2674 10854 2726 10906
rect 2738 10854 2790 10906
rect 2802 10854 2854 10906
rect 2866 10854 2918 10906
rect 7610 10854 7662 10906
rect 7674 10854 7726 10906
rect 7738 10854 7790 10906
rect 7802 10854 7854 10906
rect 7866 10854 7918 10906
rect 12610 10854 12662 10906
rect 12674 10854 12726 10906
rect 12738 10854 12790 10906
rect 12802 10854 12854 10906
rect 12866 10854 12918 10906
rect 17610 10854 17662 10906
rect 17674 10854 17726 10906
rect 17738 10854 17790 10906
rect 17802 10854 17854 10906
rect 17866 10854 17918 10906
rect 22610 10854 22662 10906
rect 22674 10854 22726 10906
rect 22738 10854 22790 10906
rect 22802 10854 22854 10906
rect 22866 10854 22918 10906
rect 27610 10854 27662 10906
rect 27674 10854 27726 10906
rect 27738 10854 27790 10906
rect 27802 10854 27854 10906
rect 27866 10854 27918 10906
rect 32610 10854 32662 10906
rect 32674 10854 32726 10906
rect 32738 10854 32790 10906
rect 32802 10854 32854 10906
rect 32866 10854 32918 10906
rect 37610 10854 37662 10906
rect 37674 10854 37726 10906
rect 37738 10854 37790 10906
rect 37802 10854 37854 10906
rect 37866 10854 37918 10906
rect 33784 10752 33836 10804
rect 36360 10684 36412 10736
rect 33140 10616 33192 10668
rect 36452 10616 36504 10668
rect 3148 10548 3200 10600
rect 22376 10480 22428 10532
rect 38384 10480 38436 10532
rect 1950 10310 2002 10362
rect 2014 10310 2066 10362
rect 2078 10310 2130 10362
rect 2142 10310 2194 10362
rect 2206 10310 2258 10362
rect 6950 10310 7002 10362
rect 7014 10310 7066 10362
rect 7078 10310 7130 10362
rect 7142 10310 7194 10362
rect 7206 10310 7258 10362
rect 11950 10310 12002 10362
rect 12014 10310 12066 10362
rect 12078 10310 12130 10362
rect 12142 10310 12194 10362
rect 12206 10310 12258 10362
rect 16950 10310 17002 10362
rect 17014 10310 17066 10362
rect 17078 10310 17130 10362
rect 17142 10310 17194 10362
rect 17206 10310 17258 10362
rect 21950 10310 22002 10362
rect 22014 10310 22066 10362
rect 22078 10310 22130 10362
rect 22142 10310 22194 10362
rect 22206 10310 22258 10362
rect 26950 10310 27002 10362
rect 27014 10310 27066 10362
rect 27078 10310 27130 10362
rect 27142 10310 27194 10362
rect 27206 10310 27258 10362
rect 31950 10310 32002 10362
rect 32014 10310 32066 10362
rect 32078 10310 32130 10362
rect 32142 10310 32194 10362
rect 32206 10310 32258 10362
rect 36950 10310 37002 10362
rect 37014 10310 37066 10362
rect 37078 10310 37130 10362
rect 37142 10310 37194 10362
rect 37206 10310 37258 10362
rect 2610 9766 2662 9818
rect 2674 9766 2726 9818
rect 2738 9766 2790 9818
rect 2802 9766 2854 9818
rect 2866 9766 2918 9818
rect 7610 9766 7662 9818
rect 7674 9766 7726 9818
rect 7738 9766 7790 9818
rect 7802 9766 7854 9818
rect 7866 9766 7918 9818
rect 12610 9766 12662 9818
rect 12674 9766 12726 9818
rect 12738 9766 12790 9818
rect 12802 9766 12854 9818
rect 12866 9766 12918 9818
rect 17610 9766 17662 9818
rect 17674 9766 17726 9818
rect 17738 9766 17790 9818
rect 17802 9766 17854 9818
rect 17866 9766 17918 9818
rect 22610 9766 22662 9818
rect 22674 9766 22726 9818
rect 22738 9766 22790 9818
rect 22802 9766 22854 9818
rect 22866 9766 22918 9818
rect 27610 9766 27662 9818
rect 27674 9766 27726 9818
rect 27738 9766 27790 9818
rect 27802 9766 27854 9818
rect 27866 9766 27918 9818
rect 32610 9766 32662 9818
rect 32674 9766 32726 9818
rect 32738 9766 32790 9818
rect 32802 9766 32854 9818
rect 32866 9766 32918 9818
rect 37610 9766 37662 9818
rect 37674 9766 37726 9818
rect 37738 9766 37790 9818
rect 37802 9766 37854 9818
rect 37866 9766 37918 9818
rect 7564 9639 7616 9648
rect 7564 9605 7573 9639
rect 7573 9605 7607 9639
rect 7607 9605 7616 9639
rect 7564 9596 7616 9605
rect 17316 9596 17368 9648
rect 19524 9596 19576 9648
rect 19984 9596 20036 9648
rect 10416 9528 10468 9580
rect 13728 9528 13780 9580
rect 9588 9324 9640 9376
rect 38844 9324 38896 9376
rect 1950 9222 2002 9274
rect 2014 9222 2066 9274
rect 2078 9222 2130 9274
rect 2142 9222 2194 9274
rect 2206 9222 2258 9274
rect 6950 9222 7002 9274
rect 7014 9222 7066 9274
rect 7078 9222 7130 9274
rect 7142 9222 7194 9274
rect 7206 9222 7258 9274
rect 11950 9222 12002 9274
rect 12014 9222 12066 9274
rect 12078 9222 12130 9274
rect 12142 9222 12194 9274
rect 12206 9222 12258 9274
rect 16950 9222 17002 9274
rect 17014 9222 17066 9274
rect 17078 9222 17130 9274
rect 17142 9222 17194 9274
rect 17206 9222 17258 9274
rect 21950 9222 22002 9274
rect 22014 9222 22066 9274
rect 22078 9222 22130 9274
rect 22142 9222 22194 9274
rect 22206 9222 22258 9274
rect 26950 9222 27002 9274
rect 27014 9222 27066 9274
rect 27078 9222 27130 9274
rect 27142 9222 27194 9274
rect 27206 9222 27258 9274
rect 31950 9222 32002 9274
rect 32014 9222 32066 9274
rect 32078 9222 32130 9274
rect 32142 9222 32194 9274
rect 32206 9222 32258 9274
rect 36950 9222 37002 9274
rect 37014 9222 37066 9274
rect 37078 9222 37130 9274
rect 37142 9222 37194 9274
rect 37206 9222 37258 9274
rect 7564 9120 7616 9172
rect 22468 9120 22520 9172
rect 33232 9120 33284 9172
rect 9312 8916 9364 8968
rect 14096 8780 14148 8832
rect 38016 8916 38068 8968
rect 38200 8848 38252 8900
rect 2610 8678 2662 8730
rect 2674 8678 2726 8730
rect 2738 8678 2790 8730
rect 2802 8678 2854 8730
rect 2866 8678 2918 8730
rect 7610 8678 7662 8730
rect 7674 8678 7726 8730
rect 7738 8678 7790 8730
rect 7802 8678 7854 8730
rect 7866 8678 7918 8730
rect 12610 8678 12662 8730
rect 12674 8678 12726 8730
rect 12738 8678 12790 8730
rect 12802 8678 12854 8730
rect 12866 8678 12918 8730
rect 17610 8678 17662 8730
rect 17674 8678 17726 8730
rect 17738 8678 17790 8730
rect 17802 8678 17854 8730
rect 17866 8678 17918 8730
rect 22610 8678 22662 8730
rect 22674 8678 22726 8730
rect 22738 8678 22790 8730
rect 22802 8678 22854 8730
rect 22866 8678 22918 8730
rect 27610 8678 27662 8730
rect 27674 8678 27726 8730
rect 27738 8678 27790 8730
rect 27802 8678 27854 8730
rect 27866 8678 27918 8730
rect 32610 8678 32662 8730
rect 32674 8678 32726 8730
rect 32738 8678 32790 8730
rect 32802 8678 32854 8730
rect 32866 8678 32918 8730
rect 37610 8678 37662 8730
rect 37674 8678 37726 8730
rect 37738 8678 37790 8730
rect 37802 8678 37854 8730
rect 37866 8678 37918 8730
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 6950 8134 7002 8186
rect 7014 8134 7066 8186
rect 7078 8134 7130 8186
rect 7142 8134 7194 8186
rect 7206 8134 7258 8186
rect 11950 8134 12002 8186
rect 12014 8134 12066 8186
rect 12078 8134 12130 8186
rect 12142 8134 12194 8186
rect 12206 8134 12258 8186
rect 16950 8134 17002 8186
rect 17014 8134 17066 8186
rect 17078 8134 17130 8186
rect 17142 8134 17194 8186
rect 17206 8134 17258 8186
rect 21950 8134 22002 8186
rect 22014 8134 22066 8186
rect 22078 8134 22130 8186
rect 22142 8134 22194 8186
rect 22206 8134 22258 8186
rect 26950 8134 27002 8186
rect 27014 8134 27066 8186
rect 27078 8134 27130 8186
rect 27142 8134 27194 8186
rect 27206 8134 27258 8186
rect 31950 8134 32002 8186
rect 32014 8134 32066 8186
rect 32078 8134 32130 8186
rect 32142 8134 32194 8186
rect 32206 8134 32258 8186
rect 36950 8134 37002 8186
rect 37014 8134 37066 8186
rect 37078 8134 37130 8186
rect 37142 8134 37194 8186
rect 37206 8134 37258 8186
rect 9496 8032 9548 8084
rect 13636 8032 13688 8084
rect 13728 7828 13780 7880
rect 18880 7871 18932 7880
rect 18880 7837 18889 7871
rect 18889 7837 18923 7871
rect 18923 7837 18932 7871
rect 18880 7828 18932 7837
rect 2610 7590 2662 7642
rect 2674 7590 2726 7642
rect 2738 7590 2790 7642
rect 2802 7590 2854 7642
rect 2866 7590 2918 7642
rect 7610 7590 7662 7642
rect 7674 7590 7726 7642
rect 7738 7590 7790 7642
rect 7802 7590 7854 7642
rect 7866 7590 7918 7642
rect 12610 7590 12662 7642
rect 12674 7590 12726 7642
rect 12738 7590 12790 7642
rect 12802 7590 12854 7642
rect 12866 7590 12918 7642
rect 17610 7590 17662 7642
rect 17674 7590 17726 7642
rect 17738 7590 17790 7642
rect 17802 7590 17854 7642
rect 17866 7590 17918 7642
rect 22610 7590 22662 7642
rect 22674 7590 22726 7642
rect 22738 7590 22790 7642
rect 22802 7590 22854 7642
rect 22866 7590 22918 7642
rect 27610 7590 27662 7642
rect 27674 7590 27726 7642
rect 27738 7590 27790 7642
rect 27802 7590 27854 7642
rect 27866 7590 27918 7642
rect 32610 7590 32662 7642
rect 32674 7590 32726 7642
rect 32738 7590 32790 7642
rect 32802 7590 32854 7642
rect 32866 7590 32918 7642
rect 37610 7590 37662 7642
rect 37674 7590 37726 7642
rect 37738 7590 37790 7642
rect 37802 7590 37854 7642
rect 37866 7590 37918 7642
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 6950 7046 7002 7098
rect 7014 7046 7066 7098
rect 7078 7046 7130 7098
rect 7142 7046 7194 7098
rect 7206 7046 7258 7098
rect 11950 7046 12002 7098
rect 12014 7046 12066 7098
rect 12078 7046 12130 7098
rect 12142 7046 12194 7098
rect 12206 7046 12258 7098
rect 16950 7046 17002 7098
rect 17014 7046 17066 7098
rect 17078 7046 17130 7098
rect 17142 7046 17194 7098
rect 17206 7046 17258 7098
rect 21950 7046 22002 7098
rect 22014 7046 22066 7098
rect 22078 7046 22130 7098
rect 22142 7046 22194 7098
rect 22206 7046 22258 7098
rect 26950 7046 27002 7098
rect 27014 7046 27066 7098
rect 27078 7046 27130 7098
rect 27142 7046 27194 7098
rect 27206 7046 27258 7098
rect 31950 7046 32002 7098
rect 32014 7046 32066 7098
rect 32078 7046 32130 7098
rect 32142 7046 32194 7098
rect 32206 7046 32258 7098
rect 36950 7046 37002 7098
rect 37014 7046 37066 7098
rect 37078 7046 37130 7098
rect 37142 7046 37194 7098
rect 37206 7046 37258 7098
rect 2610 6502 2662 6554
rect 2674 6502 2726 6554
rect 2738 6502 2790 6554
rect 2802 6502 2854 6554
rect 2866 6502 2918 6554
rect 7610 6502 7662 6554
rect 7674 6502 7726 6554
rect 7738 6502 7790 6554
rect 7802 6502 7854 6554
rect 7866 6502 7918 6554
rect 12610 6502 12662 6554
rect 12674 6502 12726 6554
rect 12738 6502 12790 6554
rect 12802 6502 12854 6554
rect 12866 6502 12918 6554
rect 17610 6502 17662 6554
rect 17674 6502 17726 6554
rect 17738 6502 17790 6554
rect 17802 6502 17854 6554
rect 17866 6502 17918 6554
rect 22610 6502 22662 6554
rect 22674 6502 22726 6554
rect 22738 6502 22790 6554
rect 22802 6502 22854 6554
rect 22866 6502 22918 6554
rect 27610 6502 27662 6554
rect 27674 6502 27726 6554
rect 27738 6502 27790 6554
rect 27802 6502 27854 6554
rect 27866 6502 27918 6554
rect 32610 6502 32662 6554
rect 32674 6502 32726 6554
rect 32738 6502 32790 6554
rect 32802 6502 32854 6554
rect 32866 6502 32918 6554
rect 37610 6502 37662 6554
rect 37674 6502 37726 6554
rect 37738 6502 37790 6554
rect 37802 6502 37854 6554
rect 37866 6502 37918 6554
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 6950 5958 7002 6010
rect 7014 5958 7066 6010
rect 7078 5958 7130 6010
rect 7142 5958 7194 6010
rect 7206 5958 7258 6010
rect 11950 5958 12002 6010
rect 12014 5958 12066 6010
rect 12078 5958 12130 6010
rect 12142 5958 12194 6010
rect 12206 5958 12258 6010
rect 16950 5958 17002 6010
rect 17014 5958 17066 6010
rect 17078 5958 17130 6010
rect 17142 5958 17194 6010
rect 17206 5958 17258 6010
rect 21950 5958 22002 6010
rect 22014 5958 22066 6010
rect 22078 5958 22130 6010
rect 22142 5958 22194 6010
rect 22206 5958 22258 6010
rect 26950 5958 27002 6010
rect 27014 5958 27066 6010
rect 27078 5958 27130 6010
rect 27142 5958 27194 6010
rect 27206 5958 27258 6010
rect 31950 5958 32002 6010
rect 32014 5958 32066 6010
rect 32078 5958 32130 6010
rect 32142 5958 32194 6010
rect 32206 5958 32258 6010
rect 36950 5958 37002 6010
rect 37014 5958 37066 6010
rect 37078 5958 37130 6010
rect 37142 5958 37194 6010
rect 37206 5958 37258 6010
rect 2610 5414 2662 5466
rect 2674 5414 2726 5466
rect 2738 5414 2790 5466
rect 2802 5414 2854 5466
rect 2866 5414 2918 5466
rect 7610 5414 7662 5466
rect 7674 5414 7726 5466
rect 7738 5414 7790 5466
rect 7802 5414 7854 5466
rect 7866 5414 7918 5466
rect 12610 5414 12662 5466
rect 12674 5414 12726 5466
rect 12738 5414 12790 5466
rect 12802 5414 12854 5466
rect 12866 5414 12918 5466
rect 17610 5414 17662 5466
rect 17674 5414 17726 5466
rect 17738 5414 17790 5466
rect 17802 5414 17854 5466
rect 17866 5414 17918 5466
rect 22610 5414 22662 5466
rect 22674 5414 22726 5466
rect 22738 5414 22790 5466
rect 22802 5414 22854 5466
rect 22866 5414 22918 5466
rect 27610 5414 27662 5466
rect 27674 5414 27726 5466
rect 27738 5414 27790 5466
rect 27802 5414 27854 5466
rect 27866 5414 27918 5466
rect 32610 5414 32662 5466
rect 32674 5414 32726 5466
rect 32738 5414 32790 5466
rect 32802 5414 32854 5466
rect 32866 5414 32918 5466
rect 37610 5414 37662 5466
rect 37674 5414 37726 5466
rect 37738 5414 37790 5466
rect 37802 5414 37854 5466
rect 37866 5414 37918 5466
rect 19984 5176 20036 5228
rect 6092 4972 6144 5024
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 6950 4870 7002 4922
rect 7014 4870 7066 4922
rect 7078 4870 7130 4922
rect 7142 4870 7194 4922
rect 7206 4870 7258 4922
rect 11950 4870 12002 4922
rect 12014 4870 12066 4922
rect 12078 4870 12130 4922
rect 12142 4870 12194 4922
rect 12206 4870 12258 4922
rect 16950 4870 17002 4922
rect 17014 4870 17066 4922
rect 17078 4870 17130 4922
rect 17142 4870 17194 4922
rect 17206 4870 17258 4922
rect 21950 4870 22002 4922
rect 22014 4870 22066 4922
rect 22078 4870 22130 4922
rect 22142 4870 22194 4922
rect 22206 4870 22258 4922
rect 26950 4870 27002 4922
rect 27014 4870 27066 4922
rect 27078 4870 27130 4922
rect 27142 4870 27194 4922
rect 27206 4870 27258 4922
rect 31950 4870 32002 4922
rect 32014 4870 32066 4922
rect 32078 4870 32130 4922
rect 32142 4870 32194 4922
rect 32206 4870 32258 4922
rect 36950 4870 37002 4922
rect 37014 4870 37066 4922
rect 37078 4870 37130 4922
rect 37142 4870 37194 4922
rect 37206 4870 37258 4922
rect 26056 4811 26108 4820
rect 26056 4777 26065 4811
rect 26065 4777 26099 4811
rect 26099 4777 26108 4811
rect 26056 4768 26108 4777
rect 28908 4700 28960 4752
rect 15844 4632 15896 4684
rect 6276 4607 6328 4616
rect 6276 4573 6285 4607
rect 6285 4573 6319 4607
rect 6319 4573 6328 4607
rect 6276 4564 6328 4573
rect 25780 4607 25832 4616
rect 25780 4573 25789 4607
rect 25789 4573 25823 4607
rect 25823 4573 25832 4607
rect 25780 4564 25832 4573
rect 6184 4471 6236 4480
rect 6184 4437 6193 4471
rect 6193 4437 6227 4471
rect 6227 4437 6236 4471
rect 6184 4428 6236 4437
rect 23756 4496 23808 4548
rect 38752 4428 38804 4480
rect 2610 4326 2662 4378
rect 2674 4326 2726 4378
rect 2738 4326 2790 4378
rect 2802 4326 2854 4378
rect 2866 4326 2918 4378
rect 7610 4326 7662 4378
rect 7674 4326 7726 4378
rect 7738 4326 7790 4378
rect 7802 4326 7854 4378
rect 7866 4326 7918 4378
rect 12610 4326 12662 4378
rect 12674 4326 12726 4378
rect 12738 4326 12790 4378
rect 12802 4326 12854 4378
rect 12866 4326 12918 4378
rect 17610 4326 17662 4378
rect 17674 4326 17726 4378
rect 17738 4326 17790 4378
rect 17802 4326 17854 4378
rect 17866 4326 17918 4378
rect 22610 4326 22662 4378
rect 22674 4326 22726 4378
rect 22738 4326 22790 4378
rect 22802 4326 22854 4378
rect 22866 4326 22918 4378
rect 27610 4326 27662 4378
rect 27674 4326 27726 4378
rect 27738 4326 27790 4378
rect 27802 4326 27854 4378
rect 27866 4326 27918 4378
rect 32610 4326 32662 4378
rect 32674 4326 32726 4378
rect 32738 4326 32790 4378
rect 32802 4326 32854 4378
rect 32866 4326 32918 4378
rect 37610 4326 37662 4378
rect 37674 4326 37726 4378
rect 37738 4326 37790 4378
rect 37802 4326 37854 4378
rect 37866 4326 37918 4378
rect 2504 3952 2556 4004
rect 14280 3952 14332 4004
rect 2872 3884 2924 3936
rect 12348 3884 12400 3936
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 6950 3782 7002 3834
rect 7014 3782 7066 3834
rect 7078 3782 7130 3834
rect 7142 3782 7194 3834
rect 7206 3782 7258 3834
rect 11950 3782 12002 3834
rect 12014 3782 12066 3834
rect 12078 3782 12130 3834
rect 12142 3782 12194 3834
rect 12206 3782 12258 3834
rect 16950 3782 17002 3834
rect 17014 3782 17066 3834
rect 17078 3782 17130 3834
rect 17142 3782 17194 3834
rect 17206 3782 17258 3834
rect 21950 3782 22002 3834
rect 22014 3782 22066 3834
rect 22078 3782 22130 3834
rect 22142 3782 22194 3834
rect 22206 3782 22258 3834
rect 26950 3782 27002 3834
rect 27014 3782 27066 3834
rect 27078 3782 27130 3834
rect 27142 3782 27194 3834
rect 27206 3782 27258 3834
rect 31950 3782 32002 3834
rect 32014 3782 32066 3834
rect 32078 3782 32130 3834
rect 32142 3782 32194 3834
rect 32206 3782 32258 3834
rect 36950 3782 37002 3834
rect 37014 3782 37066 3834
rect 37078 3782 37130 3834
rect 37142 3782 37194 3834
rect 37206 3782 37258 3834
rect 8484 3680 8536 3732
rect 29460 3680 29512 3732
rect 3056 3655 3108 3664
rect 3056 3621 3065 3655
rect 3065 3621 3099 3655
rect 3099 3621 3108 3655
rect 3056 3612 3108 3621
rect 1676 3587 1728 3596
rect 1676 3553 1685 3587
rect 1685 3553 1719 3587
rect 1719 3553 1728 3587
rect 1676 3544 1728 3553
rect 13912 3612 13964 3664
rect 2872 3519 2924 3528
rect 2872 3485 2881 3519
rect 2881 3485 2915 3519
rect 2915 3485 2924 3519
rect 2872 3476 2924 3485
rect 7380 3476 7432 3528
rect 6184 3408 6236 3460
rect 6368 3340 6420 3392
rect 7012 3340 7064 3392
rect 9496 3340 9548 3392
rect 14372 3340 14424 3392
rect 2610 3238 2662 3290
rect 2674 3238 2726 3290
rect 2738 3238 2790 3290
rect 2802 3238 2854 3290
rect 2866 3238 2918 3290
rect 7610 3238 7662 3290
rect 7674 3238 7726 3290
rect 7738 3238 7790 3290
rect 7802 3238 7854 3290
rect 7866 3238 7918 3290
rect 12610 3238 12662 3290
rect 12674 3238 12726 3290
rect 12738 3238 12790 3290
rect 12802 3238 12854 3290
rect 12866 3238 12918 3290
rect 17610 3238 17662 3290
rect 17674 3238 17726 3290
rect 17738 3238 17790 3290
rect 17802 3238 17854 3290
rect 17866 3238 17918 3290
rect 22610 3238 22662 3290
rect 22674 3238 22726 3290
rect 22738 3238 22790 3290
rect 22802 3238 22854 3290
rect 22866 3238 22918 3290
rect 27610 3238 27662 3290
rect 27674 3238 27726 3290
rect 27738 3238 27790 3290
rect 27802 3238 27854 3290
rect 27866 3238 27918 3290
rect 32610 3238 32662 3290
rect 32674 3238 32726 3290
rect 32738 3238 32790 3290
rect 32802 3238 32854 3290
rect 32866 3238 32918 3290
rect 37610 3238 37662 3290
rect 37674 3238 37726 3290
rect 37738 3238 37790 3290
rect 37802 3238 37854 3290
rect 37866 3238 37918 3290
rect 4712 3136 4764 3188
rect 7012 3068 7064 3120
rect 7288 3000 7340 3052
rect 8116 3043 8168 3052
rect 8116 3009 8125 3043
rect 8125 3009 8159 3043
rect 8159 3009 8168 3043
rect 8116 3000 8168 3009
rect 8484 3043 8536 3052
rect 8484 3009 8493 3043
rect 8493 3009 8527 3043
rect 8527 3009 8536 3043
rect 8484 3000 8536 3009
rect 8760 3043 8812 3052
rect 8760 3009 8769 3043
rect 8769 3009 8803 3043
rect 8803 3009 8812 3043
rect 8760 3000 8812 3009
rect 8300 2975 8352 2984
rect 8300 2941 8309 2975
rect 8309 2941 8343 2975
rect 8343 2941 8352 2975
rect 8300 2932 8352 2941
rect 9496 3043 9548 3052
rect 9496 3009 9505 3043
rect 9505 3009 9539 3043
rect 9539 3009 9548 3043
rect 9496 3000 9548 3009
rect 9772 2975 9824 2984
rect 9772 2941 9781 2975
rect 9781 2941 9815 2975
rect 9815 2941 9824 2975
rect 9772 2932 9824 2941
rect 14096 3000 14148 3052
rect 14280 3043 14332 3052
rect 14280 3009 14289 3043
rect 14289 3009 14323 3043
rect 14323 3009 14332 3043
rect 14280 3000 14332 3009
rect 14188 2932 14240 2984
rect 21824 3000 21876 3052
rect 29184 3000 29236 3052
rect 38292 3000 38344 3052
rect 14280 2796 14332 2848
rect 21640 2796 21692 2848
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 6950 2694 7002 2746
rect 7014 2694 7066 2746
rect 7078 2694 7130 2746
rect 7142 2694 7194 2746
rect 7206 2694 7258 2746
rect 11950 2694 12002 2746
rect 12014 2694 12066 2746
rect 12078 2694 12130 2746
rect 12142 2694 12194 2746
rect 12206 2694 12258 2746
rect 16950 2694 17002 2746
rect 17014 2694 17066 2746
rect 17078 2694 17130 2746
rect 17142 2694 17194 2746
rect 17206 2694 17258 2746
rect 21950 2694 22002 2746
rect 22014 2694 22066 2746
rect 22078 2694 22130 2746
rect 22142 2694 22194 2746
rect 22206 2694 22258 2746
rect 26950 2694 27002 2746
rect 27014 2694 27066 2746
rect 27078 2694 27130 2746
rect 27142 2694 27194 2746
rect 27206 2694 27258 2746
rect 31950 2694 32002 2746
rect 32014 2694 32066 2746
rect 32078 2694 32130 2746
rect 32142 2694 32194 2746
rect 32206 2694 32258 2746
rect 36950 2694 37002 2746
rect 37014 2694 37066 2746
rect 37078 2694 37130 2746
rect 37142 2694 37194 2746
rect 37206 2694 37258 2746
rect 36636 2592 36688 2644
rect 15200 2524 15252 2576
rect 18604 2456 18656 2508
rect 30840 2456 30892 2508
rect 2504 2388 2556 2440
rect 9128 2388 9180 2440
rect 31116 2388 31168 2440
rect 39304 2388 39356 2440
rect 10232 2320 10284 2372
rect 8024 2252 8076 2304
rect 13084 2252 13136 2304
rect 18328 2252 18380 2304
rect 23572 2252 23624 2304
rect 28816 2252 28868 2304
rect 34060 2252 34112 2304
rect 2610 2150 2662 2202
rect 2674 2150 2726 2202
rect 2738 2150 2790 2202
rect 2802 2150 2854 2202
rect 2866 2150 2918 2202
rect 7610 2150 7662 2202
rect 7674 2150 7726 2202
rect 7738 2150 7790 2202
rect 7802 2150 7854 2202
rect 7866 2150 7918 2202
rect 12610 2150 12662 2202
rect 12674 2150 12726 2202
rect 12738 2150 12790 2202
rect 12802 2150 12854 2202
rect 12866 2150 12918 2202
rect 17610 2150 17662 2202
rect 17674 2150 17726 2202
rect 17738 2150 17790 2202
rect 17802 2150 17854 2202
rect 17866 2150 17918 2202
rect 22610 2150 22662 2202
rect 22674 2150 22726 2202
rect 22738 2150 22790 2202
rect 22802 2150 22854 2202
rect 22866 2150 22918 2202
rect 27610 2150 27662 2202
rect 27674 2150 27726 2202
rect 27738 2150 27790 2202
rect 27802 2150 27854 2202
rect 27866 2150 27918 2202
rect 32610 2150 32662 2202
rect 32674 2150 32726 2202
rect 32738 2150 32790 2202
rect 32802 2150 32854 2202
rect 32866 2150 32918 2202
rect 37610 2150 37662 2202
rect 37674 2150 37726 2202
rect 37738 2150 37790 2202
rect 37802 2150 37854 2202
rect 37866 2150 37918 2202
<< metal2 >>
rect 2962 71346 3018 72000
rect 2962 71318 3096 71346
rect 2962 71200 3018 71318
rect 2610 69660 2918 69669
rect 2610 69658 2616 69660
rect 2672 69658 2696 69660
rect 2752 69658 2776 69660
rect 2832 69658 2856 69660
rect 2912 69658 2918 69660
rect 2672 69606 2674 69658
rect 2854 69606 2856 69658
rect 2610 69604 2616 69606
rect 2672 69604 2696 69606
rect 2752 69604 2776 69606
rect 2832 69604 2856 69606
rect 2912 69604 2918 69606
rect 2610 69595 2918 69604
rect 3068 69562 3096 71318
rect 8942 71200 8998 72000
rect 14922 71346 14978 72000
rect 20902 71346 20958 72000
rect 26882 71346 26938 72000
rect 32862 71346 32918 72000
rect 38842 71346 38898 72000
rect 14922 71318 15056 71346
rect 14922 71200 14978 71318
rect 7610 69660 7918 69669
rect 7610 69658 7616 69660
rect 7672 69658 7696 69660
rect 7752 69658 7776 69660
rect 7832 69658 7856 69660
rect 7912 69658 7918 69660
rect 7672 69606 7674 69658
rect 7854 69606 7856 69658
rect 7610 69604 7616 69606
rect 7672 69604 7696 69606
rect 7752 69604 7776 69606
rect 7832 69604 7856 69606
rect 7912 69604 7918 69606
rect 7610 69595 7918 69604
rect 8956 69562 8984 71200
rect 12610 69660 12918 69669
rect 12610 69658 12616 69660
rect 12672 69658 12696 69660
rect 12752 69658 12776 69660
rect 12832 69658 12856 69660
rect 12912 69658 12918 69660
rect 12672 69606 12674 69658
rect 12854 69606 12856 69658
rect 12610 69604 12616 69606
rect 12672 69604 12696 69606
rect 12752 69604 12776 69606
rect 12832 69604 12856 69606
rect 12912 69604 12918 69606
rect 12610 69595 12918 69604
rect 15028 69562 15056 71318
rect 20902 71318 21036 71346
rect 20902 71200 20958 71318
rect 17610 69660 17918 69669
rect 17610 69658 17616 69660
rect 17672 69658 17696 69660
rect 17752 69658 17776 69660
rect 17832 69658 17856 69660
rect 17912 69658 17918 69660
rect 17672 69606 17674 69658
rect 17854 69606 17856 69658
rect 17610 69604 17616 69606
rect 17672 69604 17696 69606
rect 17752 69604 17776 69606
rect 17832 69604 17856 69606
rect 17912 69604 17918 69606
rect 17610 69595 17918 69604
rect 21008 69562 21036 71318
rect 26882 71318 27016 71346
rect 26882 71200 26938 71318
rect 22610 69660 22918 69669
rect 22610 69658 22616 69660
rect 22672 69658 22696 69660
rect 22752 69658 22776 69660
rect 22832 69658 22856 69660
rect 22912 69658 22918 69660
rect 22672 69606 22674 69658
rect 22854 69606 22856 69658
rect 22610 69604 22616 69606
rect 22672 69604 22696 69606
rect 22752 69604 22776 69606
rect 22832 69604 22856 69606
rect 22912 69604 22918 69606
rect 22610 69595 22918 69604
rect 26988 69562 27016 71318
rect 32862 71318 32996 71346
rect 32862 71200 32918 71318
rect 27610 69660 27918 69669
rect 27610 69658 27616 69660
rect 27672 69658 27696 69660
rect 27752 69658 27776 69660
rect 27832 69658 27856 69660
rect 27912 69658 27918 69660
rect 27672 69606 27674 69658
rect 27854 69606 27856 69658
rect 27610 69604 27616 69606
rect 27672 69604 27696 69606
rect 27752 69604 27776 69606
rect 27832 69604 27856 69606
rect 27912 69604 27918 69606
rect 27610 69595 27918 69604
rect 32610 69660 32918 69669
rect 32610 69658 32616 69660
rect 32672 69658 32696 69660
rect 32752 69658 32776 69660
rect 32832 69658 32856 69660
rect 32912 69658 32918 69660
rect 32672 69606 32674 69658
rect 32854 69606 32856 69658
rect 32610 69604 32616 69606
rect 32672 69604 32696 69606
rect 32752 69604 32776 69606
rect 32832 69604 32856 69606
rect 32912 69604 32918 69606
rect 32610 69595 32918 69604
rect 32968 69562 32996 71318
rect 38842 71318 38976 71346
rect 38842 71200 38898 71318
rect 37610 69660 37918 69669
rect 37610 69658 37616 69660
rect 37672 69658 37696 69660
rect 37752 69658 37776 69660
rect 37832 69658 37856 69660
rect 37912 69658 37918 69660
rect 37672 69606 37674 69658
rect 37854 69606 37856 69658
rect 37610 69604 37616 69606
rect 37672 69604 37696 69606
rect 37752 69604 37776 69606
rect 37832 69604 37856 69606
rect 37912 69604 37918 69606
rect 37610 69595 37918 69604
rect 38948 69562 38976 71318
rect 3056 69556 3108 69562
rect 3056 69498 3108 69504
rect 8944 69556 8996 69562
rect 8944 69498 8996 69504
rect 15016 69556 15068 69562
rect 15016 69498 15068 69504
rect 20996 69556 21048 69562
rect 20996 69498 21048 69504
rect 26976 69556 27028 69562
rect 26976 69498 27028 69504
rect 32956 69556 33008 69562
rect 32956 69498 33008 69504
rect 38936 69556 38988 69562
rect 38936 69498 38988 69504
rect 3332 69420 3384 69426
rect 3332 69362 3384 69368
rect 9220 69420 9272 69426
rect 9220 69362 9272 69368
rect 15200 69420 15252 69426
rect 15200 69362 15252 69368
rect 21180 69420 21232 69426
rect 21180 69362 21232 69368
rect 27344 69420 27396 69426
rect 27344 69362 27396 69368
rect 33140 69420 33192 69426
rect 33140 69362 33192 69368
rect 39120 69420 39172 69426
rect 39120 69362 39172 69368
rect 1950 69116 2258 69125
rect 1950 69114 1956 69116
rect 2012 69114 2036 69116
rect 2092 69114 2116 69116
rect 2172 69114 2196 69116
rect 2252 69114 2258 69116
rect 2012 69062 2014 69114
rect 2194 69062 2196 69114
rect 1950 69060 1956 69062
rect 2012 69060 2036 69062
rect 2092 69060 2116 69062
rect 2172 69060 2196 69062
rect 2252 69060 2258 69062
rect 1950 69051 2258 69060
rect 2610 68572 2918 68581
rect 2610 68570 2616 68572
rect 2672 68570 2696 68572
rect 2752 68570 2776 68572
rect 2832 68570 2856 68572
rect 2912 68570 2918 68572
rect 2672 68518 2674 68570
rect 2854 68518 2856 68570
rect 2610 68516 2616 68518
rect 2672 68516 2696 68518
rect 2752 68516 2776 68518
rect 2832 68516 2856 68518
rect 2912 68516 2918 68518
rect 2610 68507 2918 68516
rect 1950 68028 2258 68037
rect 1950 68026 1956 68028
rect 2012 68026 2036 68028
rect 2092 68026 2116 68028
rect 2172 68026 2196 68028
rect 2252 68026 2258 68028
rect 2012 67974 2014 68026
rect 2194 67974 2196 68026
rect 1950 67972 1956 67974
rect 2012 67972 2036 67974
rect 2092 67972 2116 67974
rect 2172 67972 2196 67974
rect 2252 67972 2258 67974
rect 1950 67963 2258 67972
rect 2504 67856 2556 67862
rect 2504 67798 2556 67804
rect 2320 67720 2372 67726
rect 2320 67662 2372 67668
rect 1950 66940 2258 66949
rect 1950 66938 1956 66940
rect 2012 66938 2036 66940
rect 2092 66938 2116 66940
rect 2172 66938 2196 66940
rect 2252 66938 2258 66940
rect 2012 66886 2014 66938
rect 2194 66886 2196 66938
rect 1950 66884 1956 66886
rect 2012 66884 2036 66886
rect 2092 66884 2116 66886
rect 2172 66884 2196 66886
rect 2252 66884 2258 66886
rect 1950 66875 2258 66884
rect 1950 65852 2258 65861
rect 1950 65850 1956 65852
rect 2012 65850 2036 65852
rect 2092 65850 2116 65852
rect 2172 65850 2196 65852
rect 2252 65850 2258 65852
rect 2012 65798 2014 65850
rect 2194 65798 2196 65850
rect 1950 65796 1956 65798
rect 2012 65796 2036 65798
rect 2092 65796 2116 65798
rect 2172 65796 2196 65798
rect 2252 65796 2258 65798
rect 1950 65787 2258 65796
rect 1950 64764 2258 64773
rect 1950 64762 1956 64764
rect 2012 64762 2036 64764
rect 2092 64762 2116 64764
rect 2172 64762 2196 64764
rect 2252 64762 2258 64764
rect 2012 64710 2014 64762
rect 2194 64710 2196 64762
rect 1950 64708 1956 64710
rect 2012 64708 2036 64710
rect 2092 64708 2116 64710
rect 2172 64708 2196 64710
rect 2252 64708 2258 64710
rect 1950 64699 2258 64708
rect 1950 63676 2258 63685
rect 1950 63674 1956 63676
rect 2012 63674 2036 63676
rect 2092 63674 2116 63676
rect 2172 63674 2196 63676
rect 2252 63674 2258 63676
rect 2012 63622 2014 63674
rect 2194 63622 2196 63674
rect 1950 63620 1956 63622
rect 2012 63620 2036 63622
rect 2092 63620 2116 63622
rect 2172 63620 2196 63622
rect 2252 63620 2258 63622
rect 1950 63611 2258 63620
rect 1950 62588 2258 62597
rect 1950 62586 1956 62588
rect 2012 62586 2036 62588
rect 2092 62586 2116 62588
rect 2172 62586 2196 62588
rect 2252 62586 2258 62588
rect 2012 62534 2014 62586
rect 2194 62534 2196 62586
rect 1950 62532 1956 62534
rect 2012 62532 2036 62534
rect 2092 62532 2116 62534
rect 2172 62532 2196 62534
rect 2252 62532 2258 62534
rect 1950 62523 2258 62532
rect 1950 61500 2258 61509
rect 1950 61498 1956 61500
rect 2012 61498 2036 61500
rect 2092 61498 2116 61500
rect 2172 61498 2196 61500
rect 2252 61498 2258 61500
rect 2012 61446 2014 61498
rect 2194 61446 2196 61498
rect 1950 61444 1956 61446
rect 2012 61444 2036 61446
rect 2092 61444 2116 61446
rect 2172 61444 2196 61446
rect 2252 61444 2258 61446
rect 1950 61435 2258 61444
rect 1950 60412 2258 60421
rect 1950 60410 1956 60412
rect 2012 60410 2036 60412
rect 2092 60410 2116 60412
rect 2172 60410 2196 60412
rect 2252 60410 2258 60412
rect 2012 60358 2014 60410
rect 2194 60358 2196 60410
rect 1950 60356 1956 60358
rect 2012 60356 2036 60358
rect 2092 60356 2116 60358
rect 2172 60356 2196 60358
rect 2252 60356 2258 60358
rect 1950 60347 2258 60356
rect 1950 59324 2258 59333
rect 1950 59322 1956 59324
rect 2012 59322 2036 59324
rect 2092 59322 2116 59324
rect 2172 59322 2196 59324
rect 2252 59322 2258 59324
rect 2012 59270 2014 59322
rect 2194 59270 2196 59322
rect 1950 59268 1956 59270
rect 2012 59268 2036 59270
rect 2092 59268 2116 59270
rect 2172 59268 2196 59270
rect 2252 59268 2258 59270
rect 1950 59259 2258 59268
rect 1950 58236 2258 58245
rect 1950 58234 1956 58236
rect 2012 58234 2036 58236
rect 2092 58234 2116 58236
rect 2172 58234 2196 58236
rect 2252 58234 2258 58236
rect 2012 58182 2014 58234
rect 2194 58182 2196 58234
rect 1950 58180 1956 58182
rect 2012 58180 2036 58182
rect 2092 58180 2116 58182
rect 2172 58180 2196 58182
rect 2252 58180 2258 58182
rect 1950 58171 2258 58180
rect 1950 57148 2258 57157
rect 1950 57146 1956 57148
rect 2012 57146 2036 57148
rect 2092 57146 2116 57148
rect 2172 57146 2196 57148
rect 2252 57146 2258 57148
rect 2012 57094 2014 57146
rect 2194 57094 2196 57146
rect 1950 57092 1956 57094
rect 2012 57092 2036 57094
rect 2092 57092 2116 57094
rect 2172 57092 2196 57094
rect 2252 57092 2258 57094
rect 1950 57083 2258 57092
rect 1950 56060 2258 56069
rect 1950 56058 1956 56060
rect 2012 56058 2036 56060
rect 2092 56058 2116 56060
rect 2172 56058 2196 56060
rect 2252 56058 2258 56060
rect 2012 56006 2014 56058
rect 2194 56006 2196 56058
rect 1950 56004 1956 56006
rect 2012 56004 2036 56006
rect 2092 56004 2116 56006
rect 2172 56004 2196 56006
rect 2252 56004 2258 56006
rect 1950 55995 2258 56004
rect 1950 54972 2258 54981
rect 1950 54970 1956 54972
rect 2012 54970 2036 54972
rect 2092 54970 2116 54972
rect 2172 54970 2196 54972
rect 2252 54970 2258 54972
rect 2012 54918 2014 54970
rect 2194 54918 2196 54970
rect 1950 54916 1956 54918
rect 2012 54916 2036 54918
rect 2092 54916 2116 54918
rect 2172 54916 2196 54918
rect 2252 54916 2258 54918
rect 1950 54907 2258 54916
rect 1950 53884 2258 53893
rect 1950 53882 1956 53884
rect 2012 53882 2036 53884
rect 2092 53882 2116 53884
rect 2172 53882 2196 53884
rect 2252 53882 2258 53884
rect 2012 53830 2014 53882
rect 2194 53830 2196 53882
rect 1950 53828 1956 53830
rect 2012 53828 2036 53830
rect 2092 53828 2116 53830
rect 2172 53828 2196 53830
rect 2252 53828 2258 53830
rect 1950 53819 2258 53828
rect 1950 52796 2258 52805
rect 1950 52794 1956 52796
rect 2012 52794 2036 52796
rect 2092 52794 2116 52796
rect 2172 52794 2196 52796
rect 2252 52794 2258 52796
rect 2012 52742 2014 52794
rect 2194 52742 2196 52794
rect 1950 52740 1956 52742
rect 2012 52740 2036 52742
rect 2092 52740 2116 52742
rect 2172 52740 2196 52742
rect 2252 52740 2258 52742
rect 1950 52731 2258 52740
rect 1950 51708 2258 51717
rect 1950 51706 1956 51708
rect 2012 51706 2036 51708
rect 2092 51706 2116 51708
rect 2172 51706 2196 51708
rect 2252 51706 2258 51708
rect 2012 51654 2014 51706
rect 2194 51654 2196 51706
rect 1950 51652 1956 51654
rect 2012 51652 2036 51654
rect 2092 51652 2116 51654
rect 2172 51652 2196 51654
rect 2252 51652 2258 51654
rect 1950 51643 2258 51652
rect 1950 50620 2258 50629
rect 1950 50618 1956 50620
rect 2012 50618 2036 50620
rect 2092 50618 2116 50620
rect 2172 50618 2196 50620
rect 2252 50618 2258 50620
rect 2012 50566 2014 50618
rect 2194 50566 2196 50618
rect 1950 50564 1956 50566
rect 2012 50564 2036 50566
rect 2092 50564 2116 50566
rect 2172 50564 2196 50566
rect 2252 50564 2258 50566
rect 1950 50555 2258 50564
rect 1950 49532 2258 49541
rect 1950 49530 1956 49532
rect 2012 49530 2036 49532
rect 2092 49530 2116 49532
rect 2172 49530 2196 49532
rect 2252 49530 2258 49532
rect 2012 49478 2014 49530
rect 2194 49478 2196 49530
rect 1950 49476 1956 49478
rect 2012 49476 2036 49478
rect 2092 49476 2116 49478
rect 2172 49476 2196 49478
rect 2252 49476 2258 49478
rect 1950 49467 2258 49476
rect 1950 48444 2258 48453
rect 1950 48442 1956 48444
rect 2012 48442 2036 48444
rect 2092 48442 2116 48444
rect 2172 48442 2196 48444
rect 2252 48442 2258 48444
rect 2012 48390 2014 48442
rect 2194 48390 2196 48442
rect 1950 48388 1956 48390
rect 2012 48388 2036 48390
rect 2092 48388 2116 48390
rect 2172 48388 2196 48390
rect 2252 48388 2258 48390
rect 1950 48379 2258 48388
rect 1950 47356 2258 47365
rect 1950 47354 1956 47356
rect 2012 47354 2036 47356
rect 2092 47354 2116 47356
rect 2172 47354 2196 47356
rect 2252 47354 2258 47356
rect 2012 47302 2014 47354
rect 2194 47302 2196 47354
rect 1950 47300 1956 47302
rect 2012 47300 2036 47302
rect 2092 47300 2116 47302
rect 2172 47300 2196 47302
rect 2252 47300 2258 47302
rect 1950 47291 2258 47300
rect 1676 47048 1728 47054
rect 1676 46990 1728 46996
rect 1400 45416 1452 45422
rect 1400 45358 1452 45364
rect 1412 45082 1440 45358
rect 1400 45076 1452 45082
rect 1400 45018 1452 45024
rect 1688 18086 1716 46990
rect 1860 46912 1912 46918
rect 1860 46854 1912 46860
rect 1872 19310 1900 46854
rect 1950 46268 2258 46277
rect 1950 46266 1956 46268
rect 2012 46266 2036 46268
rect 2092 46266 2116 46268
rect 2172 46266 2196 46268
rect 2252 46266 2258 46268
rect 2012 46214 2014 46266
rect 2194 46214 2196 46266
rect 1950 46212 1956 46214
rect 2012 46212 2036 46214
rect 2092 46212 2116 46214
rect 2172 46212 2196 46214
rect 2252 46212 2258 46214
rect 1950 46203 2258 46212
rect 1950 45180 2258 45189
rect 1950 45178 1956 45180
rect 2012 45178 2036 45180
rect 2092 45178 2116 45180
rect 2172 45178 2196 45180
rect 2252 45178 2258 45180
rect 2012 45126 2014 45178
rect 2194 45126 2196 45178
rect 1950 45124 1956 45126
rect 2012 45124 2036 45126
rect 2092 45124 2116 45126
rect 2172 45124 2196 45126
rect 2252 45124 2258 45126
rect 1950 45115 2258 45124
rect 1950 44092 2258 44101
rect 1950 44090 1956 44092
rect 2012 44090 2036 44092
rect 2092 44090 2116 44092
rect 2172 44090 2196 44092
rect 2252 44090 2258 44092
rect 2012 44038 2014 44090
rect 2194 44038 2196 44090
rect 1950 44036 1956 44038
rect 2012 44036 2036 44038
rect 2092 44036 2116 44038
rect 2172 44036 2196 44038
rect 2252 44036 2258 44038
rect 1950 44027 2258 44036
rect 1950 43004 2258 43013
rect 1950 43002 1956 43004
rect 2012 43002 2036 43004
rect 2092 43002 2116 43004
rect 2172 43002 2196 43004
rect 2252 43002 2258 43004
rect 2012 42950 2014 43002
rect 2194 42950 2196 43002
rect 1950 42948 1956 42950
rect 2012 42948 2036 42950
rect 2092 42948 2116 42950
rect 2172 42948 2196 42950
rect 2252 42948 2258 42950
rect 1950 42939 2258 42948
rect 1950 41916 2258 41925
rect 1950 41914 1956 41916
rect 2012 41914 2036 41916
rect 2092 41914 2116 41916
rect 2172 41914 2196 41916
rect 2252 41914 2258 41916
rect 2012 41862 2014 41914
rect 2194 41862 2196 41914
rect 1950 41860 1956 41862
rect 2012 41860 2036 41862
rect 2092 41860 2116 41862
rect 2172 41860 2196 41862
rect 2252 41860 2258 41862
rect 1950 41851 2258 41860
rect 1950 40828 2258 40837
rect 1950 40826 1956 40828
rect 2012 40826 2036 40828
rect 2092 40826 2116 40828
rect 2172 40826 2196 40828
rect 2252 40826 2258 40828
rect 2012 40774 2014 40826
rect 2194 40774 2196 40826
rect 1950 40772 1956 40774
rect 2012 40772 2036 40774
rect 2092 40772 2116 40774
rect 2172 40772 2196 40774
rect 2252 40772 2258 40774
rect 1950 40763 2258 40772
rect 1950 39740 2258 39749
rect 1950 39738 1956 39740
rect 2012 39738 2036 39740
rect 2092 39738 2116 39740
rect 2172 39738 2196 39740
rect 2252 39738 2258 39740
rect 2012 39686 2014 39738
rect 2194 39686 2196 39738
rect 1950 39684 1956 39686
rect 2012 39684 2036 39686
rect 2092 39684 2116 39686
rect 2172 39684 2196 39686
rect 2252 39684 2258 39686
rect 1950 39675 2258 39684
rect 1950 38652 2258 38661
rect 1950 38650 1956 38652
rect 2012 38650 2036 38652
rect 2092 38650 2116 38652
rect 2172 38650 2196 38652
rect 2252 38650 2258 38652
rect 2012 38598 2014 38650
rect 2194 38598 2196 38650
rect 1950 38596 1956 38598
rect 2012 38596 2036 38598
rect 2092 38596 2116 38598
rect 2172 38596 2196 38598
rect 2252 38596 2258 38598
rect 1950 38587 2258 38596
rect 1950 37564 2258 37573
rect 1950 37562 1956 37564
rect 2012 37562 2036 37564
rect 2092 37562 2116 37564
rect 2172 37562 2196 37564
rect 2252 37562 2258 37564
rect 2012 37510 2014 37562
rect 2194 37510 2196 37562
rect 1950 37508 1956 37510
rect 2012 37508 2036 37510
rect 2092 37508 2116 37510
rect 2172 37508 2196 37510
rect 2252 37508 2258 37510
rect 1950 37499 2258 37508
rect 1950 36476 2258 36485
rect 1950 36474 1956 36476
rect 2012 36474 2036 36476
rect 2092 36474 2116 36476
rect 2172 36474 2196 36476
rect 2252 36474 2258 36476
rect 2012 36422 2014 36474
rect 2194 36422 2196 36474
rect 1950 36420 1956 36422
rect 2012 36420 2036 36422
rect 2092 36420 2116 36422
rect 2172 36420 2196 36422
rect 2252 36420 2258 36422
rect 1950 36411 2258 36420
rect 1950 35388 2258 35397
rect 1950 35386 1956 35388
rect 2012 35386 2036 35388
rect 2092 35386 2116 35388
rect 2172 35386 2196 35388
rect 2252 35386 2258 35388
rect 2012 35334 2014 35386
rect 2194 35334 2196 35386
rect 1950 35332 1956 35334
rect 2012 35332 2036 35334
rect 2092 35332 2116 35334
rect 2172 35332 2196 35334
rect 2252 35332 2258 35334
rect 1950 35323 2258 35332
rect 1950 34300 2258 34309
rect 1950 34298 1956 34300
rect 2012 34298 2036 34300
rect 2092 34298 2116 34300
rect 2172 34298 2196 34300
rect 2252 34298 2258 34300
rect 2012 34246 2014 34298
rect 2194 34246 2196 34298
rect 1950 34244 1956 34246
rect 2012 34244 2036 34246
rect 2092 34244 2116 34246
rect 2172 34244 2196 34246
rect 2252 34244 2258 34246
rect 1950 34235 2258 34244
rect 1950 33212 2258 33221
rect 1950 33210 1956 33212
rect 2012 33210 2036 33212
rect 2092 33210 2116 33212
rect 2172 33210 2196 33212
rect 2252 33210 2258 33212
rect 2012 33158 2014 33210
rect 2194 33158 2196 33210
rect 1950 33156 1956 33158
rect 2012 33156 2036 33158
rect 2092 33156 2116 33158
rect 2172 33156 2196 33158
rect 2252 33156 2258 33158
rect 1950 33147 2258 33156
rect 1950 32124 2258 32133
rect 1950 32122 1956 32124
rect 2012 32122 2036 32124
rect 2092 32122 2116 32124
rect 2172 32122 2196 32124
rect 2252 32122 2258 32124
rect 2012 32070 2014 32122
rect 2194 32070 2196 32122
rect 1950 32068 1956 32070
rect 2012 32068 2036 32070
rect 2092 32068 2116 32070
rect 2172 32068 2196 32070
rect 2252 32068 2258 32070
rect 1950 32059 2258 32068
rect 1950 31036 2258 31045
rect 1950 31034 1956 31036
rect 2012 31034 2036 31036
rect 2092 31034 2116 31036
rect 2172 31034 2196 31036
rect 2252 31034 2258 31036
rect 2012 30982 2014 31034
rect 2194 30982 2196 31034
rect 1950 30980 1956 30982
rect 2012 30980 2036 30982
rect 2092 30980 2116 30982
rect 2172 30980 2196 30982
rect 2252 30980 2258 30982
rect 1950 30971 2258 30980
rect 1950 29948 2258 29957
rect 1950 29946 1956 29948
rect 2012 29946 2036 29948
rect 2092 29946 2116 29948
rect 2172 29946 2196 29948
rect 2252 29946 2258 29948
rect 2012 29894 2014 29946
rect 2194 29894 2196 29946
rect 1950 29892 1956 29894
rect 2012 29892 2036 29894
rect 2092 29892 2116 29894
rect 2172 29892 2196 29894
rect 2252 29892 2258 29894
rect 1950 29883 2258 29892
rect 1950 28860 2258 28869
rect 1950 28858 1956 28860
rect 2012 28858 2036 28860
rect 2092 28858 2116 28860
rect 2172 28858 2196 28860
rect 2252 28858 2258 28860
rect 2012 28806 2014 28858
rect 2194 28806 2196 28858
rect 1950 28804 1956 28806
rect 2012 28804 2036 28806
rect 2092 28804 2116 28806
rect 2172 28804 2196 28806
rect 2252 28804 2258 28806
rect 1950 28795 2258 28804
rect 1950 27772 2258 27781
rect 1950 27770 1956 27772
rect 2012 27770 2036 27772
rect 2092 27770 2116 27772
rect 2172 27770 2196 27772
rect 2252 27770 2258 27772
rect 2012 27718 2014 27770
rect 2194 27718 2196 27770
rect 1950 27716 1956 27718
rect 2012 27716 2036 27718
rect 2092 27716 2116 27718
rect 2172 27716 2196 27718
rect 2252 27716 2258 27718
rect 1950 27707 2258 27716
rect 1950 26684 2258 26693
rect 1950 26682 1956 26684
rect 2012 26682 2036 26684
rect 2092 26682 2116 26684
rect 2172 26682 2196 26684
rect 2252 26682 2258 26684
rect 2012 26630 2014 26682
rect 2194 26630 2196 26682
rect 1950 26628 1956 26630
rect 2012 26628 2036 26630
rect 2092 26628 2116 26630
rect 2172 26628 2196 26630
rect 2252 26628 2258 26630
rect 1950 26619 2258 26628
rect 1950 25596 2258 25605
rect 1950 25594 1956 25596
rect 2012 25594 2036 25596
rect 2092 25594 2116 25596
rect 2172 25594 2196 25596
rect 2252 25594 2258 25596
rect 2012 25542 2014 25594
rect 2194 25542 2196 25594
rect 1950 25540 1956 25542
rect 2012 25540 2036 25542
rect 2092 25540 2116 25542
rect 2172 25540 2196 25542
rect 2252 25540 2258 25542
rect 1950 25531 2258 25540
rect 1950 24508 2258 24517
rect 1950 24506 1956 24508
rect 2012 24506 2036 24508
rect 2092 24506 2116 24508
rect 2172 24506 2196 24508
rect 2252 24506 2258 24508
rect 2012 24454 2014 24506
rect 2194 24454 2196 24506
rect 1950 24452 1956 24454
rect 2012 24452 2036 24454
rect 2092 24452 2116 24454
rect 2172 24452 2196 24454
rect 2252 24452 2258 24454
rect 1950 24443 2258 24452
rect 2332 23594 2360 67662
rect 2412 64932 2464 64938
rect 2412 64874 2464 64880
rect 2424 31210 2452 64874
rect 2516 56778 2544 67798
rect 2610 67484 2918 67493
rect 2610 67482 2616 67484
rect 2672 67482 2696 67484
rect 2752 67482 2776 67484
rect 2832 67482 2856 67484
rect 2912 67482 2918 67484
rect 2672 67430 2674 67482
rect 2854 67430 2856 67482
rect 2610 67428 2616 67430
rect 2672 67428 2696 67430
rect 2752 67428 2776 67430
rect 2832 67428 2856 67430
rect 2912 67428 2918 67430
rect 2610 67419 2918 67428
rect 2610 66396 2918 66405
rect 2610 66394 2616 66396
rect 2672 66394 2696 66396
rect 2752 66394 2776 66396
rect 2832 66394 2856 66396
rect 2912 66394 2918 66396
rect 2672 66342 2674 66394
rect 2854 66342 2856 66394
rect 2610 66340 2616 66342
rect 2672 66340 2696 66342
rect 2752 66340 2776 66342
rect 2832 66340 2856 66342
rect 2912 66340 2918 66342
rect 2610 66331 2918 66340
rect 2610 65308 2918 65317
rect 2610 65306 2616 65308
rect 2672 65306 2696 65308
rect 2752 65306 2776 65308
rect 2832 65306 2856 65308
rect 2912 65306 2918 65308
rect 2672 65254 2674 65306
rect 2854 65254 2856 65306
rect 2610 65252 2616 65254
rect 2672 65252 2696 65254
rect 2752 65252 2776 65254
rect 2832 65252 2856 65254
rect 2912 65252 2918 65254
rect 2610 65243 2918 65252
rect 2610 64220 2918 64229
rect 2610 64218 2616 64220
rect 2672 64218 2696 64220
rect 2752 64218 2776 64220
rect 2832 64218 2856 64220
rect 2912 64218 2918 64220
rect 2672 64166 2674 64218
rect 2854 64166 2856 64218
rect 2610 64164 2616 64166
rect 2672 64164 2696 64166
rect 2752 64164 2776 64166
rect 2832 64164 2856 64166
rect 2912 64164 2918 64166
rect 2610 64155 2918 64164
rect 2610 63132 2918 63141
rect 2610 63130 2616 63132
rect 2672 63130 2696 63132
rect 2752 63130 2776 63132
rect 2832 63130 2856 63132
rect 2912 63130 2918 63132
rect 2672 63078 2674 63130
rect 2854 63078 2856 63130
rect 2610 63076 2616 63078
rect 2672 63076 2696 63078
rect 2752 63076 2776 63078
rect 2832 63076 2856 63078
rect 2912 63076 2918 63078
rect 2610 63067 2918 63076
rect 2610 62044 2918 62053
rect 2610 62042 2616 62044
rect 2672 62042 2696 62044
rect 2752 62042 2776 62044
rect 2832 62042 2856 62044
rect 2912 62042 2918 62044
rect 2672 61990 2674 62042
rect 2854 61990 2856 62042
rect 2610 61988 2616 61990
rect 2672 61988 2696 61990
rect 2752 61988 2776 61990
rect 2832 61988 2856 61990
rect 2912 61988 2918 61990
rect 2610 61979 2918 61988
rect 2610 60956 2918 60965
rect 2610 60954 2616 60956
rect 2672 60954 2696 60956
rect 2752 60954 2776 60956
rect 2832 60954 2856 60956
rect 2912 60954 2918 60956
rect 2672 60902 2674 60954
rect 2854 60902 2856 60954
rect 2610 60900 2616 60902
rect 2672 60900 2696 60902
rect 2752 60900 2776 60902
rect 2832 60900 2856 60902
rect 2912 60900 2918 60902
rect 2610 60891 2918 60900
rect 2610 59868 2918 59877
rect 2610 59866 2616 59868
rect 2672 59866 2696 59868
rect 2752 59866 2776 59868
rect 2832 59866 2856 59868
rect 2912 59866 2918 59868
rect 2672 59814 2674 59866
rect 2854 59814 2856 59866
rect 2610 59812 2616 59814
rect 2672 59812 2696 59814
rect 2752 59812 2776 59814
rect 2832 59812 2856 59814
rect 2912 59812 2918 59814
rect 2610 59803 2918 59812
rect 2610 58780 2918 58789
rect 2610 58778 2616 58780
rect 2672 58778 2696 58780
rect 2752 58778 2776 58780
rect 2832 58778 2856 58780
rect 2912 58778 2918 58780
rect 2672 58726 2674 58778
rect 2854 58726 2856 58778
rect 2610 58724 2616 58726
rect 2672 58724 2696 58726
rect 2752 58724 2776 58726
rect 2832 58724 2856 58726
rect 2912 58724 2918 58726
rect 2610 58715 2918 58724
rect 3344 57866 3372 69362
rect 6950 69116 7258 69125
rect 6950 69114 6956 69116
rect 7012 69114 7036 69116
rect 7092 69114 7116 69116
rect 7172 69114 7196 69116
rect 7252 69114 7258 69116
rect 7012 69062 7014 69114
rect 7194 69062 7196 69114
rect 6950 69060 6956 69062
rect 7012 69060 7036 69062
rect 7092 69060 7116 69062
rect 7172 69060 7196 69062
rect 7252 69060 7258 69062
rect 6950 69051 7258 69060
rect 7610 68572 7918 68581
rect 7610 68570 7616 68572
rect 7672 68570 7696 68572
rect 7752 68570 7776 68572
rect 7832 68570 7856 68572
rect 7912 68570 7918 68572
rect 7672 68518 7674 68570
rect 7854 68518 7856 68570
rect 7610 68516 7616 68518
rect 7672 68516 7696 68518
rect 7752 68516 7776 68518
rect 7832 68516 7856 68518
rect 7912 68516 7918 68518
rect 7610 68507 7918 68516
rect 9128 68400 9180 68406
rect 9128 68342 9180 68348
rect 6828 68332 6880 68338
rect 6828 68274 6880 68280
rect 7288 68332 7340 68338
rect 7288 68274 7340 68280
rect 6368 67652 6420 67658
rect 6368 67594 6420 67600
rect 3608 66156 3660 66162
rect 3608 66098 3660 66104
rect 3620 63374 3648 66098
rect 5724 63980 5776 63986
rect 5724 63922 5776 63928
rect 4068 63572 4120 63578
rect 4068 63514 4120 63520
rect 3608 63368 3660 63374
rect 3608 63310 3660 63316
rect 3332 57860 3384 57866
rect 3332 57802 3384 57808
rect 2610 57692 2918 57701
rect 2610 57690 2616 57692
rect 2672 57690 2696 57692
rect 2752 57690 2776 57692
rect 2832 57690 2856 57692
rect 2912 57690 2918 57692
rect 2672 57638 2674 57690
rect 2854 57638 2856 57690
rect 2610 57636 2616 57638
rect 2672 57636 2696 57638
rect 2752 57636 2776 57638
rect 2832 57636 2856 57638
rect 2912 57636 2918 57638
rect 2610 57627 2918 57636
rect 2504 56772 2556 56778
rect 2504 56714 2556 56720
rect 2610 56604 2918 56613
rect 2610 56602 2616 56604
rect 2672 56602 2696 56604
rect 2752 56602 2776 56604
rect 2832 56602 2856 56604
rect 2912 56602 2918 56604
rect 2672 56550 2674 56602
rect 2854 56550 2856 56602
rect 2610 56548 2616 56550
rect 2672 56548 2696 56550
rect 2752 56548 2776 56550
rect 2832 56548 2856 56550
rect 2912 56548 2918 56550
rect 2610 56539 2918 56548
rect 2610 55516 2918 55525
rect 2610 55514 2616 55516
rect 2672 55514 2696 55516
rect 2752 55514 2776 55516
rect 2832 55514 2856 55516
rect 2912 55514 2918 55516
rect 2672 55462 2674 55514
rect 2854 55462 2856 55514
rect 2610 55460 2616 55462
rect 2672 55460 2696 55462
rect 2752 55460 2776 55462
rect 2832 55460 2856 55462
rect 2912 55460 2918 55462
rect 2610 55451 2918 55460
rect 2610 54428 2918 54437
rect 2610 54426 2616 54428
rect 2672 54426 2696 54428
rect 2752 54426 2776 54428
rect 2832 54426 2856 54428
rect 2912 54426 2918 54428
rect 2672 54374 2674 54426
rect 2854 54374 2856 54426
rect 2610 54372 2616 54374
rect 2672 54372 2696 54374
rect 2752 54372 2776 54374
rect 2832 54372 2856 54374
rect 2912 54372 2918 54374
rect 2610 54363 2918 54372
rect 2610 53340 2918 53349
rect 2610 53338 2616 53340
rect 2672 53338 2696 53340
rect 2752 53338 2776 53340
rect 2832 53338 2856 53340
rect 2912 53338 2918 53340
rect 2672 53286 2674 53338
rect 2854 53286 2856 53338
rect 2610 53284 2616 53286
rect 2672 53284 2696 53286
rect 2752 53284 2776 53286
rect 2832 53284 2856 53286
rect 2912 53284 2918 53286
rect 2610 53275 2918 53284
rect 2610 52252 2918 52261
rect 2610 52250 2616 52252
rect 2672 52250 2696 52252
rect 2752 52250 2776 52252
rect 2832 52250 2856 52252
rect 2912 52250 2918 52252
rect 2672 52198 2674 52250
rect 2854 52198 2856 52250
rect 2610 52196 2616 52198
rect 2672 52196 2696 52198
rect 2752 52196 2776 52198
rect 2832 52196 2856 52198
rect 2912 52196 2918 52198
rect 2610 52187 2918 52196
rect 2610 51164 2918 51173
rect 2610 51162 2616 51164
rect 2672 51162 2696 51164
rect 2752 51162 2776 51164
rect 2832 51162 2856 51164
rect 2912 51162 2918 51164
rect 2672 51110 2674 51162
rect 2854 51110 2856 51162
rect 2610 51108 2616 51110
rect 2672 51108 2696 51110
rect 2752 51108 2776 51110
rect 2832 51108 2856 51110
rect 2912 51108 2918 51110
rect 2610 51099 2918 51108
rect 2610 50076 2918 50085
rect 2610 50074 2616 50076
rect 2672 50074 2696 50076
rect 2752 50074 2776 50076
rect 2832 50074 2856 50076
rect 2912 50074 2918 50076
rect 2672 50022 2674 50074
rect 2854 50022 2856 50074
rect 2610 50020 2616 50022
rect 2672 50020 2696 50022
rect 2752 50020 2776 50022
rect 2832 50020 2856 50022
rect 2912 50020 2918 50022
rect 2610 50011 2918 50020
rect 2610 48988 2918 48997
rect 2610 48986 2616 48988
rect 2672 48986 2696 48988
rect 2752 48986 2776 48988
rect 2832 48986 2856 48988
rect 2912 48986 2918 48988
rect 2672 48934 2674 48986
rect 2854 48934 2856 48986
rect 2610 48932 2616 48934
rect 2672 48932 2696 48934
rect 2752 48932 2776 48934
rect 2832 48932 2856 48934
rect 2912 48932 2918 48934
rect 2610 48923 2918 48932
rect 3424 48204 3476 48210
rect 3424 48146 3476 48152
rect 2610 47900 2918 47909
rect 2610 47898 2616 47900
rect 2672 47898 2696 47900
rect 2752 47898 2776 47900
rect 2832 47898 2856 47900
rect 2912 47898 2918 47900
rect 2672 47846 2674 47898
rect 2854 47846 2856 47898
rect 2610 47844 2616 47846
rect 2672 47844 2696 47846
rect 2752 47844 2776 47846
rect 2832 47844 2856 47846
rect 2912 47844 2918 47846
rect 2610 47835 2918 47844
rect 2610 46812 2918 46821
rect 2610 46810 2616 46812
rect 2672 46810 2696 46812
rect 2752 46810 2776 46812
rect 2832 46810 2856 46812
rect 2912 46810 2918 46812
rect 2672 46758 2674 46810
rect 2854 46758 2856 46810
rect 2610 46756 2616 46758
rect 2672 46756 2696 46758
rect 2752 46756 2776 46758
rect 2832 46756 2856 46758
rect 2912 46756 2918 46758
rect 2610 46747 2918 46756
rect 2610 45724 2918 45733
rect 2610 45722 2616 45724
rect 2672 45722 2696 45724
rect 2752 45722 2776 45724
rect 2832 45722 2856 45724
rect 2912 45722 2918 45724
rect 2672 45670 2674 45722
rect 2854 45670 2856 45722
rect 2610 45668 2616 45670
rect 2672 45668 2696 45670
rect 2752 45668 2776 45670
rect 2832 45668 2856 45670
rect 2912 45668 2918 45670
rect 2610 45659 2918 45668
rect 3056 45552 3108 45558
rect 3056 45494 3108 45500
rect 3068 44946 3096 45494
rect 3148 45416 3200 45422
rect 3148 45358 3200 45364
rect 3056 44940 3108 44946
rect 3056 44882 3108 44888
rect 2504 44804 2556 44810
rect 2504 44746 2556 44752
rect 2412 31204 2464 31210
rect 2412 31146 2464 31152
rect 2320 23588 2372 23594
rect 2320 23530 2372 23536
rect 1950 23420 2258 23429
rect 1950 23418 1956 23420
rect 2012 23418 2036 23420
rect 2092 23418 2116 23420
rect 2172 23418 2196 23420
rect 2252 23418 2258 23420
rect 2012 23366 2014 23418
rect 2194 23366 2196 23418
rect 1950 23364 1956 23366
rect 2012 23364 2036 23366
rect 2092 23364 2116 23366
rect 2172 23364 2196 23366
rect 2252 23364 2258 23366
rect 1950 23355 2258 23364
rect 1950 22332 2258 22341
rect 1950 22330 1956 22332
rect 2012 22330 2036 22332
rect 2092 22330 2116 22332
rect 2172 22330 2196 22332
rect 2252 22330 2258 22332
rect 2012 22278 2014 22330
rect 2194 22278 2196 22330
rect 1950 22276 1956 22278
rect 2012 22276 2036 22278
rect 2092 22276 2116 22278
rect 2172 22276 2196 22278
rect 2252 22276 2258 22278
rect 1950 22267 2258 22276
rect 1950 21244 2258 21253
rect 1950 21242 1956 21244
rect 2012 21242 2036 21244
rect 2092 21242 2116 21244
rect 2172 21242 2196 21244
rect 2252 21242 2258 21244
rect 2012 21190 2014 21242
rect 2194 21190 2196 21242
rect 1950 21188 1956 21190
rect 2012 21188 2036 21190
rect 2092 21188 2116 21190
rect 2172 21188 2196 21190
rect 2252 21188 2258 21190
rect 1950 21179 2258 21188
rect 1950 20156 2258 20165
rect 1950 20154 1956 20156
rect 2012 20154 2036 20156
rect 2092 20154 2116 20156
rect 2172 20154 2196 20156
rect 2252 20154 2258 20156
rect 2012 20102 2014 20154
rect 2194 20102 2196 20154
rect 1950 20100 1956 20102
rect 2012 20100 2036 20102
rect 2092 20100 2116 20102
rect 2172 20100 2196 20102
rect 2252 20100 2258 20102
rect 1950 20091 2258 20100
rect 1860 19304 1912 19310
rect 1860 19246 1912 19252
rect 1950 19068 2258 19077
rect 1950 19066 1956 19068
rect 2012 19066 2036 19068
rect 2092 19066 2116 19068
rect 2172 19066 2196 19068
rect 2252 19066 2258 19068
rect 2012 19014 2014 19066
rect 2194 19014 2196 19066
rect 1950 19012 1956 19014
rect 2012 19012 2036 19014
rect 2092 19012 2116 19014
rect 2172 19012 2196 19014
rect 2252 19012 2258 19014
rect 1950 19003 2258 19012
rect 1676 18080 1728 18086
rect 1676 18022 1728 18028
rect 1950 17980 2258 17989
rect 1950 17978 1956 17980
rect 2012 17978 2036 17980
rect 2092 17978 2116 17980
rect 2172 17978 2196 17980
rect 2252 17978 2258 17980
rect 2012 17926 2014 17978
rect 2194 17926 2196 17978
rect 1950 17924 1956 17926
rect 2012 17924 2036 17926
rect 2092 17924 2116 17926
rect 2172 17924 2196 17926
rect 2252 17924 2258 17926
rect 1950 17915 2258 17924
rect 1676 16992 1728 16998
rect 1676 16934 1728 16940
rect 1688 3602 1716 16934
rect 1950 16892 2258 16901
rect 1950 16890 1956 16892
rect 2012 16890 2036 16892
rect 2092 16890 2116 16892
rect 2172 16890 2196 16892
rect 2252 16890 2258 16892
rect 2012 16838 2014 16890
rect 2194 16838 2196 16890
rect 1950 16836 1956 16838
rect 2012 16836 2036 16838
rect 2092 16836 2116 16838
rect 2172 16836 2196 16838
rect 2252 16836 2258 16838
rect 1950 16827 2258 16836
rect 1950 15804 2258 15813
rect 1950 15802 1956 15804
rect 2012 15802 2036 15804
rect 2092 15802 2116 15804
rect 2172 15802 2196 15804
rect 2252 15802 2258 15804
rect 2012 15750 2014 15802
rect 2194 15750 2196 15802
rect 1950 15748 1956 15750
rect 2012 15748 2036 15750
rect 2092 15748 2116 15750
rect 2172 15748 2196 15750
rect 2252 15748 2258 15750
rect 1950 15739 2258 15748
rect 1950 14716 2258 14725
rect 1950 14714 1956 14716
rect 2012 14714 2036 14716
rect 2092 14714 2116 14716
rect 2172 14714 2196 14716
rect 2252 14714 2258 14716
rect 2012 14662 2014 14714
rect 2194 14662 2196 14714
rect 1950 14660 1956 14662
rect 2012 14660 2036 14662
rect 2092 14660 2116 14662
rect 2172 14660 2196 14662
rect 2252 14660 2258 14662
rect 1950 14651 2258 14660
rect 1950 13628 2258 13637
rect 1950 13626 1956 13628
rect 2012 13626 2036 13628
rect 2092 13626 2116 13628
rect 2172 13626 2196 13628
rect 2252 13626 2258 13628
rect 2012 13574 2014 13626
rect 2194 13574 2196 13626
rect 1950 13572 1956 13574
rect 2012 13572 2036 13574
rect 2092 13572 2116 13574
rect 2172 13572 2196 13574
rect 2252 13572 2258 13574
rect 1950 13563 2258 13572
rect 1950 12540 2258 12549
rect 1950 12538 1956 12540
rect 2012 12538 2036 12540
rect 2092 12538 2116 12540
rect 2172 12538 2196 12540
rect 2252 12538 2258 12540
rect 2012 12486 2014 12538
rect 2194 12486 2196 12538
rect 1950 12484 1956 12486
rect 2012 12484 2036 12486
rect 2092 12484 2116 12486
rect 2172 12484 2196 12486
rect 2252 12484 2258 12486
rect 1950 12475 2258 12484
rect 1950 11452 2258 11461
rect 1950 11450 1956 11452
rect 2012 11450 2036 11452
rect 2092 11450 2116 11452
rect 2172 11450 2196 11452
rect 2252 11450 2258 11452
rect 2012 11398 2014 11450
rect 2194 11398 2196 11450
rect 1950 11396 1956 11398
rect 2012 11396 2036 11398
rect 2092 11396 2116 11398
rect 2172 11396 2196 11398
rect 2252 11396 2258 11398
rect 1950 11387 2258 11396
rect 1950 10364 2258 10373
rect 1950 10362 1956 10364
rect 2012 10362 2036 10364
rect 2092 10362 2116 10364
rect 2172 10362 2196 10364
rect 2252 10362 2258 10364
rect 2012 10310 2014 10362
rect 2194 10310 2196 10362
rect 1950 10308 1956 10310
rect 2012 10308 2036 10310
rect 2092 10308 2116 10310
rect 2172 10308 2196 10310
rect 2252 10308 2258 10310
rect 1950 10299 2258 10308
rect 1950 9276 2258 9285
rect 1950 9274 1956 9276
rect 2012 9274 2036 9276
rect 2092 9274 2116 9276
rect 2172 9274 2196 9276
rect 2252 9274 2258 9276
rect 2012 9222 2014 9274
rect 2194 9222 2196 9274
rect 1950 9220 1956 9222
rect 2012 9220 2036 9222
rect 2092 9220 2116 9222
rect 2172 9220 2196 9222
rect 2252 9220 2258 9222
rect 1950 9211 2258 9220
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 2516 4010 2544 44746
rect 2610 44636 2918 44645
rect 2610 44634 2616 44636
rect 2672 44634 2696 44636
rect 2752 44634 2776 44636
rect 2832 44634 2856 44636
rect 2912 44634 2918 44636
rect 2672 44582 2674 44634
rect 2854 44582 2856 44634
rect 2610 44580 2616 44582
rect 2672 44580 2696 44582
rect 2752 44580 2776 44582
rect 2832 44580 2856 44582
rect 2912 44580 2918 44582
rect 2610 44571 2918 44580
rect 2610 43548 2918 43557
rect 2610 43546 2616 43548
rect 2672 43546 2696 43548
rect 2752 43546 2776 43548
rect 2832 43546 2856 43548
rect 2912 43546 2918 43548
rect 2672 43494 2674 43546
rect 2854 43494 2856 43546
rect 2610 43492 2616 43494
rect 2672 43492 2696 43494
rect 2752 43492 2776 43494
rect 2832 43492 2856 43494
rect 2912 43492 2918 43494
rect 2610 43483 2918 43492
rect 2610 42460 2918 42469
rect 2610 42458 2616 42460
rect 2672 42458 2696 42460
rect 2752 42458 2776 42460
rect 2832 42458 2856 42460
rect 2912 42458 2918 42460
rect 2672 42406 2674 42458
rect 2854 42406 2856 42458
rect 2610 42404 2616 42406
rect 2672 42404 2696 42406
rect 2752 42404 2776 42406
rect 2832 42404 2856 42406
rect 2912 42404 2918 42406
rect 2610 42395 2918 42404
rect 2610 41372 2918 41381
rect 2610 41370 2616 41372
rect 2672 41370 2696 41372
rect 2752 41370 2776 41372
rect 2832 41370 2856 41372
rect 2912 41370 2918 41372
rect 2672 41318 2674 41370
rect 2854 41318 2856 41370
rect 2610 41316 2616 41318
rect 2672 41316 2696 41318
rect 2752 41316 2776 41318
rect 2832 41316 2856 41318
rect 2912 41316 2918 41318
rect 2610 41307 2918 41316
rect 2610 40284 2918 40293
rect 2610 40282 2616 40284
rect 2672 40282 2696 40284
rect 2752 40282 2776 40284
rect 2832 40282 2856 40284
rect 2912 40282 2918 40284
rect 2672 40230 2674 40282
rect 2854 40230 2856 40282
rect 2610 40228 2616 40230
rect 2672 40228 2696 40230
rect 2752 40228 2776 40230
rect 2832 40228 2856 40230
rect 2912 40228 2918 40230
rect 2610 40219 2918 40228
rect 2610 39196 2918 39205
rect 2610 39194 2616 39196
rect 2672 39194 2696 39196
rect 2752 39194 2776 39196
rect 2832 39194 2856 39196
rect 2912 39194 2918 39196
rect 2672 39142 2674 39194
rect 2854 39142 2856 39194
rect 2610 39140 2616 39142
rect 2672 39140 2696 39142
rect 2752 39140 2776 39142
rect 2832 39140 2856 39142
rect 2912 39140 2918 39142
rect 2610 39131 2918 39140
rect 2610 38108 2918 38117
rect 2610 38106 2616 38108
rect 2672 38106 2696 38108
rect 2752 38106 2776 38108
rect 2832 38106 2856 38108
rect 2912 38106 2918 38108
rect 2672 38054 2674 38106
rect 2854 38054 2856 38106
rect 2610 38052 2616 38054
rect 2672 38052 2696 38054
rect 2752 38052 2776 38054
rect 2832 38052 2856 38054
rect 2912 38052 2918 38054
rect 2610 38043 2918 38052
rect 2610 37020 2918 37029
rect 2610 37018 2616 37020
rect 2672 37018 2696 37020
rect 2752 37018 2776 37020
rect 2832 37018 2856 37020
rect 2912 37018 2918 37020
rect 2672 36966 2674 37018
rect 2854 36966 2856 37018
rect 2610 36964 2616 36966
rect 2672 36964 2696 36966
rect 2752 36964 2776 36966
rect 2832 36964 2856 36966
rect 2912 36964 2918 36966
rect 2610 36955 2918 36964
rect 2610 35932 2918 35941
rect 2610 35930 2616 35932
rect 2672 35930 2696 35932
rect 2752 35930 2776 35932
rect 2832 35930 2856 35932
rect 2912 35930 2918 35932
rect 2672 35878 2674 35930
rect 2854 35878 2856 35930
rect 2610 35876 2616 35878
rect 2672 35876 2696 35878
rect 2752 35876 2776 35878
rect 2832 35876 2856 35878
rect 2912 35876 2918 35878
rect 2610 35867 2918 35876
rect 2610 34844 2918 34853
rect 2610 34842 2616 34844
rect 2672 34842 2696 34844
rect 2752 34842 2776 34844
rect 2832 34842 2856 34844
rect 2912 34842 2918 34844
rect 2672 34790 2674 34842
rect 2854 34790 2856 34842
rect 2610 34788 2616 34790
rect 2672 34788 2696 34790
rect 2752 34788 2776 34790
rect 2832 34788 2856 34790
rect 2912 34788 2918 34790
rect 2610 34779 2918 34788
rect 2610 33756 2918 33765
rect 2610 33754 2616 33756
rect 2672 33754 2696 33756
rect 2752 33754 2776 33756
rect 2832 33754 2856 33756
rect 2912 33754 2918 33756
rect 2672 33702 2674 33754
rect 2854 33702 2856 33754
rect 2610 33700 2616 33702
rect 2672 33700 2696 33702
rect 2752 33700 2776 33702
rect 2832 33700 2856 33702
rect 2912 33700 2918 33702
rect 2610 33691 2918 33700
rect 2610 32668 2918 32677
rect 2610 32666 2616 32668
rect 2672 32666 2696 32668
rect 2752 32666 2776 32668
rect 2832 32666 2856 32668
rect 2912 32666 2918 32668
rect 2672 32614 2674 32666
rect 2854 32614 2856 32666
rect 2610 32612 2616 32614
rect 2672 32612 2696 32614
rect 2752 32612 2776 32614
rect 2832 32612 2856 32614
rect 2912 32612 2918 32614
rect 2610 32603 2918 32612
rect 2610 31580 2918 31589
rect 2610 31578 2616 31580
rect 2672 31578 2696 31580
rect 2752 31578 2776 31580
rect 2832 31578 2856 31580
rect 2912 31578 2918 31580
rect 2672 31526 2674 31578
rect 2854 31526 2856 31578
rect 2610 31524 2616 31526
rect 2672 31524 2696 31526
rect 2752 31524 2776 31526
rect 2832 31524 2856 31526
rect 2912 31524 2918 31526
rect 2610 31515 2918 31524
rect 2610 30492 2918 30501
rect 2610 30490 2616 30492
rect 2672 30490 2696 30492
rect 2752 30490 2776 30492
rect 2832 30490 2856 30492
rect 2912 30490 2918 30492
rect 2672 30438 2674 30490
rect 2854 30438 2856 30490
rect 2610 30436 2616 30438
rect 2672 30436 2696 30438
rect 2752 30436 2776 30438
rect 2832 30436 2856 30438
rect 2912 30436 2918 30438
rect 2610 30427 2918 30436
rect 3056 30388 3108 30394
rect 3056 30330 3108 30336
rect 2610 29404 2918 29413
rect 2610 29402 2616 29404
rect 2672 29402 2696 29404
rect 2752 29402 2776 29404
rect 2832 29402 2856 29404
rect 2912 29402 2918 29404
rect 2672 29350 2674 29402
rect 2854 29350 2856 29402
rect 2610 29348 2616 29350
rect 2672 29348 2696 29350
rect 2752 29348 2776 29350
rect 2832 29348 2856 29350
rect 2912 29348 2918 29350
rect 2610 29339 2918 29348
rect 2610 28316 2918 28325
rect 2610 28314 2616 28316
rect 2672 28314 2696 28316
rect 2752 28314 2776 28316
rect 2832 28314 2856 28316
rect 2912 28314 2918 28316
rect 2672 28262 2674 28314
rect 2854 28262 2856 28314
rect 2610 28260 2616 28262
rect 2672 28260 2696 28262
rect 2752 28260 2776 28262
rect 2832 28260 2856 28262
rect 2912 28260 2918 28262
rect 2610 28251 2918 28260
rect 2610 27228 2918 27237
rect 2610 27226 2616 27228
rect 2672 27226 2696 27228
rect 2752 27226 2776 27228
rect 2832 27226 2856 27228
rect 2912 27226 2918 27228
rect 2672 27174 2674 27226
rect 2854 27174 2856 27226
rect 2610 27172 2616 27174
rect 2672 27172 2696 27174
rect 2752 27172 2776 27174
rect 2832 27172 2856 27174
rect 2912 27172 2918 27174
rect 2610 27163 2918 27172
rect 2610 26140 2918 26149
rect 2610 26138 2616 26140
rect 2672 26138 2696 26140
rect 2752 26138 2776 26140
rect 2832 26138 2856 26140
rect 2912 26138 2918 26140
rect 2672 26086 2674 26138
rect 2854 26086 2856 26138
rect 2610 26084 2616 26086
rect 2672 26084 2696 26086
rect 2752 26084 2776 26086
rect 2832 26084 2856 26086
rect 2912 26084 2918 26086
rect 2610 26075 2918 26084
rect 2610 25052 2918 25061
rect 2610 25050 2616 25052
rect 2672 25050 2696 25052
rect 2752 25050 2776 25052
rect 2832 25050 2856 25052
rect 2912 25050 2918 25052
rect 2672 24998 2674 25050
rect 2854 24998 2856 25050
rect 2610 24996 2616 24998
rect 2672 24996 2696 24998
rect 2752 24996 2776 24998
rect 2832 24996 2856 24998
rect 2912 24996 2918 24998
rect 2610 24987 2918 24996
rect 2610 23964 2918 23973
rect 2610 23962 2616 23964
rect 2672 23962 2696 23964
rect 2752 23962 2776 23964
rect 2832 23962 2856 23964
rect 2912 23962 2918 23964
rect 2672 23910 2674 23962
rect 2854 23910 2856 23962
rect 2610 23908 2616 23910
rect 2672 23908 2696 23910
rect 2752 23908 2776 23910
rect 2832 23908 2856 23910
rect 2912 23908 2918 23910
rect 2610 23899 2918 23908
rect 2610 22876 2918 22885
rect 2610 22874 2616 22876
rect 2672 22874 2696 22876
rect 2752 22874 2776 22876
rect 2832 22874 2856 22876
rect 2912 22874 2918 22876
rect 2672 22822 2674 22874
rect 2854 22822 2856 22874
rect 2610 22820 2616 22822
rect 2672 22820 2696 22822
rect 2752 22820 2776 22822
rect 2832 22820 2856 22822
rect 2912 22820 2918 22822
rect 2610 22811 2918 22820
rect 2610 21788 2918 21797
rect 2610 21786 2616 21788
rect 2672 21786 2696 21788
rect 2752 21786 2776 21788
rect 2832 21786 2856 21788
rect 2912 21786 2918 21788
rect 2672 21734 2674 21786
rect 2854 21734 2856 21786
rect 2610 21732 2616 21734
rect 2672 21732 2696 21734
rect 2752 21732 2776 21734
rect 2832 21732 2856 21734
rect 2912 21732 2918 21734
rect 2610 21723 2918 21732
rect 2610 20700 2918 20709
rect 2610 20698 2616 20700
rect 2672 20698 2696 20700
rect 2752 20698 2776 20700
rect 2832 20698 2856 20700
rect 2912 20698 2918 20700
rect 2672 20646 2674 20698
rect 2854 20646 2856 20698
rect 2610 20644 2616 20646
rect 2672 20644 2696 20646
rect 2752 20644 2776 20646
rect 2832 20644 2856 20646
rect 2912 20644 2918 20646
rect 2610 20635 2918 20644
rect 2610 19612 2918 19621
rect 2610 19610 2616 19612
rect 2672 19610 2696 19612
rect 2752 19610 2776 19612
rect 2832 19610 2856 19612
rect 2912 19610 2918 19612
rect 2672 19558 2674 19610
rect 2854 19558 2856 19610
rect 2610 19556 2616 19558
rect 2672 19556 2696 19558
rect 2752 19556 2776 19558
rect 2832 19556 2856 19558
rect 2912 19556 2918 19558
rect 2610 19547 2918 19556
rect 2610 18524 2918 18533
rect 2610 18522 2616 18524
rect 2672 18522 2696 18524
rect 2752 18522 2776 18524
rect 2832 18522 2856 18524
rect 2912 18522 2918 18524
rect 2672 18470 2674 18522
rect 2854 18470 2856 18522
rect 2610 18468 2616 18470
rect 2672 18468 2696 18470
rect 2752 18468 2776 18470
rect 2832 18468 2856 18470
rect 2912 18468 2918 18470
rect 2610 18459 2918 18468
rect 2964 17536 3016 17542
rect 2964 17478 3016 17484
rect 2610 17436 2918 17445
rect 2610 17434 2616 17436
rect 2672 17434 2696 17436
rect 2752 17434 2776 17436
rect 2832 17434 2856 17436
rect 2912 17434 2918 17436
rect 2672 17382 2674 17434
rect 2854 17382 2856 17434
rect 2610 17380 2616 17382
rect 2672 17380 2696 17382
rect 2752 17380 2776 17382
rect 2832 17380 2856 17382
rect 2912 17380 2918 17382
rect 2610 17371 2918 17380
rect 2976 17270 3004 17478
rect 2964 17264 3016 17270
rect 2964 17206 3016 17212
rect 2610 16348 2918 16357
rect 2610 16346 2616 16348
rect 2672 16346 2696 16348
rect 2752 16346 2776 16348
rect 2832 16346 2856 16348
rect 2912 16346 2918 16348
rect 2672 16294 2674 16346
rect 2854 16294 2856 16346
rect 2610 16292 2616 16294
rect 2672 16292 2696 16294
rect 2752 16292 2776 16294
rect 2832 16292 2856 16294
rect 2912 16292 2918 16294
rect 2610 16283 2918 16292
rect 2610 15260 2918 15269
rect 2610 15258 2616 15260
rect 2672 15258 2696 15260
rect 2752 15258 2776 15260
rect 2832 15258 2856 15260
rect 2912 15258 2918 15260
rect 2672 15206 2674 15258
rect 2854 15206 2856 15258
rect 2610 15204 2616 15206
rect 2672 15204 2696 15206
rect 2752 15204 2776 15206
rect 2832 15204 2856 15206
rect 2912 15204 2918 15206
rect 2610 15195 2918 15204
rect 2610 14172 2918 14181
rect 2610 14170 2616 14172
rect 2672 14170 2696 14172
rect 2752 14170 2776 14172
rect 2832 14170 2856 14172
rect 2912 14170 2918 14172
rect 2672 14118 2674 14170
rect 2854 14118 2856 14170
rect 2610 14116 2616 14118
rect 2672 14116 2696 14118
rect 2752 14116 2776 14118
rect 2832 14116 2856 14118
rect 2912 14116 2918 14118
rect 2610 14107 2918 14116
rect 2610 13084 2918 13093
rect 2610 13082 2616 13084
rect 2672 13082 2696 13084
rect 2752 13082 2776 13084
rect 2832 13082 2856 13084
rect 2912 13082 2918 13084
rect 2672 13030 2674 13082
rect 2854 13030 2856 13082
rect 2610 13028 2616 13030
rect 2672 13028 2696 13030
rect 2752 13028 2776 13030
rect 2832 13028 2856 13030
rect 2912 13028 2918 13030
rect 2610 13019 2918 13028
rect 2610 11996 2918 12005
rect 2610 11994 2616 11996
rect 2672 11994 2696 11996
rect 2752 11994 2776 11996
rect 2832 11994 2856 11996
rect 2912 11994 2918 11996
rect 2672 11942 2674 11994
rect 2854 11942 2856 11994
rect 2610 11940 2616 11942
rect 2672 11940 2696 11942
rect 2752 11940 2776 11942
rect 2832 11940 2856 11942
rect 2912 11940 2918 11942
rect 2610 11931 2918 11940
rect 2610 10908 2918 10917
rect 2610 10906 2616 10908
rect 2672 10906 2696 10908
rect 2752 10906 2776 10908
rect 2832 10906 2856 10908
rect 2912 10906 2918 10908
rect 2672 10854 2674 10906
rect 2854 10854 2856 10906
rect 2610 10852 2616 10854
rect 2672 10852 2696 10854
rect 2752 10852 2776 10854
rect 2832 10852 2856 10854
rect 2912 10852 2918 10854
rect 2610 10843 2918 10852
rect 2610 9820 2918 9829
rect 2610 9818 2616 9820
rect 2672 9818 2696 9820
rect 2752 9818 2776 9820
rect 2832 9818 2856 9820
rect 2912 9818 2918 9820
rect 2672 9766 2674 9818
rect 2854 9766 2856 9818
rect 2610 9764 2616 9766
rect 2672 9764 2696 9766
rect 2752 9764 2776 9766
rect 2832 9764 2856 9766
rect 2912 9764 2918 9766
rect 2610 9755 2918 9764
rect 2610 8732 2918 8741
rect 2610 8730 2616 8732
rect 2672 8730 2696 8732
rect 2752 8730 2776 8732
rect 2832 8730 2856 8732
rect 2912 8730 2918 8732
rect 2672 8678 2674 8730
rect 2854 8678 2856 8730
rect 2610 8676 2616 8678
rect 2672 8676 2696 8678
rect 2752 8676 2776 8678
rect 2832 8676 2856 8678
rect 2912 8676 2918 8678
rect 2610 8667 2918 8676
rect 2610 7644 2918 7653
rect 2610 7642 2616 7644
rect 2672 7642 2696 7644
rect 2752 7642 2776 7644
rect 2832 7642 2856 7644
rect 2912 7642 2918 7644
rect 2672 7590 2674 7642
rect 2854 7590 2856 7642
rect 2610 7588 2616 7590
rect 2672 7588 2696 7590
rect 2752 7588 2776 7590
rect 2832 7588 2856 7590
rect 2912 7588 2918 7590
rect 2610 7579 2918 7588
rect 2610 6556 2918 6565
rect 2610 6554 2616 6556
rect 2672 6554 2696 6556
rect 2752 6554 2776 6556
rect 2832 6554 2856 6556
rect 2912 6554 2918 6556
rect 2672 6502 2674 6554
rect 2854 6502 2856 6554
rect 2610 6500 2616 6502
rect 2672 6500 2696 6502
rect 2752 6500 2776 6502
rect 2832 6500 2856 6502
rect 2912 6500 2918 6502
rect 2610 6491 2918 6500
rect 2610 5468 2918 5477
rect 2610 5466 2616 5468
rect 2672 5466 2696 5468
rect 2752 5466 2776 5468
rect 2832 5466 2856 5468
rect 2912 5466 2918 5468
rect 2672 5414 2674 5466
rect 2854 5414 2856 5466
rect 2610 5412 2616 5414
rect 2672 5412 2696 5414
rect 2752 5412 2776 5414
rect 2832 5412 2856 5414
rect 2912 5412 2918 5414
rect 2610 5403 2918 5412
rect 2610 4380 2918 4389
rect 2610 4378 2616 4380
rect 2672 4378 2696 4380
rect 2752 4378 2776 4380
rect 2832 4378 2856 4380
rect 2912 4378 2918 4380
rect 2672 4326 2674 4378
rect 2854 4326 2856 4378
rect 2610 4324 2616 4326
rect 2672 4324 2696 4326
rect 2752 4324 2776 4326
rect 2832 4324 2856 4326
rect 2912 4324 2918 4326
rect 2610 4315 2918 4324
rect 2504 4004 2556 4010
rect 2504 3946 2556 3952
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 1676 3596 1728 3602
rect 1676 3538 1728 3544
rect 2884 3534 2912 3878
rect 3068 3670 3096 30330
rect 3160 10606 3188 45358
rect 3436 24206 3464 48146
rect 3620 40594 3648 63310
rect 3884 57452 3936 57458
rect 3884 57394 3936 57400
rect 3896 55214 3924 57394
rect 3896 55186 4016 55214
rect 3608 40588 3660 40594
rect 3608 40530 3660 40536
rect 3988 29850 4016 55186
rect 4080 52698 4108 63514
rect 5736 57526 5764 63922
rect 5724 57520 5776 57526
rect 5724 57462 5776 57468
rect 5540 57452 5592 57458
rect 5540 57394 5592 57400
rect 4988 57384 5040 57390
rect 4988 57326 5040 57332
rect 5264 57384 5316 57390
rect 5264 57326 5316 57332
rect 5356 57384 5408 57390
rect 5356 57326 5408 57332
rect 4068 52692 4120 52698
rect 4068 52634 4120 52640
rect 4344 52420 4396 52426
rect 4344 52362 4396 52368
rect 4356 52154 4384 52362
rect 4344 52148 4396 52154
rect 4344 52090 4396 52096
rect 4068 52012 4120 52018
rect 4068 51954 4120 51960
rect 4080 48210 4108 51954
rect 5000 48550 5028 57326
rect 5276 56914 5304 57326
rect 5264 56908 5316 56914
rect 5264 56850 5316 56856
rect 5264 52896 5316 52902
rect 5264 52838 5316 52844
rect 5276 52494 5304 52838
rect 5080 52488 5132 52494
rect 5080 52430 5132 52436
rect 5264 52488 5316 52494
rect 5264 52430 5316 52436
rect 4988 48544 5040 48550
rect 4988 48486 5040 48492
rect 4068 48204 4120 48210
rect 4068 48146 4120 48152
rect 4804 43648 4856 43654
rect 4804 43590 4856 43596
rect 3976 29844 4028 29850
rect 3976 29786 4028 29792
rect 3884 29708 3936 29714
rect 3884 29650 3936 29656
rect 3896 29170 3924 29650
rect 3884 29164 3936 29170
rect 3884 29106 3936 29112
rect 4816 29102 4844 43590
rect 5092 30190 5120 52430
rect 5368 45014 5396 57326
rect 5356 45008 5408 45014
rect 5356 44950 5408 44956
rect 5552 44946 5580 57394
rect 5632 52488 5684 52494
rect 5632 52430 5684 52436
rect 5540 44940 5592 44946
rect 5540 44882 5592 44888
rect 5264 44872 5316 44878
rect 5316 44820 5488 44826
rect 5264 44814 5488 44820
rect 5276 44810 5488 44814
rect 5276 44804 5500 44810
rect 5276 44798 5448 44804
rect 5448 44746 5500 44752
rect 5552 44742 5580 44882
rect 5540 44736 5592 44742
rect 5540 44678 5592 44684
rect 5264 41472 5316 41478
rect 5264 41414 5316 41420
rect 5080 30184 5132 30190
rect 5080 30126 5132 30132
rect 5276 29170 5304 41414
rect 5644 30598 5672 52430
rect 5736 44878 5764 57462
rect 6092 57384 6144 57390
rect 6092 57326 6144 57332
rect 6104 48006 6132 57326
rect 6380 53174 6408 67594
rect 6460 66632 6512 66638
rect 6460 66574 6512 66580
rect 6472 65754 6500 66574
rect 6644 66496 6696 66502
rect 6644 66438 6696 66444
rect 6460 65748 6512 65754
rect 6460 65690 6512 65696
rect 6368 53168 6420 53174
rect 6368 53110 6420 53116
rect 6184 52352 6236 52358
rect 6184 52294 6236 52300
rect 6092 48000 6144 48006
rect 6092 47942 6144 47948
rect 5724 44872 5776 44878
rect 5724 44814 5776 44820
rect 5736 38010 5764 44814
rect 5724 38004 5776 38010
rect 5724 37946 5776 37952
rect 6196 31958 6224 52294
rect 6368 38344 6420 38350
rect 6368 38286 6420 38292
rect 6380 32570 6408 38286
rect 6368 32564 6420 32570
rect 6368 32506 6420 32512
rect 6184 31952 6236 31958
rect 6184 31894 6236 31900
rect 5632 30592 5684 30598
rect 5632 30534 5684 30540
rect 6196 29646 6224 31894
rect 6472 30666 6500 65690
rect 6656 35894 6684 66438
rect 6840 55214 6868 68274
rect 6950 68028 7258 68037
rect 6950 68026 6956 68028
rect 7012 68026 7036 68028
rect 7092 68026 7116 68028
rect 7172 68026 7196 68028
rect 7252 68026 7258 68028
rect 7012 67974 7014 68026
rect 7194 67974 7196 68026
rect 6950 67972 6956 67974
rect 7012 67972 7036 67974
rect 7092 67972 7116 67974
rect 7172 67972 7196 67974
rect 7252 67972 7258 67974
rect 6950 67963 7258 67972
rect 6950 66940 7258 66949
rect 6950 66938 6956 66940
rect 7012 66938 7036 66940
rect 7092 66938 7116 66940
rect 7172 66938 7196 66940
rect 7252 66938 7258 66940
rect 7012 66886 7014 66938
rect 7194 66886 7196 66938
rect 6950 66884 6956 66886
rect 7012 66884 7036 66886
rect 7092 66884 7116 66886
rect 7172 66884 7196 66886
rect 7252 66884 7258 66886
rect 6950 66875 7258 66884
rect 6950 65852 7258 65861
rect 6950 65850 6956 65852
rect 7012 65850 7036 65852
rect 7092 65850 7116 65852
rect 7172 65850 7196 65852
rect 7252 65850 7258 65852
rect 7012 65798 7014 65850
rect 7194 65798 7196 65850
rect 6950 65796 6956 65798
rect 7012 65796 7036 65798
rect 7092 65796 7116 65798
rect 7172 65796 7196 65798
rect 7252 65796 7258 65798
rect 6950 65787 7258 65796
rect 6950 64764 7258 64773
rect 6950 64762 6956 64764
rect 7012 64762 7036 64764
rect 7092 64762 7116 64764
rect 7172 64762 7196 64764
rect 7252 64762 7258 64764
rect 7012 64710 7014 64762
rect 7194 64710 7196 64762
rect 6950 64708 6956 64710
rect 7012 64708 7036 64710
rect 7092 64708 7116 64710
rect 7172 64708 7196 64710
rect 7252 64708 7258 64710
rect 6950 64699 7258 64708
rect 6950 63676 7258 63685
rect 6950 63674 6956 63676
rect 7012 63674 7036 63676
rect 7092 63674 7116 63676
rect 7172 63674 7196 63676
rect 7252 63674 7258 63676
rect 7012 63622 7014 63674
rect 7194 63622 7196 63674
rect 6950 63620 6956 63622
rect 7012 63620 7036 63622
rect 7092 63620 7116 63622
rect 7172 63620 7196 63622
rect 7252 63620 7258 63622
rect 6950 63611 7258 63620
rect 6950 62588 7258 62597
rect 6950 62586 6956 62588
rect 7012 62586 7036 62588
rect 7092 62586 7116 62588
rect 7172 62586 7196 62588
rect 7252 62586 7258 62588
rect 7012 62534 7014 62586
rect 7194 62534 7196 62586
rect 6950 62532 6956 62534
rect 7012 62532 7036 62534
rect 7092 62532 7116 62534
rect 7172 62532 7196 62534
rect 7252 62532 7258 62534
rect 6950 62523 7258 62532
rect 6950 61500 7258 61509
rect 6950 61498 6956 61500
rect 7012 61498 7036 61500
rect 7092 61498 7116 61500
rect 7172 61498 7196 61500
rect 7252 61498 7258 61500
rect 7012 61446 7014 61498
rect 7194 61446 7196 61498
rect 6950 61444 6956 61446
rect 7012 61444 7036 61446
rect 7092 61444 7116 61446
rect 7172 61444 7196 61446
rect 7252 61444 7258 61446
rect 6950 61435 7258 61444
rect 6950 60412 7258 60421
rect 6950 60410 6956 60412
rect 7012 60410 7036 60412
rect 7092 60410 7116 60412
rect 7172 60410 7196 60412
rect 7252 60410 7258 60412
rect 7012 60358 7014 60410
rect 7194 60358 7196 60410
rect 6950 60356 6956 60358
rect 7012 60356 7036 60358
rect 7092 60356 7116 60358
rect 7172 60356 7196 60358
rect 7252 60356 7258 60358
rect 6950 60347 7258 60356
rect 6950 59324 7258 59333
rect 6950 59322 6956 59324
rect 7012 59322 7036 59324
rect 7092 59322 7116 59324
rect 7172 59322 7196 59324
rect 7252 59322 7258 59324
rect 7012 59270 7014 59322
rect 7194 59270 7196 59322
rect 6950 59268 6956 59270
rect 7012 59268 7036 59270
rect 7092 59268 7116 59270
rect 7172 59268 7196 59270
rect 7252 59268 7258 59270
rect 6950 59259 7258 59268
rect 6950 58236 7258 58245
rect 6950 58234 6956 58236
rect 7012 58234 7036 58236
rect 7092 58234 7116 58236
rect 7172 58234 7196 58236
rect 7252 58234 7258 58236
rect 7012 58182 7014 58234
rect 7194 58182 7196 58234
rect 6950 58180 6956 58182
rect 7012 58180 7036 58182
rect 7092 58180 7116 58182
rect 7172 58180 7196 58182
rect 7252 58180 7258 58182
rect 6950 58171 7258 58180
rect 6950 57148 7258 57157
rect 6950 57146 6956 57148
rect 7012 57146 7036 57148
rect 7092 57146 7116 57148
rect 7172 57146 7196 57148
rect 7252 57146 7258 57148
rect 7012 57094 7014 57146
rect 7194 57094 7196 57146
rect 6950 57092 6956 57094
rect 7012 57092 7036 57094
rect 7092 57092 7116 57094
rect 7172 57092 7196 57094
rect 7252 57092 7258 57094
rect 6950 57083 7258 57092
rect 6950 56060 7258 56069
rect 6950 56058 6956 56060
rect 7012 56058 7036 56060
rect 7092 56058 7116 56060
rect 7172 56058 7196 56060
rect 7252 56058 7258 56060
rect 7012 56006 7014 56058
rect 7194 56006 7196 56058
rect 6950 56004 6956 56006
rect 7012 56004 7036 56006
rect 7092 56004 7116 56006
rect 7172 56004 7196 56006
rect 7252 56004 7258 56006
rect 6950 55995 7258 56004
rect 6564 35866 6684 35894
rect 6748 55186 6868 55214
rect 6460 30660 6512 30666
rect 6460 30602 6512 30608
rect 6276 30592 6328 30598
rect 6276 30534 6328 30540
rect 6184 29640 6236 29646
rect 6184 29582 6236 29588
rect 6092 29572 6144 29578
rect 6092 29514 6144 29520
rect 5264 29164 5316 29170
rect 5264 29106 5316 29112
rect 4804 29096 4856 29102
rect 4804 29038 4856 29044
rect 5724 24812 5776 24818
rect 5724 24754 5776 24760
rect 3424 24200 3476 24206
rect 3424 24142 3476 24148
rect 3240 23044 3292 23050
rect 3240 22986 3292 22992
rect 3252 22778 3280 22986
rect 3240 22772 3292 22778
rect 3240 22714 3292 22720
rect 3238 22672 3294 22681
rect 3238 22607 3240 22616
rect 3292 22607 3294 22616
rect 3240 22578 3292 22584
rect 3436 20534 3464 24142
rect 5632 22976 5684 22982
rect 5632 22918 5684 22924
rect 3516 22636 3568 22642
rect 3516 22578 3568 22584
rect 3528 22098 3556 22578
rect 5644 22574 5672 22918
rect 5632 22568 5684 22574
rect 5632 22510 5684 22516
rect 3516 22092 3568 22098
rect 3516 22034 3568 22040
rect 3424 20528 3476 20534
rect 3424 20470 3476 20476
rect 3608 18624 3660 18630
rect 3608 18566 3660 18572
rect 3620 18426 3648 18566
rect 3608 18420 3660 18426
rect 3608 18362 3660 18368
rect 3884 17672 3936 17678
rect 3884 17614 3936 17620
rect 3332 17604 3384 17610
rect 3332 17546 3384 17552
rect 3344 17338 3372 17546
rect 3332 17332 3384 17338
rect 3332 17274 3384 17280
rect 3896 17270 3924 17614
rect 3884 17264 3936 17270
rect 3884 17206 3936 17212
rect 3896 16998 3924 17206
rect 5736 17134 5764 24754
rect 5724 17128 5776 17134
rect 5724 17070 5776 17076
rect 3884 16992 3936 16998
rect 3884 16934 3936 16940
rect 4528 16992 4580 16998
rect 4528 16934 4580 16940
rect 4540 16794 4568 16934
rect 4528 16788 4580 16794
rect 4528 16730 4580 16736
rect 4712 12096 4764 12102
rect 4712 12038 4764 12044
rect 3148 10600 3200 10606
rect 3148 10542 3200 10548
rect 3056 3664 3108 3670
rect 3056 3606 3108 3612
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 2610 3292 2918 3301
rect 2610 3290 2616 3292
rect 2672 3290 2696 3292
rect 2752 3290 2776 3292
rect 2832 3290 2856 3292
rect 2912 3290 2918 3292
rect 2672 3238 2674 3290
rect 2854 3238 2856 3290
rect 2610 3236 2616 3238
rect 2672 3236 2696 3238
rect 2752 3236 2776 3238
rect 2832 3236 2856 3238
rect 2912 3236 2918 3238
rect 2610 3227 2918 3236
rect 4724 3194 4752 12038
rect 6104 5030 6132 29514
rect 6184 22500 6236 22506
rect 6184 22442 6236 22448
rect 6196 17202 6224 22442
rect 6184 17196 6236 17202
rect 6184 17138 6236 17144
rect 6092 5024 6144 5030
rect 6092 4966 6144 4972
rect 6288 4622 6316 30534
rect 6460 29504 6512 29510
rect 6460 29446 6512 29452
rect 6472 29102 6500 29446
rect 6460 29096 6512 29102
rect 6460 29038 6512 29044
rect 6472 17270 6500 29038
rect 6460 17264 6512 17270
rect 6460 17206 6512 17212
rect 6472 6914 6500 17206
rect 6564 11082 6592 35866
rect 6748 24818 6776 55186
rect 6950 54972 7258 54981
rect 6950 54970 6956 54972
rect 7012 54970 7036 54972
rect 7092 54970 7116 54972
rect 7172 54970 7196 54972
rect 7252 54970 7258 54972
rect 7012 54918 7014 54970
rect 7194 54918 7196 54970
rect 6950 54916 6956 54918
rect 7012 54916 7036 54918
rect 7092 54916 7116 54918
rect 7172 54916 7196 54918
rect 7252 54916 7258 54918
rect 6950 54907 7258 54916
rect 6950 53884 7258 53893
rect 6950 53882 6956 53884
rect 7012 53882 7036 53884
rect 7092 53882 7116 53884
rect 7172 53882 7196 53884
rect 7252 53882 7258 53884
rect 7012 53830 7014 53882
rect 7194 53830 7196 53882
rect 6950 53828 6956 53830
rect 7012 53828 7036 53830
rect 7092 53828 7116 53830
rect 7172 53828 7196 53830
rect 7252 53828 7258 53830
rect 6950 53819 7258 53828
rect 6950 52796 7258 52805
rect 6950 52794 6956 52796
rect 7012 52794 7036 52796
rect 7092 52794 7116 52796
rect 7172 52794 7196 52796
rect 7252 52794 7258 52796
rect 7012 52742 7014 52794
rect 7194 52742 7196 52794
rect 6950 52740 6956 52742
rect 7012 52740 7036 52742
rect 7092 52740 7116 52742
rect 7172 52740 7196 52742
rect 7252 52740 7258 52742
rect 6950 52731 7258 52740
rect 6950 51708 7258 51717
rect 6950 51706 6956 51708
rect 7012 51706 7036 51708
rect 7092 51706 7116 51708
rect 7172 51706 7196 51708
rect 7252 51706 7258 51708
rect 7012 51654 7014 51706
rect 7194 51654 7196 51706
rect 6950 51652 6956 51654
rect 7012 51652 7036 51654
rect 7092 51652 7116 51654
rect 7172 51652 7196 51654
rect 7252 51652 7258 51654
rect 6950 51643 7258 51652
rect 6950 50620 7258 50629
rect 6950 50618 6956 50620
rect 7012 50618 7036 50620
rect 7092 50618 7116 50620
rect 7172 50618 7196 50620
rect 7252 50618 7258 50620
rect 7012 50566 7014 50618
rect 7194 50566 7196 50618
rect 6950 50564 6956 50566
rect 7012 50564 7036 50566
rect 7092 50564 7116 50566
rect 7172 50564 7196 50566
rect 7252 50564 7258 50566
rect 6950 50555 7258 50564
rect 6950 49532 7258 49541
rect 6950 49530 6956 49532
rect 7012 49530 7036 49532
rect 7092 49530 7116 49532
rect 7172 49530 7196 49532
rect 7252 49530 7258 49532
rect 7012 49478 7014 49530
rect 7194 49478 7196 49530
rect 6950 49476 6956 49478
rect 7012 49476 7036 49478
rect 7092 49476 7116 49478
rect 7172 49476 7196 49478
rect 7252 49476 7258 49478
rect 6950 49467 7258 49476
rect 6950 48444 7258 48453
rect 6950 48442 6956 48444
rect 7012 48442 7036 48444
rect 7092 48442 7116 48444
rect 7172 48442 7196 48444
rect 7252 48442 7258 48444
rect 7012 48390 7014 48442
rect 7194 48390 7196 48442
rect 6950 48388 6956 48390
rect 7012 48388 7036 48390
rect 7092 48388 7116 48390
rect 7172 48388 7196 48390
rect 7252 48388 7258 48390
rect 6950 48379 7258 48388
rect 6828 48000 6880 48006
rect 6828 47942 6880 47948
rect 6840 32434 6868 47942
rect 6950 47356 7258 47365
rect 6950 47354 6956 47356
rect 7012 47354 7036 47356
rect 7092 47354 7116 47356
rect 7172 47354 7196 47356
rect 7252 47354 7258 47356
rect 7012 47302 7014 47354
rect 7194 47302 7196 47354
rect 6950 47300 6956 47302
rect 7012 47300 7036 47302
rect 7092 47300 7116 47302
rect 7172 47300 7196 47302
rect 7252 47300 7258 47302
rect 6950 47291 7258 47300
rect 6950 46268 7258 46277
rect 6950 46266 6956 46268
rect 7012 46266 7036 46268
rect 7092 46266 7116 46268
rect 7172 46266 7196 46268
rect 7252 46266 7258 46268
rect 7012 46214 7014 46266
rect 7194 46214 7196 46266
rect 6950 46212 6956 46214
rect 7012 46212 7036 46214
rect 7092 46212 7116 46214
rect 7172 46212 7196 46214
rect 7252 46212 7258 46214
rect 6950 46203 7258 46212
rect 6950 45180 7258 45189
rect 6950 45178 6956 45180
rect 7012 45178 7036 45180
rect 7092 45178 7116 45180
rect 7172 45178 7196 45180
rect 7252 45178 7258 45180
rect 7012 45126 7014 45178
rect 7194 45126 7196 45178
rect 6950 45124 6956 45126
rect 7012 45124 7036 45126
rect 7092 45124 7116 45126
rect 7172 45124 7196 45126
rect 7252 45124 7258 45126
rect 6950 45115 7258 45124
rect 6950 44092 7258 44101
rect 6950 44090 6956 44092
rect 7012 44090 7036 44092
rect 7092 44090 7116 44092
rect 7172 44090 7196 44092
rect 7252 44090 7258 44092
rect 7012 44038 7014 44090
rect 7194 44038 7196 44090
rect 6950 44036 6956 44038
rect 7012 44036 7036 44038
rect 7092 44036 7116 44038
rect 7172 44036 7196 44038
rect 7252 44036 7258 44038
rect 6950 44027 7258 44036
rect 6950 43004 7258 43013
rect 6950 43002 6956 43004
rect 7012 43002 7036 43004
rect 7092 43002 7116 43004
rect 7172 43002 7196 43004
rect 7252 43002 7258 43004
rect 7012 42950 7014 43002
rect 7194 42950 7196 43002
rect 6950 42948 6956 42950
rect 7012 42948 7036 42950
rect 7092 42948 7116 42950
rect 7172 42948 7196 42950
rect 7252 42948 7258 42950
rect 6950 42939 7258 42948
rect 6950 41916 7258 41925
rect 6950 41914 6956 41916
rect 7012 41914 7036 41916
rect 7092 41914 7116 41916
rect 7172 41914 7196 41916
rect 7252 41914 7258 41916
rect 7012 41862 7014 41914
rect 7194 41862 7196 41914
rect 6950 41860 6956 41862
rect 7012 41860 7036 41862
rect 7092 41860 7116 41862
rect 7172 41860 7196 41862
rect 7252 41860 7258 41862
rect 6950 41851 7258 41860
rect 6950 40828 7258 40837
rect 6950 40826 6956 40828
rect 7012 40826 7036 40828
rect 7092 40826 7116 40828
rect 7172 40826 7196 40828
rect 7252 40826 7258 40828
rect 7012 40774 7014 40826
rect 7194 40774 7196 40826
rect 6950 40772 6956 40774
rect 7012 40772 7036 40774
rect 7092 40772 7116 40774
rect 7172 40772 7196 40774
rect 7252 40772 7258 40774
rect 6950 40763 7258 40772
rect 6950 39740 7258 39749
rect 6950 39738 6956 39740
rect 7012 39738 7036 39740
rect 7092 39738 7116 39740
rect 7172 39738 7196 39740
rect 7252 39738 7258 39740
rect 7012 39686 7014 39738
rect 7194 39686 7196 39738
rect 6950 39684 6956 39686
rect 7012 39684 7036 39686
rect 7092 39684 7116 39686
rect 7172 39684 7196 39686
rect 7252 39684 7258 39686
rect 6950 39675 7258 39684
rect 6950 38652 7258 38661
rect 6950 38650 6956 38652
rect 7012 38650 7036 38652
rect 7092 38650 7116 38652
rect 7172 38650 7196 38652
rect 7252 38650 7258 38652
rect 7012 38598 7014 38650
rect 7194 38598 7196 38650
rect 6950 38596 6956 38598
rect 7012 38596 7036 38598
rect 7092 38596 7116 38598
rect 7172 38596 7196 38598
rect 7252 38596 7258 38598
rect 6950 38587 7258 38596
rect 6950 37564 7258 37573
rect 6950 37562 6956 37564
rect 7012 37562 7036 37564
rect 7092 37562 7116 37564
rect 7172 37562 7196 37564
rect 7252 37562 7258 37564
rect 7012 37510 7014 37562
rect 7194 37510 7196 37562
rect 6950 37508 6956 37510
rect 7012 37508 7036 37510
rect 7092 37508 7116 37510
rect 7172 37508 7196 37510
rect 7252 37508 7258 37510
rect 6950 37499 7258 37508
rect 6950 36476 7258 36485
rect 6950 36474 6956 36476
rect 7012 36474 7036 36476
rect 7092 36474 7116 36476
rect 7172 36474 7196 36476
rect 7252 36474 7258 36476
rect 7012 36422 7014 36474
rect 7194 36422 7196 36474
rect 6950 36420 6956 36422
rect 7012 36420 7036 36422
rect 7092 36420 7116 36422
rect 7172 36420 7196 36422
rect 7252 36420 7258 36422
rect 6950 36411 7258 36420
rect 6950 35388 7258 35397
rect 6950 35386 6956 35388
rect 7012 35386 7036 35388
rect 7092 35386 7116 35388
rect 7172 35386 7196 35388
rect 7252 35386 7258 35388
rect 7012 35334 7014 35386
rect 7194 35334 7196 35386
rect 6950 35332 6956 35334
rect 7012 35332 7036 35334
rect 7092 35332 7116 35334
rect 7172 35332 7196 35334
rect 7252 35332 7258 35334
rect 6950 35323 7258 35332
rect 6950 34300 7258 34309
rect 6950 34298 6956 34300
rect 7012 34298 7036 34300
rect 7092 34298 7116 34300
rect 7172 34298 7196 34300
rect 7252 34298 7258 34300
rect 7012 34246 7014 34298
rect 7194 34246 7196 34298
rect 6950 34244 6956 34246
rect 7012 34244 7036 34246
rect 7092 34244 7116 34246
rect 7172 34244 7196 34246
rect 7252 34244 7258 34246
rect 6950 34235 7258 34244
rect 6950 33212 7258 33221
rect 6950 33210 6956 33212
rect 7012 33210 7036 33212
rect 7092 33210 7116 33212
rect 7172 33210 7196 33212
rect 7252 33210 7258 33212
rect 7012 33158 7014 33210
rect 7194 33158 7196 33210
rect 6950 33156 6956 33158
rect 7012 33156 7036 33158
rect 7092 33156 7116 33158
rect 7172 33156 7196 33158
rect 7252 33156 7258 33158
rect 6950 33147 7258 33156
rect 6828 32428 6880 32434
rect 6828 32370 6880 32376
rect 6736 24812 6788 24818
rect 6736 24754 6788 24760
rect 6748 24614 6776 24754
rect 6736 24608 6788 24614
rect 6736 24550 6788 24556
rect 6840 22778 6868 32370
rect 6950 32124 7258 32133
rect 6950 32122 6956 32124
rect 7012 32122 7036 32124
rect 7092 32122 7116 32124
rect 7172 32122 7196 32124
rect 7252 32122 7258 32124
rect 7012 32070 7014 32122
rect 7194 32070 7196 32122
rect 6950 32068 6956 32070
rect 7012 32068 7036 32070
rect 7092 32068 7116 32070
rect 7172 32068 7196 32070
rect 7252 32068 7258 32070
rect 6950 32059 7258 32068
rect 6950 31036 7258 31045
rect 6950 31034 6956 31036
rect 7012 31034 7036 31036
rect 7092 31034 7116 31036
rect 7172 31034 7196 31036
rect 7252 31034 7258 31036
rect 7012 30982 7014 31034
rect 7194 30982 7196 31034
rect 6950 30980 6956 30982
rect 7012 30980 7036 30982
rect 7092 30980 7116 30982
rect 7172 30980 7196 30982
rect 7252 30980 7258 30982
rect 6950 30971 7258 30980
rect 6950 29948 7258 29957
rect 6950 29946 6956 29948
rect 7012 29946 7036 29948
rect 7092 29946 7116 29948
rect 7172 29946 7196 29948
rect 7252 29946 7258 29948
rect 7012 29894 7014 29946
rect 7194 29894 7196 29946
rect 6950 29892 6956 29894
rect 7012 29892 7036 29894
rect 7092 29892 7116 29894
rect 7172 29892 7196 29894
rect 7252 29892 7258 29894
rect 6950 29883 7258 29892
rect 6950 28860 7258 28869
rect 6950 28858 6956 28860
rect 7012 28858 7036 28860
rect 7092 28858 7116 28860
rect 7172 28858 7196 28860
rect 7252 28858 7258 28860
rect 7012 28806 7014 28858
rect 7194 28806 7196 28858
rect 6950 28804 6956 28806
rect 7012 28804 7036 28806
rect 7092 28804 7116 28806
rect 7172 28804 7196 28806
rect 7252 28804 7258 28806
rect 6950 28795 7258 28804
rect 6950 27772 7258 27781
rect 6950 27770 6956 27772
rect 7012 27770 7036 27772
rect 7092 27770 7116 27772
rect 7172 27770 7196 27772
rect 7252 27770 7258 27772
rect 7012 27718 7014 27770
rect 7194 27718 7196 27770
rect 6950 27716 6956 27718
rect 7012 27716 7036 27718
rect 7092 27716 7116 27718
rect 7172 27716 7196 27718
rect 7252 27716 7258 27718
rect 6950 27707 7258 27716
rect 6950 26684 7258 26693
rect 6950 26682 6956 26684
rect 7012 26682 7036 26684
rect 7092 26682 7116 26684
rect 7172 26682 7196 26684
rect 7252 26682 7258 26684
rect 7012 26630 7014 26682
rect 7194 26630 7196 26682
rect 6950 26628 6956 26630
rect 7012 26628 7036 26630
rect 7092 26628 7116 26630
rect 7172 26628 7196 26630
rect 7252 26628 7258 26630
rect 6950 26619 7258 26628
rect 6950 25596 7258 25605
rect 6950 25594 6956 25596
rect 7012 25594 7036 25596
rect 7092 25594 7116 25596
rect 7172 25594 7196 25596
rect 7252 25594 7258 25596
rect 7012 25542 7014 25594
rect 7194 25542 7196 25594
rect 6950 25540 6956 25542
rect 7012 25540 7036 25542
rect 7092 25540 7116 25542
rect 7172 25540 7196 25542
rect 7252 25540 7258 25542
rect 6950 25531 7258 25540
rect 6950 24508 7258 24517
rect 6950 24506 6956 24508
rect 7012 24506 7036 24508
rect 7092 24506 7116 24508
rect 7172 24506 7196 24508
rect 7252 24506 7258 24508
rect 7012 24454 7014 24506
rect 7194 24454 7196 24506
rect 6950 24452 6956 24454
rect 7012 24452 7036 24454
rect 7092 24452 7116 24454
rect 7172 24452 7196 24454
rect 7252 24452 7258 24454
rect 6950 24443 7258 24452
rect 6950 23420 7258 23429
rect 6950 23418 6956 23420
rect 7012 23418 7036 23420
rect 7092 23418 7116 23420
rect 7172 23418 7196 23420
rect 7252 23418 7258 23420
rect 7012 23366 7014 23418
rect 7194 23366 7196 23418
rect 6950 23364 6956 23366
rect 7012 23364 7036 23366
rect 7092 23364 7116 23366
rect 7172 23364 7196 23366
rect 7252 23364 7258 23366
rect 6950 23355 7258 23364
rect 6828 22772 6880 22778
rect 6828 22714 6880 22720
rect 6920 22772 6972 22778
rect 6920 22714 6972 22720
rect 6932 22681 6960 22714
rect 7300 22710 7328 68274
rect 9036 68128 9088 68134
rect 9036 68070 9088 68076
rect 7472 67720 7524 67726
rect 7472 67662 7524 67668
rect 7484 59022 7512 67662
rect 7610 67484 7918 67493
rect 7610 67482 7616 67484
rect 7672 67482 7696 67484
rect 7752 67482 7776 67484
rect 7832 67482 7856 67484
rect 7912 67482 7918 67484
rect 7672 67430 7674 67482
rect 7854 67430 7856 67482
rect 7610 67428 7616 67430
rect 7672 67428 7696 67430
rect 7752 67428 7776 67430
rect 7832 67428 7856 67430
rect 7912 67428 7918 67430
rect 7610 67419 7918 67428
rect 7610 66396 7918 66405
rect 7610 66394 7616 66396
rect 7672 66394 7696 66396
rect 7752 66394 7776 66396
rect 7832 66394 7856 66396
rect 7912 66394 7918 66396
rect 7672 66342 7674 66394
rect 7854 66342 7856 66394
rect 7610 66340 7616 66342
rect 7672 66340 7696 66342
rect 7752 66340 7776 66342
rect 7832 66340 7856 66342
rect 7912 66340 7918 66342
rect 7610 66331 7918 66340
rect 7610 65308 7918 65317
rect 7610 65306 7616 65308
rect 7672 65306 7696 65308
rect 7752 65306 7776 65308
rect 7832 65306 7856 65308
rect 7912 65306 7918 65308
rect 7672 65254 7674 65306
rect 7854 65254 7856 65306
rect 7610 65252 7616 65254
rect 7672 65252 7696 65254
rect 7752 65252 7776 65254
rect 7832 65252 7856 65254
rect 7912 65252 7918 65254
rect 7610 65243 7918 65252
rect 7610 64220 7918 64229
rect 7610 64218 7616 64220
rect 7672 64218 7696 64220
rect 7752 64218 7776 64220
rect 7832 64218 7856 64220
rect 7912 64218 7918 64220
rect 7672 64166 7674 64218
rect 7854 64166 7856 64218
rect 7610 64164 7616 64166
rect 7672 64164 7696 64166
rect 7752 64164 7776 64166
rect 7832 64164 7856 64166
rect 7912 64164 7918 64166
rect 7610 64155 7918 64164
rect 7610 63132 7918 63141
rect 7610 63130 7616 63132
rect 7672 63130 7696 63132
rect 7752 63130 7776 63132
rect 7832 63130 7856 63132
rect 7912 63130 7918 63132
rect 7672 63078 7674 63130
rect 7854 63078 7856 63130
rect 7610 63076 7616 63078
rect 7672 63076 7696 63078
rect 7752 63076 7776 63078
rect 7832 63076 7856 63078
rect 7912 63076 7918 63078
rect 7610 63067 7918 63076
rect 7610 62044 7918 62053
rect 7610 62042 7616 62044
rect 7672 62042 7696 62044
rect 7752 62042 7776 62044
rect 7832 62042 7856 62044
rect 7912 62042 7918 62044
rect 7672 61990 7674 62042
rect 7854 61990 7856 62042
rect 7610 61988 7616 61990
rect 7672 61988 7696 61990
rect 7752 61988 7776 61990
rect 7832 61988 7856 61990
rect 7912 61988 7918 61990
rect 7610 61979 7918 61988
rect 7610 60956 7918 60965
rect 7610 60954 7616 60956
rect 7672 60954 7696 60956
rect 7752 60954 7776 60956
rect 7832 60954 7856 60956
rect 7912 60954 7918 60956
rect 7672 60902 7674 60954
rect 7854 60902 7856 60954
rect 7610 60900 7616 60902
rect 7672 60900 7696 60902
rect 7752 60900 7776 60902
rect 7832 60900 7856 60902
rect 7912 60900 7918 60902
rect 7610 60891 7918 60900
rect 7610 59868 7918 59877
rect 7610 59866 7616 59868
rect 7672 59866 7696 59868
rect 7752 59866 7776 59868
rect 7832 59866 7856 59868
rect 7912 59866 7918 59868
rect 7672 59814 7674 59866
rect 7854 59814 7856 59866
rect 7610 59812 7616 59814
rect 7672 59812 7696 59814
rect 7752 59812 7776 59814
rect 7832 59812 7856 59814
rect 7912 59812 7918 59814
rect 7610 59803 7918 59812
rect 7472 59016 7524 59022
rect 7472 58958 7524 58964
rect 8024 58880 8076 58886
rect 8024 58822 8076 58828
rect 7610 58780 7918 58789
rect 7610 58778 7616 58780
rect 7672 58778 7696 58780
rect 7752 58778 7776 58780
rect 7832 58778 7856 58780
rect 7912 58778 7918 58780
rect 7672 58726 7674 58778
rect 7854 58726 7856 58778
rect 7610 58724 7616 58726
rect 7672 58724 7696 58726
rect 7752 58724 7776 58726
rect 7832 58724 7856 58726
rect 7912 58724 7918 58726
rect 7610 58715 7918 58724
rect 7610 57692 7918 57701
rect 7610 57690 7616 57692
rect 7672 57690 7696 57692
rect 7752 57690 7776 57692
rect 7832 57690 7856 57692
rect 7912 57690 7918 57692
rect 7672 57638 7674 57690
rect 7854 57638 7856 57690
rect 7610 57636 7616 57638
rect 7672 57636 7696 57638
rect 7752 57636 7776 57638
rect 7832 57636 7856 57638
rect 7912 57636 7918 57638
rect 7610 57627 7918 57636
rect 7380 56840 7432 56846
rect 7380 56782 7432 56788
rect 7392 55214 7420 56782
rect 7610 56604 7918 56613
rect 7610 56602 7616 56604
rect 7672 56602 7696 56604
rect 7752 56602 7776 56604
rect 7832 56602 7856 56604
rect 7912 56602 7918 56604
rect 7672 56550 7674 56602
rect 7854 56550 7856 56602
rect 7610 56548 7616 56550
rect 7672 56548 7696 56550
rect 7752 56548 7776 56550
rect 7832 56548 7856 56550
rect 7912 56548 7918 56550
rect 7610 56539 7918 56548
rect 7610 55516 7918 55525
rect 7610 55514 7616 55516
rect 7672 55514 7696 55516
rect 7752 55514 7776 55516
rect 7832 55514 7856 55516
rect 7912 55514 7918 55516
rect 7672 55462 7674 55514
rect 7854 55462 7856 55514
rect 7610 55460 7616 55462
rect 7672 55460 7696 55462
rect 7752 55460 7776 55462
rect 7832 55460 7856 55462
rect 7912 55460 7918 55462
rect 7610 55451 7918 55460
rect 7392 55186 7512 55214
rect 7380 41064 7432 41070
rect 7380 41006 7432 41012
rect 7392 40662 7420 41006
rect 7484 40934 7512 55186
rect 7610 54428 7918 54437
rect 7610 54426 7616 54428
rect 7672 54426 7696 54428
rect 7752 54426 7776 54428
rect 7832 54426 7856 54428
rect 7912 54426 7918 54428
rect 7672 54374 7674 54426
rect 7854 54374 7856 54426
rect 7610 54372 7616 54374
rect 7672 54372 7696 54374
rect 7752 54372 7776 54374
rect 7832 54372 7856 54374
rect 7912 54372 7918 54374
rect 7610 54363 7918 54372
rect 7610 53340 7918 53349
rect 7610 53338 7616 53340
rect 7672 53338 7696 53340
rect 7752 53338 7776 53340
rect 7832 53338 7856 53340
rect 7912 53338 7918 53340
rect 7672 53286 7674 53338
rect 7854 53286 7856 53338
rect 7610 53284 7616 53286
rect 7672 53284 7696 53286
rect 7752 53284 7776 53286
rect 7832 53284 7856 53286
rect 7912 53284 7918 53286
rect 7610 53275 7918 53284
rect 7610 52252 7918 52261
rect 7610 52250 7616 52252
rect 7672 52250 7696 52252
rect 7752 52250 7776 52252
rect 7832 52250 7856 52252
rect 7912 52250 7918 52252
rect 7672 52198 7674 52250
rect 7854 52198 7856 52250
rect 7610 52196 7616 52198
rect 7672 52196 7696 52198
rect 7752 52196 7776 52198
rect 7832 52196 7856 52198
rect 7912 52196 7918 52198
rect 7610 52187 7918 52196
rect 7610 51164 7918 51173
rect 7610 51162 7616 51164
rect 7672 51162 7696 51164
rect 7752 51162 7776 51164
rect 7832 51162 7856 51164
rect 7912 51162 7918 51164
rect 7672 51110 7674 51162
rect 7854 51110 7856 51162
rect 7610 51108 7616 51110
rect 7672 51108 7696 51110
rect 7752 51108 7776 51110
rect 7832 51108 7856 51110
rect 7912 51108 7918 51110
rect 7610 51099 7918 51108
rect 7610 50076 7918 50085
rect 7610 50074 7616 50076
rect 7672 50074 7696 50076
rect 7752 50074 7776 50076
rect 7832 50074 7856 50076
rect 7912 50074 7918 50076
rect 7672 50022 7674 50074
rect 7854 50022 7856 50074
rect 7610 50020 7616 50022
rect 7672 50020 7696 50022
rect 7752 50020 7776 50022
rect 7832 50020 7856 50022
rect 7912 50020 7918 50022
rect 7610 50011 7918 50020
rect 7610 48988 7918 48997
rect 7610 48986 7616 48988
rect 7672 48986 7696 48988
rect 7752 48986 7776 48988
rect 7832 48986 7856 48988
rect 7912 48986 7918 48988
rect 7672 48934 7674 48986
rect 7854 48934 7856 48986
rect 7610 48932 7616 48934
rect 7672 48932 7696 48934
rect 7752 48932 7776 48934
rect 7832 48932 7856 48934
rect 7912 48932 7918 48934
rect 7610 48923 7918 48932
rect 7610 47900 7918 47909
rect 7610 47898 7616 47900
rect 7672 47898 7696 47900
rect 7752 47898 7776 47900
rect 7832 47898 7856 47900
rect 7912 47898 7918 47900
rect 7672 47846 7674 47898
rect 7854 47846 7856 47898
rect 7610 47844 7616 47846
rect 7672 47844 7696 47846
rect 7752 47844 7776 47846
rect 7832 47844 7856 47846
rect 7912 47844 7918 47846
rect 7610 47835 7918 47844
rect 7610 46812 7918 46821
rect 7610 46810 7616 46812
rect 7672 46810 7696 46812
rect 7752 46810 7776 46812
rect 7832 46810 7856 46812
rect 7912 46810 7918 46812
rect 7672 46758 7674 46810
rect 7854 46758 7856 46810
rect 7610 46756 7616 46758
rect 7672 46756 7696 46758
rect 7752 46756 7776 46758
rect 7832 46756 7856 46758
rect 7912 46756 7918 46758
rect 7610 46747 7918 46756
rect 7610 45724 7918 45733
rect 7610 45722 7616 45724
rect 7672 45722 7696 45724
rect 7752 45722 7776 45724
rect 7832 45722 7856 45724
rect 7912 45722 7918 45724
rect 7672 45670 7674 45722
rect 7854 45670 7856 45722
rect 7610 45668 7616 45670
rect 7672 45668 7696 45670
rect 7752 45668 7776 45670
rect 7832 45668 7856 45670
rect 7912 45668 7918 45670
rect 7610 45659 7918 45668
rect 7610 44636 7918 44645
rect 7610 44634 7616 44636
rect 7672 44634 7696 44636
rect 7752 44634 7776 44636
rect 7832 44634 7856 44636
rect 7912 44634 7918 44636
rect 7672 44582 7674 44634
rect 7854 44582 7856 44634
rect 7610 44580 7616 44582
rect 7672 44580 7696 44582
rect 7752 44580 7776 44582
rect 7832 44580 7856 44582
rect 7912 44580 7918 44582
rect 7610 44571 7918 44580
rect 7610 43548 7918 43557
rect 7610 43546 7616 43548
rect 7672 43546 7696 43548
rect 7752 43546 7776 43548
rect 7832 43546 7856 43548
rect 7912 43546 7918 43548
rect 7672 43494 7674 43546
rect 7854 43494 7856 43546
rect 7610 43492 7616 43494
rect 7672 43492 7696 43494
rect 7752 43492 7776 43494
rect 7832 43492 7856 43494
rect 7912 43492 7918 43494
rect 7610 43483 7918 43492
rect 7610 42460 7918 42469
rect 7610 42458 7616 42460
rect 7672 42458 7696 42460
rect 7752 42458 7776 42460
rect 7832 42458 7856 42460
rect 7912 42458 7918 42460
rect 7672 42406 7674 42458
rect 7854 42406 7856 42458
rect 7610 42404 7616 42406
rect 7672 42404 7696 42406
rect 7752 42404 7776 42406
rect 7832 42404 7856 42406
rect 7912 42404 7918 42406
rect 7610 42395 7918 42404
rect 7610 41372 7918 41381
rect 7610 41370 7616 41372
rect 7672 41370 7696 41372
rect 7752 41370 7776 41372
rect 7832 41370 7856 41372
rect 7912 41370 7918 41372
rect 7672 41318 7674 41370
rect 7854 41318 7856 41370
rect 7610 41316 7616 41318
rect 7672 41316 7696 41318
rect 7752 41316 7776 41318
rect 7832 41316 7856 41318
rect 7912 41316 7918 41318
rect 7610 41307 7918 41316
rect 7564 41132 7616 41138
rect 7564 41074 7616 41080
rect 7472 40928 7524 40934
rect 7472 40870 7524 40876
rect 7380 40656 7432 40662
rect 7380 40598 7432 40604
rect 7576 40474 7604 41074
rect 7484 40446 7604 40474
rect 7380 31748 7432 31754
rect 7380 31690 7432 31696
rect 7392 31346 7420 31690
rect 7380 31340 7432 31346
rect 7380 31282 7432 31288
rect 7380 29164 7432 29170
rect 7380 29106 7432 29112
rect 7288 22704 7340 22710
rect 6918 22672 6974 22681
rect 7288 22646 7340 22652
rect 6918 22607 6974 22616
rect 6950 22332 7258 22341
rect 6950 22330 6956 22332
rect 7012 22330 7036 22332
rect 7092 22330 7116 22332
rect 7172 22330 7196 22332
rect 7252 22330 7258 22332
rect 7012 22278 7014 22330
rect 7194 22278 7196 22330
rect 6950 22276 6956 22278
rect 7012 22276 7036 22278
rect 7092 22276 7116 22278
rect 7172 22276 7196 22278
rect 7252 22276 7258 22278
rect 6950 22267 7258 22276
rect 7300 22234 7328 22646
rect 6920 22228 6972 22234
rect 6920 22170 6972 22176
rect 7288 22228 7340 22234
rect 7288 22170 7340 22176
rect 6932 21350 6960 22170
rect 7288 22092 7340 22098
rect 7288 22034 7340 22040
rect 6920 21344 6972 21350
rect 6920 21286 6972 21292
rect 6950 21244 7258 21253
rect 6950 21242 6956 21244
rect 7012 21242 7036 21244
rect 7092 21242 7116 21244
rect 7172 21242 7196 21244
rect 7252 21242 7258 21244
rect 7012 21190 7014 21242
rect 7194 21190 7196 21242
rect 6950 21188 6956 21190
rect 7012 21188 7036 21190
rect 7092 21188 7116 21190
rect 7172 21188 7196 21190
rect 7252 21188 7258 21190
rect 6950 21179 7258 21188
rect 6644 20392 6696 20398
rect 6644 20334 6696 20340
rect 6656 19514 6684 20334
rect 6950 20156 7258 20165
rect 6950 20154 6956 20156
rect 7012 20154 7036 20156
rect 7092 20154 7116 20156
rect 7172 20154 7196 20156
rect 7252 20154 7258 20156
rect 7012 20102 7014 20154
rect 7194 20102 7196 20154
rect 6950 20100 6956 20102
rect 7012 20100 7036 20102
rect 7092 20100 7116 20102
rect 7172 20100 7196 20102
rect 7252 20100 7258 20102
rect 6950 20091 7258 20100
rect 6644 19508 6696 19514
rect 6644 19450 6696 19456
rect 6656 19378 6684 19450
rect 6644 19372 6696 19378
rect 6644 19314 6696 19320
rect 6950 19068 7258 19077
rect 6950 19066 6956 19068
rect 7012 19066 7036 19068
rect 7092 19066 7116 19068
rect 7172 19066 7196 19068
rect 7252 19066 7258 19068
rect 7012 19014 7014 19066
rect 7194 19014 7196 19066
rect 6950 19012 6956 19014
rect 7012 19012 7036 19014
rect 7092 19012 7116 19014
rect 7172 19012 7196 19014
rect 7252 19012 7258 19014
rect 6950 19003 7258 19012
rect 6950 17980 7258 17989
rect 6950 17978 6956 17980
rect 7012 17978 7036 17980
rect 7092 17978 7116 17980
rect 7172 17978 7196 17980
rect 7252 17978 7258 17980
rect 7012 17926 7014 17978
rect 7194 17926 7196 17978
rect 6950 17924 6956 17926
rect 7012 17924 7036 17926
rect 7092 17924 7116 17926
rect 7172 17924 7196 17926
rect 7252 17924 7258 17926
rect 6950 17915 7258 17924
rect 6950 16892 7258 16901
rect 6950 16890 6956 16892
rect 7012 16890 7036 16892
rect 7092 16890 7116 16892
rect 7172 16890 7196 16892
rect 7252 16890 7258 16892
rect 7012 16838 7014 16890
rect 7194 16838 7196 16890
rect 6950 16836 6956 16838
rect 7012 16836 7036 16838
rect 7092 16836 7116 16838
rect 7172 16836 7196 16838
rect 7252 16836 7258 16838
rect 6950 16827 7258 16836
rect 6950 15804 7258 15813
rect 6950 15802 6956 15804
rect 7012 15802 7036 15804
rect 7092 15802 7116 15804
rect 7172 15802 7196 15804
rect 7252 15802 7258 15804
rect 7012 15750 7014 15802
rect 7194 15750 7196 15802
rect 6950 15748 6956 15750
rect 7012 15748 7036 15750
rect 7092 15748 7116 15750
rect 7172 15748 7196 15750
rect 7252 15748 7258 15750
rect 6950 15739 7258 15748
rect 6950 14716 7258 14725
rect 6950 14714 6956 14716
rect 7012 14714 7036 14716
rect 7092 14714 7116 14716
rect 7172 14714 7196 14716
rect 7252 14714 7258 14716
rect 7012 14662 7014 14714
rect 7194 14662 7196 14714
rect 6950 14660 6956 14662
rect 7012 14660 7036 14662
rect 7092 14660 7116 14662
rect 7172 14660 7196 14662
rect 7252 14660 7258 14662
rect 6950 14651 7258 14660
rect 6950 13628 7258 13637
rect 6950 13626 6956 13628
rect 7012 13626 7036 13628
rect 7092 13626 7116 13628
rect 7172 13626 7196 13628
rect 7252 13626 7258 13628
rect 7012 13574 7014 13626
rect 7194 13574 7196 13626
rect 6950 13572 6956 13574
rect 7012 13572 7036 13574
rect 7092 13572 7116 13574
rect 7172 13572 7196 13574
rect 7252 13572 7258 13574
rect 6950 13563 7258 13572
rect 6950 12540 7258 12549
rect 6950 12538 6956 12540
rect 7012 12538 7036 12540
rect 7092 12538 7116 12540
rect 7172 12538 7196 12540
rect 7252 12538 7258 12540
rect 7012 12486 7014 12538
rect 7194 12486 7196 12538
rect 6950 12484 6956 12486
rect 7012 12484 7036 12486
rect 7092 12484 7116 12486
rect 7172 12484 7196 12486
rect 7252 12484 7258 12486
rect 6950 12475 7258 12484
rect 6950 11452 7258 11461
rect 6950 11450 6956 11452
rect 7012 11450 7036 11452
rect 7092 11450 7116 11452
rect 7172 11450 7196 11452
rect 7252 11450 7258 11452
rect 7012 11398 7014 11450
rect 7194 11398 7196 11450
rect 6950 11396 6956 11398
rect 7012 11396 7036 11398
rect 7092 11396 7116 11398
rect 7172 11396 7196 11398
rect 7252 11396 7258 11398
rect 6950 11387 7258 11396
rect 6552 11076 6604 11082
rect 6552 11018 6604 11024
rect 6950 10364 7258 10373
rect 6950 10362 6956 10364
rect 7012 10362 7036 10364
rect 7092 10362 7116 10364
rect 7172 10362 7196 10364
rect 7252 10362 7258 10364
rect 7012 10310 7014 10362
rect 7194 10310 7196 10362
rect 6950 10308 6956 10310
rect 7012 10308 7036 10310
rect 7092 10308 7116 10310
rect 7172 10308 7196 10310
rect 7252 10308 7258 10310
rect 6950 10299 7258 10308
rect 6950 9276 7258 9285
rect 6950 9274 6956 9276
rect 7012 9274 7036 9276
rect 7092 9274 7116 9276
rect 7172 9274 7196 9276
rect 7252 9274 7258 9276
rect 7012 9222 7014 9274
rect 7194 9222 7196 9274
rect 6950 9220 6956 9222
rect 7012 9220 7036 9222
rect 7092 9220 7116 9222
rect 7172 9220 7196 9222
rect 7252 9220 7258 9222
rect 6950 9211 7258 9220
rect 6950 8188 7258 8197
rect 6950 8186 6956 8188
rect 7012 8186 7036 8188
rect 7092 8186 7116 8188
rect 7172 8186 7196 8188
rect 7252 8186 7258 8188
rect 7012 8134 7014 8186
rect 7194 8134 7196 8186
rect 6950 8132 6956 8134
rect 7012 8132 7036 8134
rect 7092 8132 7116 8134
rect 7172 8132 7196 8134
rect 7252 8132 7258 8134
rect 6950 8123 7258 8132
rect 6950 7100 7258 7109
rect 6950 7098 6956 7100
rect 7012 7098 7036 7100
rect 7092 7098 7116 7100
rect 7172 7098 7196 7100
rect 7252 7098 7258 7100
rect 7012 7046 7014 7098
rect 7194 7046 7196 7098
rect 6950 7044 6956 7046
rect 7012 7044 7036 7046
rect 7092 7044 7116 7046
rect 7172 7044 7196 7046
rect 7252 7044 7258 7046
rect 6950 7035 7258 7044
rect 6380 6886 6500 6914
rect 6276 4616 6328 4622
rect 6276 4558 6328 4564
rect 6184 4480 6236 4486
rect 6184 4422 6236 4428
rect 6196 3466 6224 4422
rect 6184 3460 6236 3466
rect 6184 3402 6236 3408
rect 6380 3398 6408 6886
rect 6950 6012 7258 6021
rect 6950 6010 6956 6012
rect 7012 6010 7036 6012
rect 7092 6010 7116 6012
rect 7172 6010 7196 6012
rect 7252 6010 7258 6012
rect 7012 5958 7014 6010
rect 7194 5958 7196 6010
rect 6950 5956 6956 5958
rect 7012 5956 7036 5958
rect 7092 5956 7116 5958
rect 7172 5956 7196 5958
rect 7252 5956 7258 5958
rect 6950 5947 7258 5956
rect 6950 4924 7258 4933
rect 6950 4922 6956 4924
rect 7012 4922 7036 4924
rect 7092 4922 7116 4924
rect 7172 4922 7196 4924
rect 7252 4922 7258 4924
rect 7012 4870 7014 4922
rect 7194 4870 7196 4922
rect 6950 4868 6956 4870
rect 7012 4868 7036 4870
rect 7092 4868 7116 4870
rect 7172 4868 7196 4870
rect 7252 4868 7258 4870
rect 6950 4859 7258 4868
rect 6950 3836 7258 3845
rect 6950 3834 6956 3836
rect 7012 3834 7036 3836
rect 7092 3834 7116 3836
rect 7172 3834 7196 3836
rect 7252 3834 7258 3836
rect 7012 3782 7014 3834
rect 7194 3782 7196 3834
rect 6950 3780 6956 3782
rect 7012 3780 7036 3782
rect 7092 3780 7116 3782
rect 7172 3780 7196 3782
rect 7252 3780 7258 3782
rect 6950 3771 7258 3780
rect 6368 3392 6420 3398
rect 6368 3334 6420 3340
rect 7012 3392 7064 3398
rect 7012 3334 7064 3340
rect 4712 3188 4764 3194
rect 4712 3130 4764 3136
rect 7024 3126 7052 3334
rect 7012 3120 7064 3126
rect 7012 3062 7064 3068
rect 7300 3058 7328 22034
rect 7392 3534 7420 29106
rect 7484 17542 7512 40446
rect 7610 40284 7918 40293
rect 7610 40282 7616 40284
rect 7672 40282 7696 40284
rect 7752 40282 7776 40284
rect 7832 40282 7856 40284
rect 7912 40282 7918 40284
rect 7672 40230 7674 40282
rect 7854 40230 7856 40282
rect 7610 40228 7616 40230
rect 7672 40228 7696 40230
rect 7752 40228 7776 40230
rect 7832 40228 7856 40230
rect 7912 40228 7918 40230
rect 7610 40219 7918 40228
rect 7610 39196 7918 39205
rect 7610 39194 7616 39196
rect 7672 39194 7696 39196
rect 7752 39194 7776 39196
rect 7832 39194 7856 39196
rect 7912 39194 7918 39196
rect 7672 39142 7674 39194
rect 7854 39142 7856 39194
rect 7610 39140 7616 39142
rect 7672 39140 7696 39142
rect 7752 39140 7776 39142
rect 7832 39140 7856 39142
rect 7912 39140 7918 39142
rect 7610 39131 7918 39140
rect 7610 38108 7918 38117
rect 7610 38106 7616 38108
rect 7672 38106 7696 38108
rect 7752 38106 7776 38108
rect 7832 38106 7856 38108
rect 7912 38106 7918 38108
rect 7672 38054 7674 38106
rect 7854 38054 7856 38106
rect 7610 38052 7616 38054
rect 7672 38052 7696 38054
rect 7752 38052 7776 38054
rect 7832 38052 7856 38054
rect 7912 38052 7918 38054
rect 7610 38043 7918 38052
rect 7610 37020 7918 37029
rect 7610 37018 7616 37020
rect 7672 37018 7696 37020
rect 7752 37018 7776 37020
rect 7832 37018 7856 37020
rect 7912 37018 7918 37020
rect 7672 36966 7674 37018
rect 7854 36966 7856 37018
rect 7610 36964 7616 36966
rect 7672 36964 7696 36966
rect 7752 36964 7776 36966
rect 7832 36964 7856 36966
rect 7912 36964 7918 36966
rect 7610 36955 7918 36964
rect 7610 35932 7918 35941
rect 7610 35930 7616 35932
rect 7672 35930 7696 35932
rect 7752 35930 7776 35932
rect 7832 35930 7856 35932
rect 7912 35930 7918 35932
rect 7672 35878 7674 35930
rect 7854 35878 7856 35930
rect 7610 35876 7616 35878
rect 7672 35876 7696 35878
rect 7752 35876 7776 35878
rect 7832 35876 7856 35878
rect 7912 35876 7918 35878
rect 7610 35867 7918 35876
rect 7610 34844 7918 34853
rect 7610 34842 7616 34844
rect 7672 34842 7696 34844
rect 7752 34842 7776 34844
rect 7832 34842 7856 34844
rect 7912 34842 7918 34844
rect 7672 34790 7674 34842
rect 7854 34790 7856 34842
rect 7610 34788 7616 34790
rect 7672 34788 7696 34790
rect 7752 34788 7776 34790
rect 7832 34788 7856 34790
rect 7912 34788 7918 34790
rect 7610 34779 7918 34788
rect 7610 33756 7918 33765
rect 7610 33754 7616 33756
rect 7672 33754 7696 33756
rect 7752 33754 7776 33756
rect 7832 33754 7856 33756
rect 7912 33754 7918 33756
rect 7672 33702 7674 33754
rect 7854 33702 7856 33754
rect 7610 33700 7616 33702
rect 7672 33700 7696 33702
rect 7752 33700 7776 33702
rect 7832 33700 7856 33702
rect 7912 33700 7918 33702
rect 7610 33691 7918 33700
rect 7610 32668 7918 32677
rect 7610 32666 7616 32668
rect 7672 32666 7696 32668
rect 7752 32666 7776 32668
rect 7832 32666 7856 32668
rect 7912 32666 7918 32668
rect 7672 32614 7674 32666
rect 7854 32614 7856 32666
rect 7610 32612 7616 32614
rect 7672 32612 7696 32614
rect 7752 32612 7776 32614
rect 7832 32612 7856 32614
rect 7912 32612 7918 32614
rect 7610 32603 7918 32612
rect 7610 31580 7918 31589
rect 7610 31578 7616 31580
rect 7672 31578 7696 31580
rect 7752 31578 7776 31580
rect 7832 31578 7856 31580
rect 7912 31578 7918 31580
rect 7672 31526 7674 31578
rect 7854 31526 7856 31578
rect 7610 31524 7616 31526
rect 7672 31524 7696 31526
rect 7752 31524 7776 31526
rect 7832 31524 7856 31526
rect 7912 31524 7918 31526
rect 7610 31515 7918 31524
rect 7610 30492 7918 30501
rect 7610 30490 7616 30492
rect 7672 30490 7696 30492
rect 7752 30490 7776 30492
rect 7832 30490 7856 30492
rect 7912 30490 7918 30492
rect 7672 30438 7674 30490
rect 7854 30438 7856 30490
rect 7610 30436 7616 30438
rect 7672 30436 7696 30438
rect 7752 30436 7776 30438
rect 7832 30436 7856 30438
rect 7912 30436 7918 30438
rect 7610 30427 7918 30436
rect 7610 29404 7918 29413
rect 7610 29402 7616 29404
rect 7672 29402 7696 29404
rect 7752 29402 7776 29404
rect 7832 29402 7856 29404
rect 7912 29402 7918 29404
rect 7672 29350 7674 29402
rect 7854 29350 7856 29402
rect 7610 29348 7616 29350
rect 7672 29348 7696 29350
rect 7752 29348 7776 29350
rect 7832 29348 7856 29350
rect 7912 29348 7918 29350
rect 7610 29339 7918 29348
rect 7610 28316 7918 28325
rect 7610 28314 7616 28316
rect 7672 28314 7696 28316
rect 7752 28314 7776 28316
rect 7832 28314 7856 28316
rect 7912 28314 7918 28316
rect 7672 28262 7674 28314
rect 7854 28262 7856 28314
rect 7610 28260 7616 28262
rect 7672 28260 7696 28262
rect 7752 28260 7776 28262
rect 7832 28260 7856 28262
rect 7912 28260 7918 28262
rect 7610 28251 7918 28260
rect 7610 27228 7918 27237
rect 7610 27226 7616 27228
rect 7672 27226 7696 27228
rect 7752 27226 7776 27228
rect 7832 27226 7856 27228
rect 7912 27226 7918 27228
rect 7672 27174 7674 27226
rect 7854 27174 7856 27226
rect 7610 27172 7616 27174
rect 7672 27172 7696 27174
rect 7752 27172 7776 27174
rect 7832 27172 7856 27174
rect 7912 27172 7918 27174
rect 7610 27163 7918 27172
rect 7610 26140 7918 26149
rect 7610 26138 7616 26140
rect 7672 26138 7696 26140
rect 7752 26138 7776 26140
rect 7832 26138 7856 26140
rect 7912 26138 7918 26140
rect 7672 26086 7674 26138
rect 7854 26086 7856 26138
rect 7610 26084 7616 26086
rect 7672 26084 7696 26086
rect 7752 26084 7776 26086
rect 7832 26084 7856 26086
rect 7912 26084 7918 26086
rect 7610 26075 7918 26084
rect 7610 25052 7918 25061
rect 7610 25050 7616 25052
rect 7672 25050 7696 25052
rect 7752 25050 7776 25052
rect 7832 25050 7856 25052
rect 7912 25050 7918 25052
rect 7672 24998 7674 25050
rect 7854 24998 7856 25050
rect 7610 24996 7616 24998
rect 7672 24996 7696 24998
rect 7752 24996 7776 24998
rect 7832 24996 7856 24998
rect 7912 24996 7918 24998
rect 7610 24987 7918 24996
rect 7610 23964 7918 23973
rect 7610 23962 7616 23964
rect 7672 23962 7696 23964
rect 7752 23962 7776 23964
rect 7832 23962 7856 23964
rect 7912 23962 7918 23964
rect 7672 23910 7674 23962
rect 7854 23910 7856 23962
rect 7610 23908 7616 23910
rect 7672 23908 7696 23910
rect 7752 23908 7776 23910
rect 7832 23908 7856 23910
rect 7912 23908 7918 23910
rect 7610 23899 7918 23908
rect 7610 22876 7918 22885
rect 7610 22874 7616 22876
rect 7672 22874 7696 22876
rect 7752 22874 7776 22876
rect 7832 22874 7856 22876
rect 7912 22874 7918 22876
rect 7672 22822 7674 22874
rect 7854 22822 7856 22874
rect 7610 22820 7616 22822
rect 7672 22820 7696 22822
rect 7752 22820 7776 22822
rect 7832 22820 7856 22822
rect 7912 22820 7918 22822
rect 7610 22811 7918 22820
rect 7610 21788 7918 21797
rect 7610 21786 7616 21788
rect 7672 21786 7696 21788
rect 7752 21786 7776 21788
rect 7832 21786 7856 21788
rect 7912 21786 7918 21788
rect 7672 21734 7674 21786
rect 7854 21734 7856 21786
rect 7610 21732 7616 21734
rect 7672 21732 7696 21734
rect 7752 21732 7776 21734
rect 7832 21732 7856 21734
rect 7912 21732 7918 21734
rect 7610 21723 7918 21732
rect 7610 20700 7918 20709
rect 7610 20698 7616 20700
rect 7672 20698 7696 20700
rect 7752 20698 7776 20700
rect 7832 20698 7856 20700
rect 7912 20698 7918 20700
rect 7672 20646 7674 20698
rect 7854 20646 7856 20698
rect 7610 20644 7616 20646
rect 7672 20644 7696 20646
rect 7752 20644 7776 20646
rect 7832 20644 7856 20646
rect 7912 20644 7918 20646
rect 7610 20635 7918 20644
rect 7610 19612 7918 19621
rect 7610 19610 7616 19612
rect 7672 19610 7696 19612
rect 7752 19610 7776 19612
rect 7832 19610 7856 19612
rect 7912 19610 7918 19612
rect 7672 19558 7674 19610
rect 7854 19558 7856 19610
rect 7610 19556 7616 19558
rect 7672 19556 7696 19558
rect 7752 19556 7776 19558
rect 7832 19556 7856 19558
rect 7912 19556 7918 19558
rect 7610 19547 7918 19556
rect 7610 18524 7918 18533
rect 7610 18522 7616 18524
rect 7672 18522 7696 18524
rect 7752 18522 7776 18524
rect 7832 18522 7856 18524
rect 7912 18522 7918 18524
rect 7672 18470 7674 18522
rect 7854 18470 7856 18522
rect 7610 18468 7616 18470
rect 7672 18468 7696 18470
rect 7752 18468 7776 18470
rect 7832 18468 7856 18470
rect 7912 18468 7918 18470
rect 7610 18459 7918 18468
rect 7472 17536 7524 17542
rect 7472 17478 7524 17484
rect 7610 17436 7918 17445
rect 7610 17434 7616 17436
rect 7672 17434 7696 17436
rect 7752 17434 7776 17436
rect 7832 17434 7856 17436
rect 7912 17434 7918 17436
rect 7672 17382 7674 17434
rect 7854 17382 7856 17434
rect 7610 17380 7616 17382
rect 7672 17380 7696 17382
rect 7752 17380 7776 17382
rect 7832 17380 7856 17382
rect 7912 17380 7918 17382
rect 7610 17371 7918 17380
rect 7610 16348 7918 16357
rect 7610 16346 7616 16348
rect 7672 16346 7696 16348
rect 7752 16346 7776 16348
rect 7832 16346 7856 16348
rect 7912 16346 7918 16348
rect 7672 16294 7674 16346
rect 7854 16294 7856 16346
rect 7610 16292 7616 16294
rect 7672 16292 7696 16294
rect 7752 16292 7776 16294
rect 7832 16292 7856 16294
rect 7912 16292 7918 16294
rect 7610 16283 7918 16292
rect 7610 15260 7918 15269
rect 7610 15258 7616 15260
rect 7672 15258 7696 15260
rect 7752 15258 7776 15260
rect 7832 15258 7856 15260
rect 7912 15258 7918 15260
rect 7672 15206 7674 15258
rect 7854 15206 7856 15258
rect 7610 15204 7616 15206
rect 7672 15204 7696 15206
rect 7752 15204 7776 15206
rect 7832 15204 7856 15206
rect 7912 15204 7918 15206
rect 7610 15195 7918 15204
rect 7610 14172 7918 14181
rect 7610 14170 7616 14172
rect 7672 14170 7696 14172
rect 7752 14170 7776 14172
rect 7832 14170 7856 14172
rect 7912 14170 7918 14172
rect 7672 14118 7674 14170
rect 7854 14118 7856 14170
rect 7610 14116 7616 14118
rect 7672 14116 7696 14118
rect 7752 14116 7776 14118
rect 7832 14116 7856 14118
rect 7912 14116 7918 14118
rect 7610 14107 7918 14116
rect 8036 14006 8064 58822
rect 8300 57588 8352 57594
rect 8300 57530 8352 57536
rect 8312 56710 8340 57530
rect 8392 56908 8444 56914
rect 8392 56850 8444 56856
rect 8300 56704 8352 56710
rect 8300 56646 8352 56652
rect 8312 50794 8340 56646
rect 8404 54194 8432 56850
rect 8392 54188 8444 54194
rect 8392 54130 8444 54136
rect 8300 50788 8352 50794
rect 8300 50730 8352 50736
rect 8404 46730 8432 54130
rect 8668 54120 8720 54126
rect 8668 54062 8720 54068
rect 8484 50788 8536 50794
rect 8484 50730 8536 50736
rect 8312 46702 8432 46730
rect 8312 45626 8340 46702
rect 8300 45620 8352 45626
rect 8300 45562 8352 45568
rect 8312 45490 8340 45562
rect 8300 45484 8352 45490
rect 8300 45426 8352 45432
rect 8496 44810 8524 50730
rect 8484 44804 8536 44810
rect 8484 44746 8536 44752
rect 8300 41132 8352 41138
rect 8300 41074 8352 41080
rect 8208 41064 8260 41070
rect 8208 41006 8260 41012
rect 8116 39364 8168 39370
rect 8116 39306 8168 39312
rect 8024 14000 8076 14006
rect 8024 13942 8076 13948
rect 7610 13084 7918 13093
rect 7610 13082 7616 13084
rect 7672 13082 7696 13084
rect 7752 13082 7776 13084
rect 7832 13082 7856 13084
rect 7912 13082 7918 13084
rect 7672 13030 7674 13082
rect 7854 13030 7856 13082
rect 7610 13028 7616 13030
rect 7672 13028 7696 13030
rect 7752 13028 7776 13030
rect 7832 13028 7856 13030
rect 7912 13028 7918 13030
rect 7610 13019 7918 13028
rect 7610 11996 7918 12005
rect 7610 11994 7616 11996
rect 7672 11994 7696 11996
rect 7752 11994 7776 11996
rect 7832 11994 7856 11996
rect 7912 11994 7918 11996
rect 7672 11942 7674 11994
rect 7854 11942 7856 11994
rect 7610 11940 7616 11942
rect 7672 11940 7696 11942
rect 7752 11940 7776 11942
rect 7832 11940 7856 11942
rect 7912 11940 7918 11942
rect 7610 11931 7918 11940
rect 7610 10908 7918 10917
rect 7610 10906 7616 10908
rect 7672 10906 7696 10908
rect 7752 10906 7776 10908
rect 7832 10906 7856 10908
rect 7912 10906 7918 10908
rect 7672 10854 7674 10906
rect 7854 10854 7856 10906
rect 7610 10852 7616 10854
rect 7672 10852 7696 10854
rect 7752 10852 7776 10854
rect 7832 10852 7856 10854
rect 7912 10852 7918 10854
rect 7610 10843 7918 10852
rect 7610 9820 7918 9829
rect 7610 9818 7616 9820
rect 7672 9818 7696 9820
rect 7752 9818 7776 9820
rect 7832 9818 7856 9820
rect 7912 9818 7918 9820
rect 7672 9766 7674 9818
rect 7854 9766 7856 9818
rect 7610 9764 7616 9766
rect 7672 9764 7696 9766
rect 7752 9764 7776 9766
rect 7832 9764 7856 9766
rect 7912 9764 7918 9766
rect 7610 9755 7918 9764
rect 7564 9648 7616 9654
rect 7562 9616 7564 9625
rect 7616 9616 7618 9625
rect 7562 9551 7618 9560
rect 7576 9178 7604 9551
rect 7564 9172 7616 9178
rect 7564 9114 7616 9120
rect 7610 8732 7918 8741
rect 7610 8730 7616 8732
rect 7672 8730 7696 8732
rect 7752 8730 7776 8732
rect 7832 8730 7856 8732
rect 7912 8730 7918 8732
rect 7672 8678 7674 8730
rect 7854 8678 7856 8730
rect 7610 8676 7616 8678
rect 7672 8676 7696 8678
rect 7752 8676 7776 8678
rect 7832 8676 7856 8678
rect 7912 8676 7918 8678
rect 7610 8667 7918 8676
rect 7610 7644 7918 7653
rect 7610 7642 7616 7644
rect 7672 7642 7696 7644
rect 7752 7642 7776 7644
rect 7832 7642 7856 7644
rect 7912 7642 7918 7644
rect 7672 7590 7674 7642
rect 7854 7590 7856 7642
rect 7610 7588 7616 7590
rect 7672 7588 7696 7590
rect 7752 7588 7776 7590
rect 7832 7588 7856 7590
rect 7912 7588 7918 7590
rect 7610 7579 7918 7588
rect 7610 6556 7918 6565
rect 7610 6554 7616 6556
rect 7672 6554 7696 6556
rect 7752 6554 7776 6556
rect 7832 6554 7856 6556
rect 7912 6554 7918 6556
rect 7672 6502 7674 6554
rect 7854 6502 7856 6554
rect 7610 6500 7616 6502
rect 7672 6500 7696 6502
rect 7752 6500 7776 6502
rect 7832 6500 7856 6502
rect 7912 6500 7918 6502
rect 7610 6491 7918 6500
rect 7610 5468 7918 5477
rect 7610 5466 7616 5468
rect 7672 5466 7696 5468
rect 7752 5466 7776 5468
rect 7832 5466 7856 5468
rect 7912 5466 7918 5468
rect 7672 5414 7674 5466
rect 7854 5414 7856 5466
rect 7610 5412 7616 5414
rect 7672 5412 7696 5414
rect 7752 5412 7776 5414
rect 7832 5412 7856 5414
rect 7912 5412 7918 5414
rect 7610 5403 7918 5412
rect 7610 4380 7918 4389
rect 7610 4378 7616 4380
rect 7672 4378 7696 4380
rect 7752 4378 7776 4380
rect 7832 4378 7856 4380
rect 7912 4378 7918 4380
rect 7672 4326 7674 4378
rect 7854 4326 7856 4378
rect 7610 4324 7616 4326
rect 7672 4324 7696 4326
rect 7752 4324 7776 4326
rect 7832 4324 7856 4326
rect 7912 4324 7918 4326
rect 7610 4315 7918 4324
rect 7380 3528 7432 3534
rect 7380 3470 7432 3476
rect 7610 3292 7918 3301
rect 7610 3290 7616 3292
rect 7672 3290 7696 3292
rect 7752 3290 7776 3292
rect 7832 3290 7856 3292
rect 7912 3290 7918 3292
rect 7672 3238 7674 3290
rect 7854 3238 7856 3290
rect 7610 3236 7616 3238
rect 7672 3236 7696 3238
rect 7752 3236 7776 3238
rect 7832 3236 7856 3238
rect 7912 3236 7918 3238
rect 7610 3227 7918 3236
rect 8128 3058 8156 39306
rect 8220 31346 8248 41006
rect 8312 36922 8340 41074
rect 8392 38888 8444 38894
rect 8392 38830 8444 38836
rect 8300 36916 8352 36922
rect 8300 36858 8352 36864
rect 8404 36854 8432 38830
rect 8392 36848 8444 36854
rect 8392 36790 8444 36796
rect 8496 36174 8524 44746
rect 8484 36168 8536 36174
rect 8484 36110 8536 36116
rect 8680 34542 8708 54062
rect 9048 49094 9076 68070
rect 9140 66162 9168 68342
rect 9128 66156 9180 66162
rect 9128 66098 9180 66104
rect 9036 49088 9088 49094
rect 9036 49030 9088 49036
rect 9048 45554 9076 49030
rect 8772 45526 9076 45554
rect 8668 34536 8720 34542
rect 8668 34478 8720 34484
rect 8208 31340 8260 31346
rect 8208 31282 8260 31288
rect 8484 29844 8536 29850
rect 8484 29786 8536 29792
rect 8300 29640 8352 29646
rect 8300 29582 8352 29588
rect 8312 28558 8340 29582
rect 8496 29510 8524 29786
rect 8484 29504 8536 29510
rect 8484 29446 8536 29452
rect 8300 28552 8352 28558
rect 8300 28494 8352 28500
rect 8208 28416 8260 28422
rect 8208 28358 8260 28364
rect 8300 28416 8352 28422
rect 8300 28358 8352 28364
rect 8220 19854 8248 28358
rect 8312 22642 8340 28358
rect 8392 27124 8444 27130
rect 8392 27066 8444 27072
rect 8300 22636 8352 22642
rect 8300 22578 8352 22584
rect 8208 19848 8260 19854
rect 8208 19790 8260 19796
rect 7288 3052 7340 3058
rect 7288 2994 7340 3000
rect 8116 3052 8168 3058
rect 8116 2994 8168 3000
rect 8312 2990 8340 22578
rect 8404 22098 8432 27066
rect 8668 26988 8720 26994
rect 8668 26930 8720 26936
rect 8680 22574 8708 26930
rect 8668 22568 8720 22574
rect 8668 22510 8720 22516
rect 8392 22092 8444 22098
rect 8392 22034 8444 22040
rect 8680 19378 8708 22510
rect 8668 19372 8720 19378
rect 8668 19314 8720 19320
rect 8680 17610 8708 19314
rect 8668 17604 8720 17610
rect 8668 17546 8720 17552
rect 8484 3732 8536 3738
rect 8484 3674 8536 3680
rect 8496 3058 8524 3674
rect 8772 3058 8800 45526
rect 9232 38418 9260 69362
rect 11950 69116 12258 69125
rect 11950 69114 11956 69116
rect 12012 69114 12036 69116
rect 12092 69114 12116 69116
rect 12172 69114 12196 69116
rect 12252 69114 12258 69116
rect 12012 69062 12014 69114
rect 12194 69062 12196 69114
rect 11950 69060 11956 69062
rect 12012 69060 12036 69062
rect 12092 69060 12116 69062
rect 12172 69060 12196 69062
rect 12252 69060 12258 69062
rect 11950 69051 12258 69060
rect 12610 68572 12918 68581
rect 12610 68570 12616 68572
rect 12672 68570 12696 68572
rect 12752 68570 12776 68572
rect 12832 68570 12856 68572
rect 12912 68570 12918 68572
rect 12672 68518 12674 68570
rect 12854 68518 12856 68570
rect 12610 68516 12616 68518
rect 12672 68516 12696 68518
rect 12752 68516 12776 68518
rect 12832 68516 12856 68518
rect 12912 68516 12918 68518
rect 12610 68507 12918 68516
rect 9588 68196 9640 68202
rect 9588 68138 9640 68144
rect 9312 68128 9364 68134
rect 9312 68070 9364 68076
rect 9220 38412 9272 38418
rect 9220 38354 9272 38360
rect 9220 36780 9272 36786
rect 9220 36722 9272 36728
rect 9232 33658 9260 36722
rect 9220 33652 9272 33658
rect 9220 33594 9272 33600
rect 9036 30864 9088 30870
rect 9036 30806 9088 30812
rect 9048 30705 9076 30806
rect 9034 30696 9090 30705
rect 9034 30631 9090 30640
rect 9220 26784 9272 26790
rect 9220 26726 9272 26732
rect 9232 18154 9260 26726
rect 9220 18148 9272 18154
rect 9220 18090 9272 18096
rect 9128 17604 9180 17610
rect 9128 17546 9180 17552
rect 8484 3052 8536 3058
rect 8484 2994 8536 3000
rect 8760 3052 8812 3058
rect 8760 2994 8812 3000
rect 8300 2984 8352 2990
rect 8300 2926 8352 2932
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 6950 2748 7258 2757
rect 6950 2746 6956 2748
rect 7012 2746 7036 2748
rect 7092 2746 7116 2748
rect 7172 2746 7196 2748
rect 7252 2746 7258 2748
rect 7012 2694 7014 2746
rect 7194 2694 7196 2746
rect 6950 2692 6956 2694
rect 7012 2692 7036 2694
rect 7092 2692 7116 2694
rect 7172 2692 7196 2694
rect 7252 2692 7258 2694
rect 6950 2683 7258 2692
rect 9140 2446 9168 17546
rect 9324 8974 9352 68070
rect 9600 55214 9628 68138
rect 11950 68028 12258 68037
rect 11950 68026 11956 68028
rect 12012 68026 12036 68028
rect 12092 68026 12116 68028
rect 12172 68026 12196 68028
rect 12252 68026 12258 68028
rect 12012 67974 12014 68026
rect 12194 67974 12196 68026
rect 11950 67972 11956 67974
rect 12012 67972 12036 67974
rect 12092 67972 12116 67974
rect 12172 67972 12196 67974
rect 12252 67972 12258 67974
rect 11950 67963 12258 67972
rect 12610 67484 12918 67493
rect 12610 67482 12616 67484
rect 12672 67482 12696 67484
rect 12752 67482 12776 67484
rect 12832 67482 12856 67484
rect 12912 67482 12918 67484
rect 12672 67430 12674 67482
rect 12854 67430 12856 67482
rect 12610 67428 12616 67430
rect 12672 67428 12696 67430
rect 12752 67428 12776 67430
rect 12832 67428 12856 67430
rect 12912 67428 12918 67430
rect 12610 67419 12918 67428
rect 14280 67244 14332 67250
rect 14280 67186 14332 67192
rect 14188 67176 14240 67182
rect 14188 67118 14240 67124
rect 11950 66940 12258 66949
rect 11950 66938 11956 66940
rect 12012 66938 12036 66940
rect 12092 66938 12116 66940
rect 12172 66938 12196 66940
rect 12252 66938 12258 66940
rect 12012 66886 12014 66938
rect 12194 66886 12196 66938
rect 11950 66884 11956 66886
rect 12012 66884 12036 66886
rect 12092 66884 12116 66886
rect 12172 66884 12196 66886
rect 12252 66884 12258 66886
rect 11950 66875 12258 66884
rect 12610 66396 12918 66405
rect 12610 66394 12616 66396
rect 12672 66394 12696 66396
rect 12752 66394 12776 66396
rect 12832 66394 12856 66396
rect 12912 66394 12918 66396
rect 12672 66342 12674 66394
rect 12854 66342 12856 66394
rect 12610 66340 12616 66342
rect 12672 66340 12696 66342
rect 12752 66340 12776 66342
rect 12832 66340 12856 66342
rect 12912 66340 12918 66342
rect 12610 66331 12918 66340
rect 11950 65852 12258 65861
rect 11950 65850 11956 65852
rect 12012 65850 12036 65852
rect 12092 65850 12116 65852
rect 12172 65850 12196 65852
rect 12252 65850 12258 65852
rect 12012 65798 12014 65850
rect 12194 65798 12196 65850
rect 11950 65796 11956 65798
rect 12012 65796 12036 65798
rect 12092 65796 12116 65798
rect 12172 65796 12196 65798
rect 12252 65796 12258 65798
rect 11950 65787 12258 65796
rect 12610 65308 12918 65317
rect 12610 65306 12616 65308
rect 12672 65306 12696 65308
rect 12752 65306 12776 65308
rect 12832 65306 12856 65308
rect 12912 65306 12918 65308
rect 12672 65254 12674 65306
rect 12854 65254 12856 65306
rect 12610 65252 12616 65254
rect 12672 65252 12696 65254
rect 12752 65252 12776 65254
rect 12832 65252 12856 65254
rect 12912 65252 12918 65254
rect 12610 65243 12918 65252
rect 10692 65000 10744 65006
rect 10692 64942 10744 64948
rect 10784 65000 10836 65006
rect 10784 64942 10836 64948
rect 10968 65000 11020 65006
rect 10968 64942 11020 64948
rect 10508 57928 10560 57934
rect 10508 57870 10560 57876
rect 10520 56846 10548 57870
rect 10508 56840 10560 56846
rect 10508 56782 10560 56788
rect 9508 55186 9628 55214
rect 9404 48748 9456 48754
rect 9404 48690 9456 48696
rect 9416 36378 9444 48690
rect 9404 36372 9456 36378
rect 9404 36314 9456 36320
rect 9508 35894 9536 55186
rect 9772 54188 9824 54194
rect 9772 54130 9824 54136
rect 9588 45960 9640 45966
rect 9588 45902 9640 45908
rect 9600 45626 9628 45902
rect 9588 45620 9640 45626
rect 9588 45562 9640 45568
rect 9600 38894 9628 45562
rect 9588 38888 9640 38894
rect 9588 38830 9640 38836
rect 9508 35866 9628 35894
rect 9496 30796 9548 30802
rect 9496 30738 9548 30744
rect 9312 8968 9364 8974
rect 9312 8910 9364 8916
rect 9508 8090 9536 30738
rect 9600 25498 9628 35866
rect 9588 25492 9640 25498
rect 9588 25434 9640 25440
rect 9680 23792 9732 23798
rect 9680 23734 9732 23740
rect 9588 22228 9640 22234
rect 9588 22170 9640 22176
rect 9600 19514 9628 22170
rect 9588 19508 9640 19514
rect 9588 19450 9640 19456
rect 9600 18834 9628 19450
rect 9588 18828 9640 18834
rect 9588 18770 9640 18776
rect 9600 13870 9628 18770
rect 9588 13864 9640 13870
rect 9588 13806 9640 13812
rect 9600 9382 9628 13806
rect 9588 9376 9640 9382
rect 9588 9318 9640 9324
rect 9496 8084 9548 8090
rect 9496 8026 9548 8032
rect 9692 6914 9720 23734
rect 9784 14074 9812 54130
rect 10416 52012 10468 52018
rect 10416 51954 10468 51960
rect 10232 51944 10284 51950
rect 10232 51886 10284 51892
rect 9864 27940 9916 27946
rect 9864 27882 9916 27888
rect 9876 22982 9904 27882
rect 9864 22976 9916 22982
rect 9864 22918 9916 22924
rect 9864 18692 9916 18698
rect 9864 18634 9916 18640
rect 9876 18426 9904 18634
rect 9864 18420 9916 18426
rect 9864 18362 9916 18368
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 9692 6886 9812 6914
rect 9496 3392 9548 3398
rect 9496 3334 9548 3340
rect 9508 3058 9536 3334
rect 9496 3052 9548 3058
rect 9496 2994 9548 3000
rect 9784 2990 9812 6886
rect 9772 2984 9824 2990
rect 9772 2926 9824 2932
rect 2504 2440 2556 2446
rect 2504 2382 2556 2388
rect 9128 2440 9180 2446
rect 9128 2382 9180 2388
rect 2516 1306 2544 2382
rect 10244 2378 10272 51886
rect 10324 47048 10376 47054
rect 10324 46990 10376 46996
rect 10336 23118 10364 46990
rect 10428 45082 10456 51954
rect 10416 45076 10468 45082
rect 10416 45018 10468 45024
rect 10428 44946 10456 45018
rect 10416 44940 10468 44946
rect 10416 44882 10468 44888
rect 10520 33658 10548 56782
rect 10600 40724 10652 40730
rect 10600 40666 10652 40672
rect 10508 33652 10560 33658
rect 10508 33594 10560 33600
rect 10416 33312 10468 33318
rect 10416 33254 10468 33260
rect 10324 23112 10376 23118
rect 10324 23054 10376 23060
rect 10428 9586 10456 33254
rect 10612 27946 10640 40666
rect 10704 34134 10732 64942
rect 10796 57934 10824 64942
rect 10784 57928 10836 57934
rect 10784 57870 10836 57876
rect 10784 51332 10836 51338
rect 10784 51274 10836 51280
rect 10796 40730 10824 51274
rect 10980 49842 11008 64942
rect 11950 64764 12258 64773
rect 11950 64762 11956 64764
rect 12012 64762 12036 64764
rect 12092 64762 12116 64764
rect 12172 64762 12196 64764
rect 12252 64762 12258 64764
rect 12012 64710 12014 64762
rect 12194 64710 12196 64762
rect 11950 64708 11956 64710
rect 12012 64708 12036 64710
rect 12092 64708 12116 64710
rect 12172 64708 12196 64710
rect 12252 64708 12258 64710
rect 11950 64699 12258 64708
rect 11060 64456 11112 64462
rect 11060 64398 11112 64404
rect 12348 64456 12400 64462
rect 12348 64398 12400 64404
rect 11072 52154 11100 64398
rect 11796 64320 11848 64326
rect 11796 64262 11848 64268
rect 11244 62348 11296 62354
rect 11244 62290 11296 62296
rect 11060 52148 11112 52154
rect 11060 52090 11112 52096
rect 11256 51406 11284 62290
rect 11336 62144 11388 62150
rect 11336 62086 11388 62092
rect 11244 51400 11296 51406
rect 11244 51342 11296 51348
rect 11348 51338 11376 62086
rect 11704 51468 11756 51474
rect 11704 51410 11756 51416
rect 11336 51332 11388 51338
rect 11336 51274 11388 51280
rect 11612 51264 11664 51270
rect 11612 51206 11664 51212
rect 10968 49836 11020 49842
rect 10968 49778 11020 49784
rect 10784 40724 10836 40730
rect 10784 40666 10836 40672
rect 11624 35894 11652 51206
rect 11532 35866 11652 35894
rect 10692 34128 10744 34134
rect 10692 34070 10744 34076
rect 10704 33318 10732 34070
rect 10692 33312 10744 33318
rect 10692 33254 10744 33260
rect 11336 30660 11388 30666
rect 11336 30602 11388 30608
rect 11348 30394 11376 30602
rect 11336 30388 11388 30394
rect 11336 30330 11388 30336
rect 11532 30326 11560 35866
rect 11612 30796 11664 30802
rect 11612 30738 11664 30744
rect 11520 30320 11572 30326
rect 11520 30262 11572 30268
rect 11532 28558 11560 30262
rect 11624 29714 11652 30738
rect 11716 30258 11744 51410
rect 11808 31770 11836 64262
rect 11950 63676 12258 63685
rect 11950 63674 11956 63676
rect 12012 63674 12036 63676
rect 12092 63674 12116 63676
rect 12172 63674 12196 63676
rect 12252 63674 12258 63676
rect 12012 63622 12014 63674
rect 12194 63622 12196 63674
rect 11950 63620 11956 63622
rect 12012 63620 12036 63622
rect 12092 63620 12116 63622
rect 12172 63620 12196 63622
rect 12252 63620 12258 63622
rect 11950 63611 12258 63620
rect 11950 62588 12258 62597
rect 11950 62586 11956 62588
rect 12012 62586 12036 62588
rect 12092 62586 12116 62588
rect 12172 62586 12196 62588
rect 12252 62586 12258 62588
rect 12012 62534 12014 62586
rect 12194 62534 12196 62586
rect 11950 62532 11956 62534
rect 12012 62532 12036 62534
rect 12092 62532 12116 62534
rect 12172 62532 12196 62534
rect 12252 62532 12258 62534
rect 11950 62523 12258 62532
rect 11950 61500 12258 61509
rect 11950 61498 11956 61500
rect 12012 61498 12036 61500
rect 12092 61498 12116 61500
rect 12172 61498 12196 61500
rect 12252 61498 12258 61500
rect 12012 61446 12014 61498
rect 12194 61446 12196 61498
rect 11950 61444 11956 61446
rect 12012 61444 12036 61446
rect 12092 61444 12116 61446
rect 12172 61444 12196 61446
rect 12252 61444 12258 61446
rect 11950 61435 12258 61444
rect 11950 60412 12258 60421
rect 11950 60410 11956 60412
rect 12012 60410 12036 60412
rect 12092 60410 12116 60412
rect 12172 60410 12196 60412
rect 12252 60410 12258 60412
rect 12012 60358 12014 60410
rect 12194 60358 12196 60410
rect 11950 60356 11956 60358
rect 12012 60356 12036 60358
rect 12092 60356 12116 60358
rect 12172 60356 12196 60358
rect 12252 60356 12258 60358
rect 11950 60347 12258 60356
rect 11950 59324 12258 59333
rect 11950 59322 11956 59324
rect 12012 59322 12036 59324
rect 12092 59322 12116 59324
rect 12172 59322 12196 59324
rect 12252 59322 12258 59324
rect 12012 59270 12014 59322
rect 12194 59270 12196 59322
rect 11950 59268 11956 59270
rect 12012 59268 12036 59270
rect 12092 59268 12116 59270
rect 12172 59268 12196 59270
rect 12252 59268 12258 59270
rect 11950 59259 12258 59268
rect 11950 58236 12258 58245
rect 11950 58234 11956 58236
rect 12012 58234 12036 58236
rect 12092 58234 12116 58236
rect 12172 58234 12196 58236
rect 12252 58234 12258 58236
rect 12012 58182 12014 58234
rect 12194 58182 12196 58234
rect 11950 58180 11956 58182
rect 12012 58180 12036 58182
rect 12092 58180 12116 58182
rect 12172 58180 12196 58182
rect 12252 58180 12258 58182
rect 11950 58171 12258 58180
rect 11950 57148 12258 57157
rect 11950 57146 11956 57148
rect 12012 57146 12036 57148
rect 12092 57146 12116 57148
rect 12172 57146 12196 57148
rect 12252 57146 12258 57148
rect 12012 57094 12014 57146
rect 12194 57094 12196 57146
rect 11950 57092 11956 57094
rect 12012 57092 12036 57094
rect 12092 57092 12116 57094
rect 12172 57092 12196 57094
rect 12252 57092 12258 57094
rect 11950 57083 12258 57092
rect 11950 56060 12258 56069
rect 11950 56058 11956 56060
rect 12012 56058 12036 56060
rect 12092 56058 12116 56060
rect 12172 56058 12196 56060
rect 12252 56058 12258 56060
rect 12012 56006 12014 56058
rect 12194 56006 12196 56058
rect 11950 56004 11956 56006
rect 12012 56004 12036 56006
rect 12092 56004 12116 56006
rect 12172 56004 12196 56006
rect 12252 56004 12258 56006
rect 11950 55995 12258 56004
rect 12360 55894 12388 64398
rect 12610 64220 12918 64229
rect 12610 64218 12616 64220
rect 12672 64218 12696 64220
rect 12752 64218 12776 64220
rect 12832 64218 12856 64220
rect 12912 64218 12918 64220
rect 12672 64166 12674 64218
rect 12854 64166 12856 64218
rect 12610 64164 12616 64166
rect 12672 64164 12696 64166
rect 12752 64164 12776 64166
rect 12832 64164 12856 64166
rect 12912 64164 12918 64166
rect 12610 64155 12918 64164
rect 14096 63776 14148 63782
rect 14096 63718 14148 63724
rect 12610 63132 12918 63141
rect 12610 63130 12616 63132
rect 12672 63130 12696 63132
rect 12752 63130 12776 63132
rect 12832 63130 12856 63132
rect 12912 63130 12918 63132
rect 12672 63078 12674 63130
rect 12854 63078 12856 63130
rect 12610 63076 12616 63078
rect 12672 63076 12696 63078
rect 12752 63076 12776 63078
rect 12832 63076 12856 63078
rect 12912 63076 12918 63078
rect 12610 63067 12918 63076
rect 12610 62044 12918 62053
rect 12610 62042 12616 62044
rect 12672 62042 12696 62044
rect 12752 62042 12776 62044
rect 12832 62042 12856 62044
rect 12912 62042 12918 62044
rect 12672 61990 12674 62042
rect 12854 61990 12856 62042
rect 12610 61988 12616 61990
rect 12672 61988 12696 61990
rect 12752 61988 12776 61990
rect 12832 61988 12856 61990
rect 12912 61988 12918 61990
rect 12610 61979 12918 61988
rect 12610 60956 12918 60965
rect 12610 60954 12616 60956
rect 12672 60954 12696 60956
rect 12752 60954 12776 60956
rect 12832 60954 12856 60956
rect 12912 60954 12918 60956
rect 12672 60902 12674 60954
rect 12854 60902 12856 60954
rect 12610 60900 12616 60902
rect 12672 60900 12696 60902
rect 12752 60900 12776 60902
rect 12832 60900 12856 60902
rect 12912 60900 12918 60902
rect 12610 60891 12918 60900
rect 12610 59868 12918 59877
rect 12610 59866 12616 59868
rect 12672 59866 12696 59868
rect 12752 59866 12776 59868
rect 12832 59866 12856 59868
rect 12912 59866 12918 59868
rect 12672 59814 12674 59866
rect 12854 59814 12856 59866
rect 12610 59812 12616 59814
rect 12672 59812 12696 59814
rect 12752 59812 12776 59814
rect 12832 59812 12856 59814
rect 12912 59812 12918 59814
rect 12610 59803 12918 59812
rect 12610 58780 12918 58789
rect 12610 58778 12616 58780
rect 12672 58778 12696 58780
rect 12752 58778 12776 58780
rect 12832 58778 12856 58780
rect 12912 58778 12918 58780
rect 12672 58726 12674 58778
rect 12854 58726 12856 58778
rect 12610 58724 12616 58726
rect 12672 58724 12696 58726
rect 12752 58724 12776 58726
rect 12832 58724 12856 58726
rect 12912 58724 12918 58726
rect 12610 58715 12918 58724
rect 12610 57692 12918 57701
rect 12610 57690 12616 57692
rect 12672 57690 12696 57692
rect 12752 57690 12776 57692
rect 12832 57690 12856 57692
rect 12912 57690 12918 57692
rect 12672 57638 12674 57690
rect 12854 57638 12856 57690
rect 12610 57636 12616 57638
rect 12672 57636 12696 57638
rect 12752 57636 12776 57638
rect 12832 57636 12856 57638
rect 12912 57636 12918 57638
rect 12610 57627 12918 57636
rect 12610 56604 12918 56613
rect 12610 56602 12616 56604
rect 12672 56602 12696 56604
rect 12752 56602 12776 56604
rect 12832 56602 12856 56604
rect 12912 56602 12918 56604
rect 12672 56550 12674 56602
rect 12854 56550 12856 56602
rect 12610 56548 12616 56550
rect 12672 56548 12696 56550
rect 12752 56548 12776 56550
rect 12832 56548 12856 56550
rect 12912 56548 12918 56550
rect 12610 56539 12918 56548
rect 12348 55888 12400 55894
rect 12348 55830 12400 55836
rect 12610 55516 12918 55525
rect 12610 55514 12616 55516
rect 12672 55514 12696 55516
rect 12752 55514 12776 55516
rect 12832 55514 12856 55516
rect 12912 55514 12918 55516
rect 12672 55462 12674 55514
rect 12854 55462 12856 55514
rect 12610 55460 12616 55462
rect 12672 55460 12696 55462
rect 12752 55460 12776 55462
rect 12832 55460 12856 55462
rect 12912 55460 12918 55462
rect 12610 55451 12918 55460
rect 11950 54972 12258 54981
rect 11950 54970 11956 54972
rect 12012 54970 12036 54972
rect 12092 54970 12116 54972
rect 12172 54970 12196 54972
rect 12252 54970 12258 54972
rect 12012 54918 12014 54970
rect 12194 54918 12196 54970
rect 11950 54916 11956 54918
rect 12012 54916 12036 54918
rect 12092 54916 12116 54918
rect 12172 54916 12196 54918
rect 12252 54916 12258 54918
rect 11950 54907 12258 54916
rect 12610 54428 12918 54437
rect 12610 54426 12616 54428
rect 12672 54426 12696 54428
rect 12752 54426 12776 54428
rect 12832 54426 12856 54428
rect 12912 54426 12918 54428
rect 12672 54374 12674 54426
rect 12854 54374 12856 54426
rect 12610 54372 12616 54374
rect 12672 54372 12696 54374
rect 12752 54372 12776 54374
rect 12832 54372 12856 54374
rect 12912 54372 12918 54374
rect 12610 54363 12918 54372
rect 13820 53984 13872 53990
rect 13820 53926 13872 53932
rect 11950 53884 12258 53893
rect 11950 53882 11956 53884
rect 12012 53882 12036 53884
rect 12092 53882 12116 53884
rect 12172 53882 12196 53884
rect 12252 53882 12258 53884
rect 12012 53830 12014 53882
rect 12194 53830 12196 53882
rect 11950 53828 11956 53830
rect 12012 53828 12036 53830
rect 12092 53828 12116 53830
rect 12172 53828 12196 53830
rect 12252 53828 12258 53830
rect 11950 53819 12258 53828
rect 13544 53576 13596 53582
rect 13544 53518 13596 53524
rect 12610 53340 12918 53349
rect 12610 53338 12616 53340
rect 12672 53338 12696 53340
rect 12752 53338 12776 53340
rect 12832 53338 12856 53340
rect 12912 53338 12918 53340
rect 12672 53286 12674 53338
rect 12854 53286 12856 53338
rect 12610 53284 12616 53286
rect 12672 53284 12696 53286
rect 12752 53284 12776 53286
rect 12832 53284 12856 53286
rect 12912 53284 12918 53286
rect 12610 53275 12918 53284
rect 11950 52796 12258 52805
rect 11950 52794 11956 52796
rect 12012 52794 12036 52796
rect 12092 52794 12116 52796
rect 12172 52794 12196 52796
rect 12252 52794 12258 52796
rect 12012 52742 12014 52794
rect 12194 52742 12196 52794
rect 11950 52740 11956 52742
rect 12012 52740 12036 52742
rect 12092 52740 12116 52742
rect 12172 52740 12196 52742
rect 12252 52740 12258 52742
rect 11950 52731 12258 52740
rect 12610 52252 12918 52261
rect 12610 52250 12616 52252
rect 12672 52250 12696 52252
rect 12752 52250 12776 52252
rect 12832 52250 12856 52252
rect 12912 52250 12918 52252
rect 12672 52198 12674 52250
rect 12854 52198 12856 52250
rect 12610 52196 12616 52198
rect 12672 52196 12696 52198
rect 12752 52196 12776 52198
rect 12832 52196 12856 52198
rect 12912 52196 12918 52198
rect 12610 52187 12918 52196
rect 12348 52148 12400 52154
rect 12348 52090 12400 52096
rect 11950 51708 12258 51717
rect 11950 51706 11956 51708
rect 12012 51706 12036 51708
rect 12092 51706 12116 51708
rect 12172 51706 12196 51708
rect 12252 51706 12258 51708
rect 12012 51654 12014 51706
rect 12194 51654 12196 51706
rect 11950 51652 11956 51654
rect 12012 51652 12036 51654
rect 12092 51652 12116 51654
rect 12172 51652 12196 51654
rect 12252 51652 12258 51654
rect 11950 51643 12258 51652
rect 11950 50620 12258 50629
rect 11950 50618 11956 50620
rect 12012 50618 12036 50620
rect 12092 50618 12116 50620
rect 12172 50618 12196 50620
rect 12252 50618 12258 50620
rect 12012 50566 12014 50618
rect 12194 50566 12196 50618
rect 11950 50564 11956 50566
rect 12012 50564 12036 50566
rect 12092 50564 12116 50566
rect 12172 50564 12196 50566
rect 12252 50564 12258 50566
rect 11950 50555 12258 50564
rect 11950 49532 12258 49541
rect 11950 49530 11956 49532
rect 12012 49530 12036 49532
rect 12092 49530 12116 49532
rect 12172 49530 12196 49532
rect 12252 49530 12258 49532
rect 12012 49478 12014 49530
rect 12194 49478 12196 49530
rect 11950 49476 11956 49478
rect 12012 49476 12036 49478
rect 12092 49476 12116 49478
rect 12172 49476 12196 49478
rect 12252 49476 12258 49478
rect 11950 49467 12258 49476
rect 11950 48444 12258 48453
rect 11950 48442 11956 48444
rect 12012 48442 12036 48444
rect 12092 48442 12116 48444
rect 12172 48442 12196 48444
rect 12252 48442 12258 48444
rect 12012 48390 12014 48442
rect 12194 48390 12196 48442
rect 11950 48388 11956 48390
rect 12012 48388 12036 48390
rect 12092 48388 12116 48390
rect 12172 48388 12196 48390
rect 12252 48388 12258 48390
rect 11950 48379 12258 48388
rect 11950 47356 12258 47365
rect 11950 47354 11956 47356
rect 12012 47354 12036 47356
rect 12092 47354 12116 47356
rect 12172 47354 12196 47356
rect 12252 47354 12258 47356
rect 12012 47302 12014 47354
rect 12194 47302 12196 47354
rect 11950 47300 11956 47302
rect 12012 47300 12036 47302
rect 12092 47300 12116 47302
rect 12172 47300 12196 47302
rect 12252 47300 12258 47302
rect 11950 47291 12258 47300
rect 11950 46268 12258 46277
rect 11950 46266 11956 46268
rect 12012 46266 12036 46268
rect 12092 46266 12116 46268
rect 12172 46266 12196 46268
rect 12252 46266 12258 46268
rect 12012 46214 12014 46266
rect 12194 46214 12196 46266
rect 11950 46212 11956 46214
rect 12012 46212 12036 46214
rect 12092 46212 12116 46214
rect 12172 46212 12196 46214
rect 12252 46212 12258 46214
rect 11950 46203 12258 46212
rect 11950 45180 12258 45189
rect 11950 45178 11956 45180
rect 12012 45178 12036 45180
rect 12092 45178 12116 45180
rect 12172 45178 12196 45180
rect 12252 45178 12258 45180
rect 12012 45126 12014 45178
rect 12194 45126 12196 45178
rect 11950 45124 11956 45126
rect 12012 45124 12036 45126
rect 12092 45124 12116 45126
rect 12172 45124 12196 45126
rect 12252 45124 12258 45126
rect 11950 45115 12258 45124
rect 11950 44092 12258 44101
rect 11950 44090 11956 44092
rect 12012 44090 12036 44092
rect 12092 44090 12116 44092
rect 12172 44090 12196 44092
rect 12252 44090 12258 44092
rect 12012 44038 12014 44090
rect 12194 44038 12196 44090
rect 11950 44036 11956 44038
rect 12012 44036 12036 44038
rect 12092 44036 12116 44038
rect 12172 44036 12196 44038
rect 12252 44036 12258 44038
rect 11950 44027 12258 44036
rect 11950 43004 12258 43013
rect 11950 43002 11956 43004
rect 12012 43002 12036 43004
rect 12092 43002 12116 43004
rect 12172 43002 12196 43004
rect 12252 43002 12258 43004
rect 12012 42950 12014 43002
rect 12194 42950 12196 43002
rect 11950 42948 11956 42950
rect 12012 42948 12036 42950
rect 12092 42948 12116 42950
rect 12172 42948 12196 42950
rect 12252 42948 12258 42950
rect 11950 42939 12258 42948
rect 11950 41916 12258 41925
rect 11950 41914 11956 41916
rect 12012 41914 12036 41916
rect 12092 41914 12116 41916
rect 12172 41914 12196 41916
rect 12252 41914 12258 41916
rect 12012 41862 12014 41914
rect 12194 41862 12196 41914
rect 11950 41860 11956 41862
rect 12012 41860 12036 41862
rect 12092 41860 12116 41862
rect 12172 41860 12196 41862
rect 12252 41860 12258 41862
rect 11950 41851 12258 41860
rect 11950 40828 12258 40837
rect 11950 40826 11956 40828
rect 12012 40826 12036 40828
rect 12092 40826 12116 40828
rect 12172 40826 12196 40828
rect 12252 40826 12258 40828
rect 12012 40774 12014 40826
rect 12194 40774 12196 40826
rect 11950 40772 11956 40774
rect 12012 40772 12036 40774
rect 12092 40772 12116 40774
rect 12172 40772 12196 40774
rect 12252 40772 12258 40774
rect 11950 40763 12258 40772
rect 11950 39740 12258 39749
rect 11950 39738 11956 39740
rect 12012 39738 12036 39740
rect 12092 39738 12116 39740
rect 12172 39738 12196 39740
rect 12252 39738 12258 39740
rect 12012 39686 12014 39738
rect 12194 39686 12196 39738
rect 11950 39684 11956 39686
rect 12012 39684 12036 39686
rect 12092 39684 12116 39686
rect 12172 39684 12196 39686
rect 12252 39684 12258 39686
rect 11950 39675 12258 39684
rect 11950 38652 12258 38661
rect 11950 38650 11956 38652
rect 12012 38650 12036 38652
rect 12092 38650 12116 38652
rect 12172 38650 12196 38652
rect 12252 38650 12258 38652
rect 12012 38598 12014 38650
rect 12194 38598 12196 38650
rect 11950 38596 11956 38598
rect 12012 38596 12036 38598
rect 12092 38596 12116 38598
rect 12172 38596 12196 38598
rect 12252 38596 12258 38598
rect 11950 38587 12258 38596
rect 11950 37564 12258 37573
rect 11950 37562 11956 37564
rect 12012 37562 12036 37564
rect 12092 37562 12116 37564
rect 12172 37562 12196 37564
rect 12252 37562 12258 37564
rect 12012 37510 12014 37562
rect 12194 37510 12196 37562
rect 11950 37508 11956 37510
rect 12012 37508 12036 37510
rect 12092 37508 12116 37510
rect 12172 37508 12196 37510
rect 12252 37508 12258 37510
rect 11950 37499 12258 37508
rect 11950 36476 12258 36485
rect 11950 36474 11956 36476
rect 12012 36474 12036 36476
rect 12092 36474 12116 36476
rect 12172 36474 12196 36476
rect 12252 36474 12258 36476
rect 12012 36422 12014 36474
rect 12194 36422 12196 36474
rect 11950 36420 11956 36422
rect 12012 36420 12036 36422
rect 12092 36420 12116 36422
rect 12172 36420 12196 36422
rect 12252 36420 12258 36422
rect 11950 36411 12258 36420
rect 11950 35388 12258 35397
rect 11950 35386 11956 35388
rect 12012 35386 12036 35388
rect 12092 35386 12116 35388
rect 12172 35386 12196 35388
rect 12252 35386 12258 35388
rect 12012 35334 12014 35386
rect 12194 35334 12196 35386
rect 11950 35332 11956 35334
rect 12012 35332 12036 35334
rect 12092 35332 12116 35334
rect 12172 35332 12196 35334
rect 12252 35332 12258 35334
rect 11950 35323 12258 35332
rect 11950 34300 12258 34309
rect 11950 34298 11956 34300
rect 12012 34298 12036 34300
rect 12092 34298 12116 34300
rect 12172 34298 12196 34300
rect 12252 34298 12258 34300
rect 12012 34246 12014 34298
rect 12194 34246 12196 34298
rect 11950 34244 11956 34246
rect 12012 34244 12036 34246
rect 12092 34244 12116 34246
rect 12172 34244 12196 34246
rect 12252 34244 12258 34246
rect 11950 34235 12258 34244
rect 11950 33212 12258 33221
rect 11950 33210 11956 33212
rect 12012 33210 12036 33212
rect 12092 33210 12116 33212
rect 12172 33210 12196 33212
rect 12252 33210 12258 33212
rect 12012 33158 12014 33210
rect 12194 33158 12196 33210
rect 11950 33156 11956 33158
rect 12012 33156 12036 33158
rect 12092 33156 12116 33158
rect 12172 33156 12196 33158
rect 12252 33156 12258 33158
rect 11950 33147 12258 33156
rect 11950 32124 12258 32133
rect 11950 32122 11956 32124
rect 12012 32122 12036 32124
rect 12092 32122 12116 32124
rect 12172 32122 12196 32124
rect 12252 32122 12258 32124
rect 12012 32070 12014 32122
rect 12194 32070 12196 32122
rect 11950 32068 11956 32070
rect 12012 32068 12036 32070
rect 12092 32068 12116 32070
rect 12172 32068 12196 32070
rect 12252 32068 12258 32070
rect 11950 32059 12258 32068
rect 12360 31906 12388 52090
rect 12610 51164 12918 51173
rect 12610 51162 12616 51164
rect 12672 51162 12696 51164
rect 12752 51162 12776 51164
rect 12832 51162 12856 51164
rect 12912 51162 12918 51164
rect 12672 51110 12674 51162
rect 12854 51110 12856 51162
rect 12610 51108 12616 51110
rect 12672 51108 12696 51110
rect 12752 51108 12776 51110
rect 12832 51108 12856 51110
rect 12912 51108 12918 51110
rect 12610 51099 12918 51108
rect 13084 50924 13136 50930
rect 13084 50866 13136 50872
rect 12440 50856 12492 50862
rect 12440 50798 12492 50804
rect 12452 48754 12480 50798
rect 12992 50788 13044 50794
rect 12992 50730 13044 50736
rect 12610 50076 12918 50085
rect 12610 50074 12616 50076
rect 12672 50074 12696 50076
rect 12752 50074 12776 50076
rect 12832 50074 12856 50076
rect 12912 50074 12918 50076
rect 12672 50022 12674 50074
rect 12854 50022 12856 50074
rect 12610 50020 12616 50022
rect 12672 50020 12696 50022
rect 12752 50020 12776 50022
rect 12832 50020 12856 50022
rect 12912 50020 12918 50022
rect 12610 50011 12918 50020
rect 12610 48988 12918 48997
rect 12610 48986 12616 48988
rect 12672 48986 12696 48988
rect 12752 48986 12776 48988
rect 12832 48986 12856 48988
rect 12912 48986 12918 48988
rect 12672 48934 12674 48986
rect 12854 48934 12856 48986
rect 12610 48932 12616 48934
rect 12672 48932 12696 48934
rect 12752 48932 12776 48934
rect 12832 48932 12856 48934
rect 12912 48932 12918 48934
rect 12610 48923 12918 48932
rect 12440 48748 12492 48754
rect 12440 48690 12492 48696
rect 12610 47900 12918 47909
rect 12610 47898 12616 47900
rect 12672 47898 12696 47900
rect 12752 47898 12776 47900
rect 12832 47898 12856 47900
rect 12912 47898 12918 47900
rect 12672 47846 12674 47898
rect 12854 47846 12856 47898
rect 12610 47844 12616 47846
rect 12672 47844 12696 47846
rect 12752 47844 12776 47846
rect 12832 47844 12856 47846
rect 12912 47844 12918 47846
rect 12610 47835 12918 47844
rect 12610 46812 12918 46821
rect 12610 46810 12616 46812
rect 12672 46810 12696 46812
rect 12752 46810 12776 46812
rect 12832 46810 12856 46812
rect 12912 46810 12918 46812
rect 12672 46758 12674 46810
rect 12854 46758 12856 46810
rect 12610 46756 12616 46758
rect 12672 46756 12696 46758
rect 12752 46756 12776 46758
rect 12832 46756 12856 46758
rect 12912 46756 12918 46758
rect 12610 46747 12918 46756
rect 12610 45724 12918 45733
rect 12610 45722 12616 45724
rect 12672 45722 12696 45724
rect 12752 45722 12776 45724
rect 12832 45722 12856 45724
rect 12912 45722 12918 45724
rect 12672 45670 12674 45722
rect 12854 45670 12856 45722
rect 12610 45668 12616 45670
rect 12672 45668 12696 45670
rect 12752 45668 12776 45670
rect 12832 45668 12856 45670
rect 12912 45668 12918 45670
rect 12610 45659 12918 45668
rect 12610 44636 12918 44645
rect 12610 44634 12616 44636
rect 12672 44634 12696 44636
rect 12752 44634 12776 44636
rect 12832 44634 12856 44636
rect 12912 44634 12918 44636
rect 12672 44582 12674 44634
rect 12854 44582 12856 44634
rect 12610 44580 12616 44582
rect 12672 44580 12696 44582
rect 12752 44580 12776 44582
rect 12832 44580 12856 44582
rect 12912 44580 12918 44582
rect 12610 44571 12918 44580
rect 12610 43548 12918 43557
rect 12610 43546 12616 43548
rect 12672 43546 12696 43548
rect 12752 43546 12776 43548
rect 12832 43546 12856 43548
rect 12912 43546 12918 43548
rect 12672 43494 12674 43546
rect 12854 43494 12856 43546
rect 12610 43492 12616 43494
rect 12672 43492 12696 43494
rect 12752 43492 12776 43494
rect 12832 43492 12856 43494
rect 12912 43492 12918 43494
rect 12610 43483 12918 43492
rect 12610 42460 12918 42469
rect 12610 42458 12616 42460
rect 12672 42458 12696 42460
rect 12752 42458 12776 42460
rect 12832 42458 12856 42460
rect 12912 42458 12918 42460
rect 12672 42406 12674 42458
rect 12854 42406 12856 42458
rect 12610 42404 12616 42406
rect 12672 42404 12696 42406
rect 12752 42404 12776 42406
rect 12832 42404 12856 42406
rect 12912 42404 12918 42406
rect 12610 42395 12918 42404
rect 12610 41372 12918 41381
rect 12610 41370 12616 41372
rect 12672 41370 12696 41372
rect 12752 41370 12776 41372
rect 12832 41370 12856 41372
rect 12912 41370 12918 41372
rect 12672 41318 12674 41370
rect 12854 41318 12856 41370
rect 12610 41316 12616 41318
rect 12672 41316 12696 41318
rect 12752 41316 12776 41318
rect 12832 41316 12856 41318
rect 12912 41316 12918 41318
rect 12610 41307 12918 41316
rect 12610 40284 12918 40293
rect 12610 40282 12616 40284
rect 12672 40282 12696 40284
rect 12752 40282 12776 40284
rect 12832 40282 12856 40284
rect 12912 40282 12918 40284
rect 12672 40230 12674 40282
rect 12854 40230 12856 40282
rect 12610 40228 12616 40230
rect 12672 40228 12696 40230
rect 12752 40228 12776 40230
rect 12832 40228 12856 40230
rect 12912 40228 12918 40230
rect 12610 40219 12918 40228
rect 12610 39196 12918 39205
rect 12610 39194 12616 39196
rect 12672 39194 12696 39196
rect 12752 39194 12776 39196
rect 12832 39194 12856 39196
rect 12912 39194 12918 39196
rect 12672 39142 12674 39194
rect 12854 39142 12856 39194
rect 12610 39140 12616 39142
rect 12672 39140 12696 39142
rect 12752 39140 12776 39142
rect 12832 39140 12856 39142
rect 12912 39140 12918 39142
rect 12610 39131 12918 39140
rect 13004 38826 13032 50730
rect 12992 38820 13044 38826
rect 12992 38762 13044 38768
rect 12610 38108 12918 38117
rect 12610 38106 12616 38108
rect 12672 38106 12696 38108
rect 12752 38106 12776 38108
rect 12832 38106 12856 38108
rect 12912 38106 12918 38108
rect 12672 38054 12674 38106
rect 12854 38054 12856 38106
rect 12610 38052 12616 38054
rect 12672 38052 12696 38054
rect 12752 38052 12776 38054
rect 12832 38052 12856 38054
rect 12912 38052 12918 38054
rect 12610 38043 12918 38052
rect 12610 37020 12918 37029
rect 12610 37018 12616 37020
rect 12672 37018 12696 37020
rect 12752 37018 12776 37020
rect 12832 37018 12856 37020
rect 12912 37018 12918 37020
rect 12672 36966 12674 37018
rect 12854 36966 12856 37018
rect 12610 36964 12616 36966
rect 12672 36964 12696 36966
rect 12752 36964 12776 36966
rect 12832 36964 12856 36966
rect 12912 36964 12918 36966
rect 12610 36955 12918 36964
rect 12610 35932 12918 35941
rect 12610 35930 12616 35932
rect 12672 35930 12696 35932
rect 12752 35930 12776 35932
rect 12832 35930 12856 35932
rect 12912 35930 12918 35932
rect 12672 35878 12674 35930
rect 12854 35878 12856 35930
rect 12610 35876 12616 35878
rect 12672 35876 12696 35878
rect 12752 35876 12776 35878
rect 12832 35876 12856 35878
rect 12912 35876 12918 35878
rect 12610 35867 12918 35876
rect 12610 34844 12918 34853
rect 12610 34842 12616 34844
rect 12672 34842 12696 34844
rect 12752 34842 12776 34844
rect 12832 34842 12856 34844
rect 12912 34842 12918 34844
rect 12672 34790 12674 34842
rect 12854 34790 12856 34842
rect 12610 34788 12616 34790
rect 12672 34788 12696 34790
rect 12752 34788 12776 34790
rect 12832 34788 12856 34790
rect 12912 34788 12918 34790
rect 12610 34779 12918 34788
rect 12610 33756 12918 33765
rect 12610 33754 12616 33756
rect 12672 33754 12696 33756
rect 12752 33754 12776 33756
rect 12832 33754 12856 33756
rect 12912 33754 12918 33756
rect 12672 33702 12674 33754
rect 12854 33702 12856 33754
rect 12610 33700 12616 33702
rect 12672 33700 12696 33702
rect 12752 33700 12776 33702
rect 12832 33700 12856 33702
rect 12912 33700 12918 33702
rect 12610 33691 12918 33700
rect 12610 32668 12918 32677
rect 12610 32666 12616 32668
rect 12672 32666 12696 32668
rect 12752 32666 12776 32668
rect 12832 32666 12856 32668
rect 12912 32666 12918 32668
rect 12672 32614 12674 32666
rect 12854 32614 12856 32666
rect 12610 32612 12616 32614
rect 12672 32612 12696 32614
rect 12752 32612 12776 32614
rect 12832 32612 12856 32614
rect 12912 32612 12918 32614
rect 12610 32603 12918 32612
rect 13096 32502 13124 50866
rect 13556 41818 13584 53518
rect 13832 52018 13860 53926
rect 13820 52012 13872 52018
rect 13820 51954 13872 51960
rect 13820 47592 13872 47598
rect 13820 47534 13872 47540
rect 13832 47122 13860 47534
rect 13820 47116 13872 47122
rect 13820 47058 13872 47064
rect 13544 41812 13596 41818
rect 13544 41754 13596 41760
rect 13832 41614 13860 47058
rect 13820 41608 13872 41614
rect 13820 41550 13872 41556
rect 13084 32496 13136 32502
rect 13084 32438 13136 32444
rect 12360 31878 12480 31906
rect 11808 31742 12388 31770
rect 11950 31036 12258 31045
rect 11950 31034 11956 31036
rect 12012 31034 12036 31036
rect 12092 31034 12116 31036
rect 12172 31034 12196 31036
rect 12252 31034 12258 31036
rect 12012 30982 12014 31034
rect 12194 30982 12196 31034
rect 11950 30980 11956 30982
rect 12012 30980 12036 30982
rect 12092 30980 12116 30982
rect 12172 30980 12196 30982
rect 12252 30980 12258 30982
rect 11950 30971 12258 30980
rect 11704 30252 11756 30258
rect 11704 30194 11756 30200
rect 11612 29708 11664 29714
rect 11612 29650 11664 29656
rect 11520 28552 11572 28558
rect 11520 28494 11572 28500
rect 10600 27940 10652 27946
rect 10600 27882 10652 27888
rect 11624 25362 11652 29650
rect 11716 28490 11744 30194
rect 11950 29948 12258 29957
rect 11950 29946 11956 29948
rect 12012 29946 12036 29948
rect 12092 29946 12116 29948
rect 12172 29946 12196 29948
rect 12252 29946 12258 29948
rect 12012 29894 12014 29946
rect 12194 29894 12196 29946
rect 11950 29892 11956 29894
rect 12012 29892 12036 29894
rect 12092 29892 12116 29894
rect 12172 29892 12196 29894
rect 12252 29892 12258 29894
rect 11950 29883 12258 29892
rect 11950 28860 12258 28869
rect 11950 28858 11956 28860
rect 12012 28858 12036 28860
rect 12092 28858 12116 28860
rect 12172 28858 12196 28860
rect 12252 28858 12258 28860
rect 12012 28806 12014 28858
rect 12194 28806 12196 28858
rect 11950 28804 11956 28806
rect 12012 28804 12036 28806
rect 12092 28804 12116 28806
rect 12172 28804 12196 28806
rect 12252 28804 12258 28806
rect 11950 28795 12258 28804
rect 11704 28484 11756 28490
rect 11704 28426 11756 28432
rect 11950 27772 12258 27781
rect 11950 27770 11956 27772
rect 12012 27770 12036 27772
rect 12092 27770 12116 27772
rect 12172 27770 12196 27772
rect 12252 27770 12258 27772
rect 12012 27718 12014 27770
rect 12194 27718 12196 27770
rect 11950 27716 11956 27718
rect 12012 27716 12036 27718
rect 12092 27716 12116 27718
rect 12172 27716 12196 27718
rect 12252 27716 12258 27718
rect 11950 27707 12258 27716
rect 12360 27538 12388 31742
rect 12452 29170 12480 31878
rect 12610 31580 12918 31589
rect 12610 31578 12616 31580
rect 12672 31578 12696 31580
rect 12752 31578 12776 31580
rect 12832 31578 12856 31580
rect 12912 31578 12918 31580
rect 12672 31526 12674 31578
rect 12854 31526 12856 31578
rect 12610 31524 12616 31526
rect 12672 31524 12696 31526
rect 12752 31524 12776 31526
rect 12832 31524 12856 31526
rect 12912 31524 12918 31526
rect 12610 31515 12918 31524
rect 14108 30938 14136 63718
rect 14200 41070 14228 67118
rect 14292 45422 14320 67186
rect 15016 67176 15068 67182
rect 15016 67118 15068 67124
rect 15028 64462 15056 67118
rect 15016 64456 15068 64462
rect 15016 64398 15068 64404
rect 14372 63980 14424 63986
rect 14372 63922 14424 63928
rect 14384 50250 14412 63922
rect 14740 54188 14792 54194
rect 14740 54130 14792 54136
rect 14372 50244 14424 50250
rect 14372 50186 14424 50192
rect 14464 49156 14516 49162
rect 14464 49098 14516 49104
rect 14280 45416 14332 45422
rect 14280 45358 14332 45364
rect 14292 44198 14320 45358
rect 14280 44192 14332 44198
rect 14280 44134 14332 44140
rect 14280 41608 14332 41614
rect 14280 41550 14332 41556
rect 14188 41064 14240 41070
rect 14188 41006 14240 41012
rect 14188 39432 14240 39438
rect 14188 39374 14240 39380
rect 14200 39098 14228 39374
rect 14188 39092 14240 39098
rect 14188 39034 14240 39040
rect 14292 37262 14320 41550
rect 14280 37256 14332 37262
rect 14280 37198 14332 37204
rect 14292 35894 14320 37198
rect 14200 35866 14320 35894
rect 14096 30932 14148 30938
rect 14096 30874 14148 30880
rect 12610 30492 12918 30501
rect 12610 30490 12616 30492
rect 12672 30490 12696 30492
rect 12752 30490 12776 30492
rect 12832 30490 12856 30492
rect 12912 30490 12918 30492
rect 12672 30438 12674 30490
rect 12854 30438 12856 30490
rect 12610 30436 12616 30438
rect 12672 30436 12696 30438
rect 12752 30436 12776 30438
rect 12832 30436 12856 30438
rect 12912 30436 12918 30438
rect 12610 30427 12918 30436
rect 14200 29714 14228 35866
rect 14372 33652 14424 33658
rect 14372 33594 14424 33600
rect 14188 29708 14240 29714
rect 14188 29650 14240 29656
rect 14280 29708 14332 29714
rect 14280 29650 14332 29656
rect 13912 29640 13964 29646
rect 13912 29582 13964 29588
rect 12610 29404 12918 29413
rect 12610 29402 12616 29404
rect 12672 29402 12696 29404
rect 12752 29402 12776 29404
rect 12832 29402 12856 29404
rect 12912 29402 12918 29404
rect 12672 29350 12674 29402
rect 12854 29350 12856 29402
rect 12610 29348 12616 29350
rect 12672 29348 12696 29350
rect 12752 29348 12776 29350
rect 12832 29348 12856 29350
rect 12912 29348 12918 29350
rect 12610 29339 12918 29348
rect 12440 29164 12492 29170
rect 12440 29106 12492 29112
rect 12348 27532 12400 27538
rect 12348 27474 12400 27480
rect 12452 27418 12480 29106
rect 12610 28316 12918 28325
rect 12610 28314 12616 28316
rect 12672 28314 12696 28316
rect 12752 28314 12776 28316
rect 12832 28314 12856 28316
rect 12912 28314 12918 28316
rect 12672 28262 12674 28314
rect 12854 28262 12856 28314
rect 12610 28260 12616 28262
rect 12672 28260 12696 28262
rect 12752 28260 12776 28262
rect 12832 28260 12856 28262
rect 12912 28260 12918 28262
rect 12610 28251 12918 28260
rect 12360 27390 12480 27418
rect 11950 26684 12258 26693
rect 11950 26682 11956 26684
rect 12012 26682 12036 26684
rect 12092 26682 12116 26684
rect 12172 26682 12196 26684
rect 12252 26682 12258 26684
rect 12012 26630 12014 26682
rect 12194 26630 12196 26682
rect 11950 26628 11956 26630
rect 12012 26628 12036 26630
rect 12092 26628 12116 26630
rect 12172 26628 12196 26630
rect 12252 26628 12258 26630
rect 11950 26619 12258 26628
rect 11950 25596 12258 25605
rect 11950 25594 11956 25596
rect 12012 25594 12036 25596
rect 12092 25594 12116 25596
rect 12172 25594 12196 25596
rect 12252 25594 12258 25596
rect 12012 25542 12014 25594
rect 12194 25542 12196 25594
rect 11950 25540 11956 25542
rect 12012 25540 12036 25542
rect 12092 25540 12116 25542
rect 12172 25540 12196 25542
rect 12252 25540 12258 25542
rect 11950 25531 12258 25540
rect 11612 25356 11664 25362
rect 11612 25298 11664 25304
rect 11624 22234 11652 25298
rect 11950 24508 12258 24517
rect 11950 24506 11956 24508
rect 12012 24506 12036 24508
rect 12092 24506 12116 24508
rect 12172 24506 12196 24508
rect 12252 24506 12258 24508
rect 12012 24454 12014 24506
rect 12194 24454 12196 24506
rect 11950 24452 11956 24454
rect 12012 24452 12036 24454
rect 12092 24452 12116 24454
rect 12172 24452 12196 24454
rect 12252 24452 12258 24454
rect 11950 24443 12258 24452
rect 11950 23420 12258 23429
rect 11950 23418 11956 23420
rect 12012 23418 12036 23420
rect 12092 23418 12116 23420
rect 12172 23418 12196 23420
rect 12252 23418 12258 23420
rect 12012 23366 12014 23418
rect 12194 23366 12196 23418
rect 11950 23364 11956 23366
rect 12012 23364 12036 23366
rect 12092 23364 12116 23366
rect 12172 23364 12196 23366
rect 12252 23364 12258 23366
rect 11950 23355 12258 23364
rect 11950 22332 12258 22341
rect 11950 22330 11956 22332
rect 12012 22330 12036 22332
rect 12092 22330 12116 22332
rect 12172 22330 12196 22332
rect 12252 22330 12258 22332
rect 12012 22278 12014 22330
rect 12194 22278 12196 22330
rect 11950 22276 11956 22278
rect 12012 22276 12036 22278
rect 12092 22276 12116 22278
rect 12172 22276 12196 22278
rect 12252 22276 12258 22278
rect 11950 22267 12258 22276
rect 11612 22228 11664 22234
rect 11612 22170 11664 22176
rect 11058 21992 11114 22001
rect 11058 21927 11060 21936
rect 11112 21927 11114 21936
rect 11060 21898 11112 21904
rect 11950 21244 12258 21253
rect 11950 21242 11956 21244
rect 12012 21242 12036 21244
rect 12092 21242 12116 21244
rect 12172 21242 12196 21244
rect 12252 21242 12258 21244
rect 12012 21190 12014 21242
rect 12194 21190 12196 21242
rect 11950 21188 11956 21190
rect 12012 21188 12036 21190
rect 12092 21188 12116 21190
rect 12172 21188 12196 21190
rect 12252 21188 12258 21190
rect 11950 21179 12258 21188
rect 11950 20156 12258 20165
rect 11950 20154 11956 20156
rect 12012 20154 12036 20156
rect 12092 20154 12116 20156
rect 12172 20154 12196 20156
rect 12252 20154 12258 20156
rect 12012 20102 12014 20154
rect 12194 20102 12196 20154
rect 11950 20100 11956 20102
rect 12012 20100 12036 20102
rect 12092 20100 12116 20102
rect 12172 20100 12196 20102
rect 12252 20100 12258 20102
rect 11950 20091 12258 20100
rect 11950 19068 12258 19077
rect 11950 19066 11956 19068
rect 12012 19066 12036 19068
rect 12092 19066 12116 19068
rect 12172 19066 12196 19068
rect 12252 19066 12258 19068
rect 12012 19014 12014 19066
rect 12194 19014 12196 19066
rect 11950 19012 11956 19014
rect 12012 19012 12036 19014
rect 12092 19012 12116 19014
rect 12172 19012 12196 19014
rect 12252 19012 12258 19014
rect 11950 19003 12258 19012
rect 11950 17980 12258 17989
rect 11950 17978 11956 17980
rect 12012 17978 12036 17980
rect 12092 17978 12116 17980
rect 12172 17978 12196 17980
rect 12252 17978 12258 17980
rect 12012 17926 12014 17978
rect 12194 17926 12196 17978
rect 11950 17924 11956 17926
rect 12012 17924 12036 17926
rect 12092 17924 12116 17926
rect 12172 17924 12196 17926
rect 12252 17924 12258 17926
rect 11950 17915 12258 17924
rect 11950 16892 12258 16901
rect 11950 16890 11956 16892
rect 12012 16890 12036 16892
rect 12092 16890 12116 16892
rect 12172 16890 12196 16892
rect 12252 16890 12258 16892
rect 12012 16838 12014 16890
rect 12194 16838 12196 16890
rect 11950 16836 11956 16838
rect 12012 16836 12036 16838
rect 12092 16836 12116 16838
rect 12172 16836 12196 16838
rect 12252 16836 12258 16838
rect 11950 16827 12258 16836
rect 11950 15804 12258 15813
rect 11950 15802 11956 15804
rect 12012 15802 12036 15804
rect 12092 15802 12116 15804
rect 12172 15802 12196 15804
rect 12252 15802 12258 15804
rect 12012 15750 12014 15802
rect 12194 15750 12196 15802
rect 11950 15748 11956 15750
rect 12012 15748 12036 15750
rect 12092 15748 12116 15750
rect 12172 15748 12196 15750
rect 12252 15748 12258 15750
rect 11950 15739 12258 15748
rect 11950 14716 12258 14725
rect 11950 14714 11956 14716
rect 12012 14714 12036 14716
rect 12092 14714 12116 14716
rect 12172 14714 12196 14716
rect 12252 14714 12258 14716
rect 12012 14662 12014 14714
rect 12194 14662 12196 14714
rect 11950 14660 11956 14662
rect 12012 14660 12036 14662
rect 12092 14660 12116 14662
rect 12172 14660 12196 14662
rect 12252 14660 12258 14662
rect 11950 14651 12258 14660
rect 11950 13628 12258 13637
rect 11950 13626 11956 13628
rect 12012 13626 12036 13628
rect 12092 13626 12116 13628
rect 12172 13626 12196 13628
rect 12252 13626 12258 13628
rect 12012 13574 12014 13626
rect 12194 13574 12196 13626
rect 11950 13572 11956 13574
rect 12012 13572 12036 13574
rect 12092 13572 12116 13574
rect 12172 13572 12196 13574
rect 12252 13572 12258 13574
rect 11950 13563 12258 13572
rect 11950 12540 12258 12549
rect 11950 12538 11956 12540
rect 12012 12538 12036 12540
rect 12092 12538 12116 12540
rect 12172 12538 12196 12540
rect 12252 12538 12258 12540
rect 12012 12486 12014 12538
rect 12194 12486 12196 12538
rect 11950 12484 11956 12486
rect 12012 12484 12036 12486
rect 12092 12484 12116 12486
rect 12172 12484 12196 12486
rect 12252 12484 12258 12486
rect 11950 12475 12258 12484
rect 11950 11452 12258 11461
rect 11950 11450 11956 11452
rect 12012 11450 12036 11452
rect 12092 11450 12116 11452
rect 12172 11450 12196 11452
rect 12252 11450 12258 11452
rect 12012 11398 12014 11450
rect 12194 11398 12196 11450
rect 11950 11396 11956 11398
rect 12012 11396 12036 11398
rect 12092 11396 12116 11398
rect 12172 11396 12196 11398
rect 12252 11396 12258 11398
rect 11950 11387 12258 11396
rect 11950 10364 12258 10373
rect 11950 10362 11956 10364
rect 12012 10362 12036 10364
rect 12092 10362 12116 10364
rect 12172 10362 12196 10364
rect 12252 10362 12258 10364
rect 12012 10310 12014 10362
rect 12194 10310 12196 10362
rect 11950 10308 11956 10310
rect 12012 10308 12036 10310
rect 12092 10308 12116 10310
rect 12172 10308 12196 10310
rect 12252 10308 12258 10310
rect 11950 10299 12258 10308
rect 10416 9580 10468 9586
rect 10416 9522 10468 9528
rect 11950 9276 12258 9285
rect 11950 9274 11956 9276
rect 12012 9274 12036 9276
rect 12092 9274 12116 9276
rect 12172 9274 12196 9276
rect 12252 9274 12258 9276
rect 12012 9222 12014 9274
rect 12194 9222 12196 9274
rect 11950 9220 11956 9222
rect 12012 9220 12036 9222
rect 12092 9220 12116 9222
rect 12172 9220 12196 9222
rect 12252 9220 12258 9222
rect 11950 9211 12258 9220
rect 11950 8188 12258 8197
rect 11950 8186 11956 8188
rect 12012 8186 12036 8188
rect 12092 8186 12116 8188
rect 12172 8186 12196 8188
rect 12252 8186 12258 8188
rect 12012 8134 12014 8186
rect 12194 8134 12196 8186
rect 11950 8132 11956 8134
rect 12012 8132 12036 8134
rect 12092 8132 12116 8134
rect 12172 8132 12196 8134
rect 12252 8132 12258 8134
rect 11950 8123 12258 8132
rect 11950 7100 12258 7109
rect 11950 7098 11956 7100
rect 12012 7098 12036 7100
rect 12092 7098 12116 7100
rect 12172 7098 12196 7100
rect 12252 7098 12258 7100
rect 12012 7046 12014 7098
rect 12194 7046 12196 7098
rect 11950 7044 11956 7046
rect 12012 7044 12036 7046
rect 12092 7044 12116 7046
rect 12172 7044 12196 7046
rect 12252 7044 12258 7046
rect 11950 7035 12258 7044
rect 11950 6012 12258 6021
rect 11950 6010 11956 6012
rect 12012 6010 12036 6012
rect 12092 6010 12116 6012
rect 12172 6010 12196 6012
rect 12252 6010 12258 6012
rect 12012 5958 12014 6010
rect 12194 5958 12196 6010
rect 11950 5956 11956 5958
rect 12012 5956 12036 5958
rect 12092 5956 12116 5958
rect 12172 5956 12196 5958
rect 12252 5956 12258 5958
rect 11950 5947 12258 5956
rect 11950 4924 12258 4933
rect 11950 4922 11956 4924
rect 12012 4922 12036 4924
rect 12092 4922 12116 4924
rect 12172 4922 12196 4924
rect 12252 4922 12258 4924
rect 12012 4870 12014 4922
rect 12194 4870 12196 4922
rect 11950 4868 11956 4870
rect 12012 4868 12036 4870
rect 12092 4868 12116 4870
rect 12172 4868 12196 4870
rect 12252 4868 12258 4870
rect 11950 4859 12258 4868
rect 12360 3942 12388 27390
rect 12610 27228 12918 27237
rect 12610 27226 12616 27228
rect 12672 27226 12696 27228
rect 12752 27226 12776 27228
rect 12832 27226 12856 27228
rect 12912 27226 12918 27228
rect 12672 27174 12674 27226
rect 12854 27174 12856 27226
rect 12610 27172 12616 27174
rect 12672 27172 12696 27174
rect 12752 27172 12776 27174
rect 12832 27172 12856 27174
rect 12912 27172 12918 27174
rect 12610 27163 12918 27172
rect 12610 26140 12918 26149
rect 12610 26138 12616 26140
rect 12672 26138 12696 26140
rect 12752 26138 12776 26140
rect 12832 26138 12856 26140
rect 12912 26138 12918 26140
rect 12672 26086 12674 26138
rect 12854 26086 12856 26138
rect 12610 26084 12616 26086
rect 12672 26084 12696 26086
rect 12752 26084 12776 26086
rect 12832 26084 12856 26086
rect 12912 26084 12918 26086
rect 12610 26075 12918 26084
rect 12610 25052 12918 25061
rect 12610 25050 12616 25052
rect 12672 25050 12696 25052
rect 12752 25050 12776 25052
rect 12832 25050 12856 25052
rect 12912 25050 12918 25052
rect 12672 24998 12674 25050
rect 12854 24998 12856 25050
rect 12610 24996 12616 24998
rect 12672 24996 12696 24998
rect 12752 24996 12776 24998
rect 12832 24996 12856 24998
rect 12912 24996 12918 24998
rect 12610 24987 12918 24996
rect 12610 23964 12918 23973
rect 12610 23962 12616 23964
rect 12672 23962 12696 23964
rect 12752 23962 12776 23964
rect 12832 23962 12856 23964
rect 12912 23962 12918 23964
rect 12672 23910 12674 23962
rect 12854 23910 12856 23962
rect 12610 23908 12616 23910
rect 12672 23908 12696 23910
rect 12752 23908 12776 23910
rect 12832 23908 12856 23910
rect 12912 23908 12918 23910
rect 12610 23899 12918 23908
rect 12610 22876 12918 22885
rect 12610 22874 12616 22876
rect 12672 22874 12696 22876
rect 12752 22874 12776 22876
rect 12832 22874 12856 22876
rect 12912 22874 12918 22876
rect 12672 22822 12674 22874
rect 12854 22822 12856 22874
rect 12610 22820 12616 22822
rect 12672 22820 12696 22822
rect 12752 22820 12776 22822
rect 12832 22820 12856 22822
rect 12912 22820 12918 22822
rect 12610 22811 12918 22820
rect 12610 21788 12918 21797
rect 12610 21786 12616 21788
rect 12672 21786 12696 21788
rect 12752 21786 12776 21788
rect 12832 21786 12856 21788
rect 12912 21786 12918 21788
rect 12672 21734 12674 21786
rect 12854 21734 12856 21786
rect 12610 21732 12616 21734
rect 12672 21732 12696 21734
rect 12752 21732 12776 21734
rect 12832 21732 12856 21734
rect 12912 21732 12918 21734
rect 12610 21723 12918 21732
rect 12610 20700 12918 20709
rect 12610 20698 12616 20700
rect 12672 20698 12696 20700
rect 12752 20698 12776 20700
rect 12832 20698 12856 20700
rect 12912 20698 12918 20700
rect 12672 20646 12674 20698
rect 12854 20646 12856 20698
rect 12610 20644 12616 20646
rect 12672 20644 12696 20646
rect 12752 20644 12776 20646
rect 12832 20644 12856 20646
rect 12912 20644 12918 20646
rect 12610 20635 12918 20644
rect 12610 19612 12918 19621
rect 12610 19610 12616 19612
rect 12672 19610 12696 19612
rect 12752 19610 12776 19612
rect 12832 19610 12856 19612
rect 12912 19610 12918 19612
rect 12672 19558 12674 19610
rect 12854 19558 12856 19610
rect 12610 19556 12616 19558
rect 12672 19556 12696 19558
rect 12752 19556 12776 19558
rect 12832 19556 12856 19558
rect 12912 19556 12918 19558
rect 12610 19547 12918 19556
rect 12610 18524 12918 18533
rect 12610 18522 12616 18524
rect 12672 18522 12696 18524
rect 12752 18522 12776 18524
rect 12832 18522 12856 18524
rect 12912 18522 12918 18524
rect 12672 18470 12674 18522
rect 12854 18470 12856 18522
rect 12610 18468 12616 18470
rect 12672 18468 12696 18470
rect 12752 18468 12776 18470
rect 12832 18468 12856 18470
rect 12912 18468 12918 18470
rect 12610 18459 12918 18468
rect 12610 17436 12918 17445
rect 12610 17434 12616 17436
rect 12672 17434 12696 17436
rect 12752 17434 12776 17436
rect 12832 17434 12856 17436
rect 12912 17434 12918 17436
rect 12672 17382 12674 17434
rect 12854 17382 12856 17434
rect 12610 17380 12616 17382
rect 12672 17380 12696 17382
rect 12752 17380 12776 17382
rect 12832 17380 12856 17382
rect 12912 17380 12918 17382
rect 12610 17371 12918 17380
rect 12610 16348 12918 16357
rect 12610 16346 12616 16348
rect 12672 16346 12696 16348
rect 12752 16346 12776 16348
rect 12832 16346 12856 16348
rect 12912 16346 12918 16348
rect 12672 16294 12674 16346
rect 12854 16294 12856 16346
rect 12610 16292 12616 16294
rect 12672 16292 12696 16294
rect 12752 16292 12776 16294
rect 12832 16292 12856 16294
rect 12912 16292 12918 16294
rect 12610 16283 12918 16292
rect 12610 15260 12918 15269
rect 12610 15258 12616 15260
rect 12672 15258 12696 15260
rect 12752 15258 12776 15260
rect 12832 15258 12856 15260
rect 12912 15258 12918 15260
rect 12672 15206 12674 15258
rect 12854 15206 12856 15258
rect 12610 15204 12616 15206
rect 12672 15204 12696 15206
rect 12752 15204 12776 15206
rect 12832 15204 12856 15206
rect 12912 15204 12918 15206
rect 12610 15195 12918 15204
rect 12610 14172 12918 14181
rect 12610 14170 12616 14172
rect 12672 14170 12696 14172
rect 12752 14170 12776 14172
rect 12832 14170 12856 14172
rect 12912 14170 12918 14172
rect 12672 14118 12674 14170
rect 12854 14118 12856 14170
rect 12610 14116 12616 14118
rect 12672 14116 12696 14118
rect 12752 14116 12776 14118
rect 12832 14116 12856 14118
rect 12912 14116 12918 14118
rect 12610 14107 12918 14116
rect 13636 13728 13688 13734
rect 13636 13670 13688 13676
rect 12610 13084 12918 13093
rect 12610 13082 12616 13084
rect 12672 13082 12696 13084
rect 12752 13082 12776 13084
rect 12832 13082 12856 13084
rect 12912 13082 12918 13084
rect 12672 13030 12674 13082
rect 12854 13030 12856 13082
rect 12610 13028 12616 13030
rect 12672 13028 12696 13030
rect 12752 13028 12776 13030
rect 12832 13028 12856 13030
rect 12912 13028 12918 13030
rect 12610 13019 12918 13028
rect 12610 11996 12918 12005
rect 12610 11994 12616 11996
rect 12672 11994 12696 11996
rect 12752 11994 12776 11996
rect 12832 11994 12856 11996
rect 12912 11994 12918 11996
rect 12672 11942 12674 11994
rect 12854 11942 12856 11994
rect 12610 11940 12616 11942
rect 12672 11940 12696 11942
rect 12752 11940 12776 11942
rect 12832 11940 12856 11942
rect 12912 11940 12918 11942
rect 12610 11931 12918 11940
rect 12610 10908 12918 10917
rect 12610 10906 12616 10908
rect 12672 10906 12696 10908
rect 12752 10906 12776 10908
rect 12832 10906 12856 10908
rect 12912 10906 12918 10908
rect 12672 10854 12674 10906
rect 12854 10854 12856 10906
rect 12610 10852 12616 10854
rect 12672 10852 12696 10854
rect 12752 10852 12776 10854
rect 12832 10852 12856 10854
rect 12912 10852 12918 10854
rect 12610 10843 12918 10852
rect 12610 9820 12918 9829
rect 12610 9818 12616 9820
rect 12672 9818 12696 9820
rect 12752 9818 12776 9820
rect 12832 9818 12856 9820
rect 12912 9818 12918 9820
rect 12672 9766 12674 9818
rect 12854 9766 12856 9818
rect 12610 9764 12616 9766
rect 12672 9764 12696 9766
rect 12752 9764 12776 9766
rect 12832 9764 12856 9766
rect 12912 9764 12918 9766
rect 12610 9755 12918 9764
rect 12610 8732 12918 8741
rect 12610 8730 12616 8732
rect 12672 8730 12696 8732
rect 12752 8730 12776 8732
rect 12832 8730 12856 8732
rect 12912 8730 12918 8732
rect 12672 8678 12674 8730
rect 12854 8678 12856 8730
rect 12610 8676 12616 8678
rect 12672 8676 12696 8678
rect 12752 8676 12776 8678
rect 12832 8676 12856 8678
rect 12912 8676 12918 8678
rect 12610 8667 12918 8676
rect 13648 8090 13676 13670
rect 13728 9580 13780 9586
rect 13728 9522 13780 9528
rect 13636 8084 13688 8090
rect 13636 8026 13688 8032
rect 13740 7886 13768 9522
rect 13728 7880 13780 7886
rect 13728 7822 13780 7828
rect 12610 7644 12918 7653
rect 12610 7642 12616 7644
rect 12672 7642 12696 7644
rect 12752 7642 12776 7644
rect 12832 7642 12856 7644
rect 12912 7642 12918 7644
rect 12672 7590 12674 7642
rect 12854 7590 12856 7642
rect 12610 7588 12616 7590
rect 12672 7588 12696 7590
rect 12752 7588 12776 7590
rect 12832 7588 12856 7590
rect 12912 7588 12918 7590
rect 12610 7579 12918 7588
rect 12610 6556 12918 6565
rect 12610 6554 12616 6556
rect 12672 6554 12696 6556
rect 12752 6554 12776 6556
rect 12832 6554 12856 6556
rect 12912 6554 12918 6556
rect 12672 6502 12674 6554
rect 12854 6502 12856 6554
rect 12610 6500 12616 6502
rect 12672 6500 12696 6502
rect 12752 6500 12776 6502
rect 12832 6500 12856 6502
rect 12912 6500 12918 6502
rect 12610 6491 12918 6500
rect 12610 5468 12918 5477
rect 12610 5466 12616 5468
rect 12672 5466 12696 5468
rect 12752 5466 12776 5468
rect 12832 5466 12856 5468
rect 12912 5466 12918 5468
rect 12672 5414 12674 5466
rect 12854 5414 12856 5466
rect 12610 5412 12616 5414
rect 12672 5412 12696 5414
rect 12752 5412 12776 5414
rect 12832 5412 12856 5414
rect 12912 5412 12918 5414
rect 12610 5403 12918 5412
rect 12610 4380 12918 4389
rect 12610 4378 12616 4380
rect 12672 4378 12696 4380
rect 12752 4378 12776 4380
rect 12832 4378 12856 4380
rect 12912 4378 12918 4380
rect 12672 4326 12674 4378
rect 12854 4326 12856 4378
rect 12610 4324 12616 4326
rect 12672 4324 12696 4326
rect 12752 4324 12776 4326
rect 12832 4324 12856 4326
rect 12912 4324 12918 4326
rect 12610 4315 12918 4324
rect 12348 3936 12400 3942
rect 12348 3878 12400 3884
rect 11950 3836 12258 3845
rect 11950 3834 11956 3836
rect 12012 3834 12036 3836
rect 12092 3834 12116 3836
rect 12172 3834 12196 3836
rect 12252 3834 12258 3836
rect 12012 3782 12014 3834
rect 12194 3782 12196 3834
rect 11950 3780 11956 3782
rect 12012 3780 12036 3782
rect 12092 3780 12116 3782
rect 12172 3780 12196 3782
rect 12252 3780 12258 3782
rect 11950 3771 12258 3780
rect 13924 3670 13952 29582
rect 14096 25356 14148 25362
rect 14096 25298 14148 25304
rect 14108 15502 14136 25298
rect 14200 23118 14228 29650
rect 14292 27130 14320 29650
rect 14384 28994 14412 33594
rect 14476 29238 14504 49098
rect 14554 45928 14610 45937
rect 14554 45863 14556 45872
rect 14608 45863 14610 45872
rect 14556 45834 14608 45840
rect 14648 44192 14700 44198
rect 14648 44134 14700 44140
rect 14660 31482 14688 44134
rect 14648 31476 14700 31482
rect 14648 31418 14700 31424
rect 14556 30864 14608 30870
rect 14556 30806 14608 30812
rect 14464 29232 14516 29238
rect 14464 29174 14516 29180
rect 14384 28966 14504 28994
rect 14280 27124 14332 27130
rect 14280 27066 14332 27072
rect 14280 24132 14332 24138
rect 14280 24074 14332 24080
rect 14188 23112 14240 23118
rect 14188 23054 14240 23060
rect 14292 16658 14320 24074
rect 14476 19334 14504 28966
rect 14568 24138 14596 30806
rect 14556 24132 14608 24138
rect 14556 24074 14608 24080
rect 14384 19306 14504 19334
rect 14280 16652 14332 16658
rect 14280 16594 14332 16600
rect 14384 15502 14412 19306
rect 14752 16590 14780 54130
rect 14832 50244 14884 50250
rect 14832 50186 14884 50192
rect 14844 45558 14872 50186
rect 15028 49162 15056 64398
rect 15108 49836 15160 49842
rect 15108 49778 15160 49784
rect 15016 49156 15068 49162
rect 15016 49098 15068 49104
rect 14832 45552 14884 45558
rect 14832 45494 14884 45500
rect 14924 41608 14976 41614
rect 14924 41550 14976 41556
rect 14832 33924 14884 33930
rect 14832 33866 14884 33872
rect 14844 25362 14872 33866
rect 14936 33522 14964 41550
rect 15120 33930 15148 49778
rect 15108 33924 15160 33930
rect 15108 33866 15160 33872
rect 14924 33516 14976 33522
rect 14924 33458 14976 33464
rect 14832 25356 14884 25362
rect 14832 25298 14884 25304
rect 14740 16584 14792 16590
rect 14740 16526 14792 16532
rect 15016 16584 15068 16590
rect 15016 16526 15068 16532
rect 15028 16250 15056 16526
rect 15016 16244 15068 16250
rect 15016 16186 15068 16192
rect 14096 15496 14148 15502
rect 14096 15438 14148 15444
rect 14372 15496 14424 15502
rect 14372 15438 14424 15444
rect 14108 8838 14136 15438
rect 14188 15360 14240 15366
rect 14188 15302 14240 15308
rect 14096 8832 14148 8838
rect 14096 8774 14148 8780
rect 13912 3664 13964 3670
rect 13912 3606 13964 3612
rect 12610 3292 12918 3301
rect 12610 3290 12616 3292
rect 12672 3290 12696 3292
rect 12752 3290 12776 3292
rect 12832 3290 12856 3292
rect 12912 3290 12918 3292
rect 12672 3238 12674 3290
rect 12854 3238 12856 3290
rect 12610 3236 12616 3238
rect 12672 3236 12696 3238
rect 12752 3236 12776 3238
rect 12832 3236 12856 3238
rect 12912 3236 12918 3238
rect 12610 3227 12918 3236
rect 14108 3058 14136 8774
rect 14096 3052 14148 3058
rect 14096 2994 14148 3000
rect 14200 2990 14228 15302
rect 14280 4004 14332 4010
rect 14280 3946 14332 3952
rect 14292 3058 14320 3946
rect 14384 3398 14412 15438
rect 14372 3392 14424 3398
rect 14372 3334 14424 3340
rect 14280 3052 14332 3058
rect 14280 2994 14332 3000
rect 14188 2984 14240 2990
rect 14188 2926 14240 2932
rect 14292 2854 14320 2994
rect 14280 2848 14332 2854
rect 14280 2790 14332 2796
rect 11950 2748 12258 2757
rect 11950 2746 11956 2748
rect 12012 2746 12036 2748
rect 12092 2746 12116 2748
rect 12172 2746 12196 2748
rect 12252 2746 12258 2748
rect 12012 2694 12014 2746
rect 12194 2694 12196 2746
rect 11950 2692 11956 2694
rect 12012 2692 12036 2694
rect 12092 2692 12116 2694
rect 12172 2692 12196 2694
rect 12252 2692 12258 2694
rect 11950 2683 12258 2692
rect 15212 2582 15240 69362
rect 16950 69116 17258 69125
rect 16950 69114 16956 69116
rect 17012 69114 17036 69116
rect 17092 69114 17116 69116
rect 17172 69114 17196 69116
rect 17252 69114 17258 69116
rect 17012 69062 17014 69114
rect 17194 69062 17196 69114
rect 16950 69060 16956 69062
rect 17012 69060 17036 69062
rect 17092 69060 17116 69062
rect 17172 69060 17196 69062
rect 17252 69060 17258 69062
rect 16950 69051 17258 69060
rect 16488 68740 16540 68746
rect 16488 68682 16540 68688
rect 16500 64394 16528 68682
rect 16672 68672 16724 68678
rect 16672 68614 16724 68620
rect 16684 64462 16712 68614
rect 17610 68572 17918 68581
rect 17610 68570 17616 68572
rect 17672 68570 17696 68572
rect 17752 68570 17776 68572
rect 17832 68570 17856 68572
rect 17912 68570 17918 68572
rect 17672 68518 17674 68570
rect 17854 68518 17856 68570
rect 17610 68516 17616 68518
rect 17672 68516 17696 68518
rect 17752 68516 17776 68518
rect 17832 68516 17856 68518
rect 17912 68516 17918 68518
rect 17610 68507 17918 68516
rect 18696 68400 18748 68406
rect 18696 68342 18748 68348
rect 16950 68028 17258 68037
rect 16950 68026 16956 68028
rect 17012 68026 17036 68028
rect 17092 68026 17116 68028
rect 17172 68026 17196 68028
rect 17252 68026 17258 68028
rect 17012 67974 17014 68026
rect 17194 67974 17196 68026
rect 16950 67972 16956 67974
rect 17012 67972 17036 67974
rect 17092 67972 17116 67974
rect 17172 67972 17196 67974
rect 17252 67972 17258 67974
rect 16950 67963 17258 67972
rect 17610 67484 17918 67493
rect 17610 67482 17616 67484
rect 17672 67482 17696 67484
rect 17752 67482 17776 67484
rect 17832 67482 17856 67484
rect 17912 67482 17918 67484
rect 17672 67430 17674 67482
rect 17854 67430 17856 67482
rect 17610 67428 17616 67430
rect 17672 67428 17696 67430
rect 17752 67428 17776 67430
rect 17832 67428 17856 67430
rect 17912 67428 17918 67430
rect 17610 67419 17918 67428
rect 17316 67176 17368 67182
rect 17316 67118 17368 67124
rect 16950 66940 17258 66949
rect 16950 66938 16956 66940
rect 17012 66938 17036 66940
rect 17092 66938 17116 66940
rect 17172 66938 17196 66940
rect 17252 66938 17258 66940
rect 17012 66886 17014 66938
rect 17194 66886 17196 66938
rect 16950 66884 16956 66886
rect 17012 66884 17036 66886
rect 17092 66884 17116 66886
rect 17172 66884 17196 66886
rect 17252 66884 17258 66886
rect 16950 66875 17258 66884
rect 16950 65852 17258 65861
rect 16950 65850 16956 65852
rect 17012 65850 17036 65852
rect 17092 65850 17116 65852
rect 17172 65850 17196 65852
rect 17252 65850 17258 65852
rect 17012 65798 17014 65850
rect 17194 65798 17196 65850
rect 16950 65796 16956 65798
rect 17012 65796 17036 65798
rect 17092 65796 17116 65798
rect 17172 65796 17196 65798
rect 17252 65796 17258 65798
rect 16950 65787 17258 65796
rect 16950 64764 17258 64773
rect 16950 64762 16956 64764
rect 17012 64762 17036 64764
rect 17092 64762 17116 64764
rect 17172 64762 17196 64764
rect 17252 64762 17258 64764
rect 17012 64710 17014 64762
rect 17194 64710 17196 64762
rect 16950 64708 16956 64710
rect 17012 64708 17036 64710
rect 17092 64708 17116 64710
rect 17172 64708 17196 64710
rect 17252 64708 17258 64710
rect 16950 64699 17258 64708
rect 16672 64456 16724 64462
rect 16672 64398 16724 64404
rect 16488 64388 16540 64394
rect 16488 64330 16540 64336
rect 15660 63980 15712 63986
rect 15660 63922 15712 63928
rect 15292 63776 15344 63782
rect 15292 63718 15344 63724
rect 15304 29646 15332 63718
rect 15384 45892 15436 45898
rect 15384 45834 15436 45840
rect 15396 41614 15424 45834
rect 15384 41608 15436 41614
rect 15384 41550 15436 41556
rect 15568 41472 15620 41478
rect 15568 41414 15620 41420
rect 15476 34604 15528 34610
rect 15476 34546 15528 34552
rect 15384 32768 15436 32774
rect 15384 32710 15436 32716
rect 15292 29640 15344 29646
rect 15292 29582 15344 29588
rect 15396 29306 15424 32710
rect 15384 29300 15436 29306
rect 15384 29242 15436 29248
rect 15488 16590 15516 34546
rect 15580 24410 15608 41414
rect 15568 24404 15620 24410
rect 15568 24346 15620 24352
rect 15672 17066 15700 63922
rect 15936 52488 15988 52494
rect 15936 52430 15988 52436
rect 15948 48074 15976 52430
rect 15936 48068 15988 48074
rect 15936 48010 15988 48016
rect 15844 40452 15896 40458
rect 15844 40394 15896 40400
rect 15856 27402 15884 40394
rect 15948 35494 15976 48010
rect 16120 41268 16172 41274
rect 16120 41210 16172 41216
rect 16132 40458 16160 41210
rect 16120 40452 16172 40458
rect 16120 40394 16172 40400
rect 15936 35488 15988 35494
rect 15936 35430 15988 35436
rect 15948 34610 15976 35430
rect 15936 34604 15988 34610
rect 15936 34546 15988 34552
rect 16500 32774 16528 64330
rect 16580 64320 16632 64326
rect 16580 64262 16632 64268
rect 16592 64122 16620 64262
rect 16580 64116 16632 64122
rect 16580 64058 16632 64064
rect 16580 51400 16632 51406
rect 16580 51342 16632 51348
rect 16488 32768 16540 32774
rect 16488 32710 16540 32716
rect 16592 31142 16620 51342
rect 16684 41274 16712 64398
rect 16764 64320 16816 64326
rect 16764 64262 16816 64268
rect 16672 41268 16724 41274
rect 16672 41210 16724 41216
rect 16776 40526 16804 64262
rect 16950 63676 17258 63685
rect 16950 63674 16956 63676
rect 17012 63674 17036 63676
rect 17092 63674 17116 63676
rect 17172 63674 17196 63676
rect 17252 63674 17258 63676
rect 17012 63622 17014 63674
rect 17194 63622 17196 63674
rect 16950 63620 16956 63622
rect 17012 63620 17036 63622
rect 17092 63620 17116 63622
rect 17172 63620 17196 63622
rect 17252 63620 17258 63622
rect 16950 63611 17258 63620
rect 16950 62588 17258 62597
rect 16950 62586 16956 62588
rect 17012 62586 17036 62588
rect 17092 62586 17116 62588
rect 17172 62586 17196 62588
rect 17252 62586 17258 62588
rect 17012 62534 17014 62586
rect 17194 62534 17196 62586
rect 16950 62532 16956 62534
rect 17012 62532 17036 62534
rect 17092 62532 17116 62534
rect 17172 62532 17196 62534
rect 17252 62532 17258 62534
rect 16950 62523 17258 62532
rect 16950 61500 17258 61509
rect 16950 61498 16956 61500
rect 17012 61498 17036 61500
rect 17092 61498 17116 61500
rect 17172 61498 17196 61500
rect 17252 61498 17258 61500
rect 17012 61446 17014 61498
rect 17194 61446 17196 61498
rect 16950 61444 16956 61446
rect 17012 61444 17036 61446
rect 17092 61444 17116 61446
rect 17172 61444 17196 61446
rect 17252 61444 17258 61446
rect 16950 61435 17258 61444
rect 16950 60412 17258 60421
rect 16950 60410 16956 60412
rect 17012 60410 17036 60412
rect 17092 60410 17116 60412
rect 17172 60410 17196 60412
rect 17252 60410 17258 60412
rect 17012 60358 17014 60410
rect 17194 60358 17196 60410
rect 16950 60356 16956 60358
rect 17012 60356 17036 60358
rect 17092 60356 17116 60358
rect 17172 60356 17196 60358
rect 17252 60356 17258 60358
rect 16950 60347 17258 60356
rect 16950 59324 17258 59333
rect 16950 59322 16956 59324
rect 17012 59322 17036 59324
rect 17092 59322 17116 59324
rect 17172 59322 17196 59324
rect 17252 59322 17258 59324
rect 17012 59270 17014 59322
rect 17194 59270 17196 59322
rect 16950 59268 16956 59270
rect 17012 59268 17036 59270
rect 17092 59268 17116 59270
rect 17172 59268 17196 59270
rect 17252 59268 17258 59270
rect 16950 59259 17258 59268
rect 16950 58236 17258 58245
rect 16950 58234 16956 58236
rect 17012 58234 17036 58236
rect 17092 58234 17116 58236
rect 17172 58234 17196 58236
rect 17252 58234 17258 58236
rect 17012 58182 17014 58234
rect 17194 58182 17196 58234
rect 16950 58180 16956 58182
rect 17012 58180 17036 58182
rect 17092 58180 17116 58182
rect 17172 58180 17196 58182
rect 17252 58180 17258 58182
rect 16950 58171 17258 58180
rect 16950 57148 17258 57157
rect 16950 57146 16956 57148
rect 17012 57146 17036 57148
rect 17092 57146 17116 57148
rect 17172 57146 17196 57148
rect 17252 57146 17258 57148
rect 17012 57094 17014 57146
rect 17194 57094 17196 57146
rect 16950 57092 16956 57094
rect 17012 57092 17036 57094
rect 17092 57092 17116 57094
rect 17172 57092 17196 57094
rect 17252 57092 17258 57094
rect 16950 57083 17258 57092
rect 16950 56060 17258 56069
rect 16950 56058 16956 56060
rect 17012 56058 17036 56060
rect 17092 56058 17116 56060
rect 17172 56058 17196 56060
rect 17252 56058 17258 56060
rect 17012 56006 17014 56058
rect 17194 56006 17196 56058
rect 16950 56004 16956 56006
rect 17012 56004 17036 56006
rect 17092 56004 17116 56006
rect 17172 56004 17196 56006
rect 17252 56004 17258 56006
rect 16950 55995 17258 56004
rect 16856 55344 16908 55350
rect 16856 55286 16908 55292
rect 16868 51406 16896 55286
rect 16950 54972 17258 54981
rect 16950 54970 16956 54972
rect 17012 54970 17036 54972
rect 17092 54970 17116 54972
rect 17172 54970 17196 54972
rect 17252 54970 17258 54972
rect 17012 54918 17014 54970
rect 17194 54918 17196 54970
rect 16950 54916 16956 54918
rect 17012 54916 17036 54918
rect 17092 54916 17116 54918
rect 17172 54916 17196 54918
rect 17252 54916 17258 54918
rect 16950 54907 17258 54916
rect 16950 53884 17258 53893
rect 16950 53882 16956 53884
rect 17012 53882 17036 53884
rect 17092 53882 17116 53884
rect 17172 53882 17196 53884
rect 17252 53882 17258 53884
rect 17012 53830 17014 53882
rect 17194 53830 17196 53882
rect 16950 53828 16956 53830
rect 17012 53828 17036 53830
rect 17092 53828 17116 53830
rect 17172 53828 17196 53830
rect 17252 53828 17258 53830
rect 16950 53819 17258 53828
rect 17328 53446 17356 67118
rect 17610 66396 17918 66405
rect 17610 66394 17616 66396
rect 17672 66394 17696 66396
rect 17752 66394 17776 66396
rect 17832 66394 17856 66396
rect 17912 66394 17918 66396
rect 17672 66342 17674 66394
rect 17854 66342 17856 66394
rect 17610 66340 17616 66342
rect 17672 66340 17696 66342
rect 17752 66340 17776 66342
rect 17832 66340 17856 66342
rect 17912 66340 17918 66342
rect 17610 66331 17918 66340
rect 17610 65308 17918 65317
rect 17610 65306 17616 65308
rect 17672 65306 17696 65308
rect 17752 65306 17776 65308
rect 17832 65306 17856 65308
rect 17912 65306 17918 65308
rect 17672 65254 17674 65306
rect 17854 65254 17856 65306
rect 17610 65252 17616 65254
rect 17672 65252 17696 65254
rect 17752 65252 17776 65254
rect 17832 65252 17856 65254
rect 17912 65252 17918 65254
rect 17610 65243 17918 65252
rect 17408 65136 17460 65142
rect 17408 65078 17460 65084
rect 17420 63510 17448 65078
rect 17500 64524 17552 64530
rect 17500 64466 17552 64472
rect 17408 63504 17460 63510
rect 17408 63446 17460 63452
rect 17408 54052 17460 54058
rect 17408 53994 17460 54000
rect 17316 53440 17368 53446
rect 17316 53382 17368 53388
rect 16950 52796 17258 52805
rect 16950 52794 16956 52796
rect 17012 52794 17036 52796
rect 17092 52794 17116 52796
rect 17172 52794 17196 52796
rect 17252 52794 17258 52796
rect 17012 52742 17014 52794
rect 17194 52742 17196 52794
rect 16950 52740 16956 52742
rect 17012 52740 17036 52742
rect 17092 52740 17116 52742
rect 17172 52740 17196 52742
rect 17252 52740 17258 52742
rect 16950 52731 17258 52740
rect 16950 51708 17258 51717
rect 16950 51706 16956 51708
rect 17012 51706 17036 51708
rect 17092 51706 17116 51708
rect 17172 51706 17196 51708
rect 17252 51706 17258 51708
rect 17012 51654 17014 51706
rect 17194 51654 17196 51706
rect 16950 51652 16956 51654
rect 17012 51652 17036 51654
rect 17092 51652 17116 51654
rect 17172 51652 17196 51654
rect 17252 51652 17258 51654
rect 16950 51643 17258 51652
rect 17328 51406 17356 53382
rect 16856 51400 16908 51406
rect 16856 51342 16908 51348
rect 17316 51400 17368 51406
rect 17316 51342 17368 51348
rect 16868 45490 16896 51342
rect 16950 50620 17258 50629
rect 16950 50618 16956 50620
rect 17012 50618 17036 50620
rect 17092 50618 17116 50620
rect 17172 50618 17196 50620
rect 17252 50618 17258 50620
rect 17012 50566 17014 50618
rect 17194 50566 17196 50618
rect 16950 50564 16956 50566
rect 17012 50564 17036 50566
rect 17092 50564 17116 50566
rect 17172 50564 17196 50566
rect 17252 50564 17258 50566
rect 16950 50555 17258 50564
rect 16950 49532 17258 49541
rect 16950 49530 16956 49532
rect 17012 49530 17036 49532
rect 17092 49530 17116 49532
rect 17172 49530 17196 49532
rect 17252 49530 17258 49532
rect 17012 49478 17014 49530
rect 17194 49478 17196 49530
rect 16950 49476 16956 49478
rect 17012 49476 17036 49478
rect 17092 49476 17116 49478
rect 17172 49476 17196 49478
rect 17252 49476 17258 49478
rect 16950 49467 17258 49476
rect 16950 48444 17258 48453
rect 16950 48442 16956 48444
rect 17012 48442 17036 48444
rect 17092 48442 17116 48444
rect 17172 48442 17196 48444
rect 17252 48442 17258 48444
rect 17012 48390 17014 48442
rect 17194 48390 17196 48442
rect 16950 48388 16956 48390
rect 17012 48388 17036 48390
rect 17092 48388 17116 48390
rect 17172 48388 17196 48390
rect 17252 48388 17258 48390
rect 16950 48379 17258 48388
rect 16950 47356 17258 47365
rect 16950 47354 16956 47356
rect 17012 47354 17036 47356
rect 17092 47354 17116 47356
rect 17172 47354 17196 47356
rect 17252 47354 17258 47356
rect 17012 47302 17014 47354
rect 17194 47302 17196 47354
rect 16950 47300 16956 47302
rect 17012 47300 17036 47302
rect 17092 47300 17116 47302
rect 17172 47300 17196 47302
rect 17252 47300 17258 47302
rect 16950 47291 17258 47300
rect 16950 46268 17258 46277
rect 16950 46266 16956 46268
rect 17012 46266 17036 46268
rect 17092 46266 17116 46268
rect 17172 46266 17196 46268
rect 17252 46266 17258 46268
rect 17012 46214 17014 46266
rect 17194 46214 17196 46266
rect 16950 46212 16956 46214
rect 17012 46212 17036 46214
rect 17092 46212 17116 46214
rect 17172 46212 17196 46214
rect 17252 46212 17258 46214
rect 16950 46203 17258 46212
rect 16856 45484 16908 45490
rect 16856 45426 16908 45432
rect 16868 44198 16896 45426
rect 16950 45180 17258 45189
rect 16950 45178 16956 45180
rect 17012 45178 17036 45180
rect 17092 45178 17116 45180
rect 17172 45178 17196 45180
rect 17252 45178 17258 45180
rect 17012 45126 17014 45178
rect 17194 45126 17196 45178
rect 16950 45124 16956 45126
rect 17012 45124 17036 45126
rect 17092 45124 17116 45126
rect 17172 45124 17196 45126
rect 17252 45124 17258 45126
rect 16950 45115 17258 45124
rect 16856 44192 16908 44198
rect 16856 44134 16908 44140
rect 17316 44192 17368 44198
rect 17316 44134 17368 44140
rect 16950 44092 17258 44101
rect 16950 44090 16956 44092
rect 17012 44090 17036 44092
rect 17092 44090 17116 44092
rect 17172 44090 17196 44092
rect 17252 44090 17258 44092
rect 17012 44038 17014 44090
rect 17194 44038 17196 44090
rect 16950 44036 16956 44038
rect 17012 44036 17036 44038
rect 17092 44036 17116 44038
rect 17172 44036 17196 44038
rect 17252 44036 17258 44038
rect 16950 44027 17258 44036
rect 16950 43004 17258 43013
rect 16950 43002 16956 43004
rect 17012 43002 17036 43004
rect 17092 43002 17116 43004
rect 17172 43002 17196 43004
rect 17252 43002 17258 43004
rect 17012 42950 17014 43002
rect 17194 42950 17196 43002
rect 16950 42948 16956 42950
rect 17012 42948 17036 42950
rect 17092 42948 17116 42950
rect 17172 42948 17196 42950
rect 17252 42948 17258 42950
rect 16950 42939 17258 42948
rect 16950 41916 17258 41925
rect 16950 41914 16956 41916
rect 17012 41914 17036 41916
rect 17092 41914 17116 41916
rect 17172 41914 17196 41916
rect 17252 41914 17258 41916
rect 17012 41862 17014 41914
rect 17194 41862 17196 41914
rect 16950 41860 16956 41862
rect 17012 41860 17036 41862
rect 17092 41860 17116 41862
rect 17172 41860 17196 41862
rect 17252 41860 17258 41862
rect 16950 41851 17258 41860
rect 16950 40828 17258 40837
rect 16950 40826 16956 40828
rect 17012 40826 17036 40828
rect 17092 40826 17116 40828
rect 17172 40826 17196 40828
rect 17252 40826 17258 40828
rect 17012 40774 17014 40826
rect 17194 40774 17196 40826
rect 16950 40772 16956 40774
rect 17012 40772 17036 40774
rect 17092 40772 17116 40774
rect 17172 40772 17196 40774
rect 17252 40772 17258 40774
rect 16950 40763 17258 40772
rect 16764 40520 16816 40526
rect 16764 40462 16816 40468
rect 16950 39740 17258 39749
rect 16950 39738 16956 39740
rect 17012 39738 17036 39740
rect 17092 39738 17116 39740
rect 17172 39738 17196 39740
rect 17252 39738 17258 39740
rect 17012 39686 17014 39738
rect 17194 39686 17196 39738
rect 16950 39684 16956 39686
rect 17012 39684 17036 39686
rect 17092 39684 17116 39686
rect 17172 39684 17196 39686
rect 17252 39684 17258 39686
rect 16950 39675 17258 39684
rect 16950 38652 17258 38661
rect 16950 38650 16956 38652
rect 17012 38650 17036 38652
rect 17092 38650 17116 38652
rect 17172 38650 17196 38652
rect 17252 38650 17258 38652
rect 17012 38598 17014 38650
rect 17194 38598 17196 38650
rect 16950 38596 16956 38598
rect 17012 38596 17036 38598
rect 17092 38596 17116 38598
rect 17172 38596 17196 38598
rect 17252 38596 17258 38598
rect 16950 38587 17258 38596
rect 16950 37564 17258 37573
rect 16950 37562 16956 37564
rect 17012 37562 17036 37564
rect 17092 37562 17116 37564
rect 17172 37562 17196 37564
rect 17252 37562 17258 37564
rect 17012 37510 17014 37562
rect 17194 37510 17196 37562
rect 16950 37508 16956 37510
rect 17012 37508 17036 37510
rect 17092 37508 17116 37510
rect 17172 37508 17196 37510
rect 17252 37508 17258 37510
rect 16950 37499 17258 37508
rect 16950 36476 17258 36485
rect 16950 36474 16956 36476
rect 17012 36474 17036 36476
rect 17092 36474 17116 36476
rect 17172 36474 17196 36476
rect 17252 36474 17258 36476
rect 17012 36422 17014 36474
rect 17194 36422 17196 36474
rect 16950 36420 16956 36422
rect 17012 36420 17036 36422
rect 17092 36420 17116 36422
rect 17172 36420 17196 36422
rect 17252 36420 17258 36422
rect 16950 36411 17258 36420
rect 16950 35388 17258 35397
rect 16950 35386 16956 35388
rect 17012 35386 17036 35388
rect 17092 35386 17116 35388
rect 17172 35386 17196 35388
rect 17252 35386 17258 35388
rect 17012 35334 17014 35386
rect 17194 35334 17196 35386
rect 16950 35332 16956 35334
rect 17012 35332 17036 35334
rect 17092 35332 17116 35334
rect 17172 35332 17196 35334
rect 17252 35332 17258 35334
rect 16950 35323 17258 35332
rect 16950 34300 17258 34309
rect 16950 34298 16956 34300
rect 17012 34298 17036 34300
rect 17092 34298 17116 34300
rect 17172 34298 17196 34300
rect 17252 34298 17258 34300
rect 17012 34246 17014 34298
rect 17194 34246 17196 34298
rect 16950 34244 16956 34246
rect 17012 34244 17036 34246
rect 17092 34244 17116 34246
rect 17172 34244 17196 34246
rect 17252 34244 17258 34246
rect 16950 34235 17258 34244
rect 16950 33212 17258 33221
rect 16950 33210 16956 33212
rect 17012 33210 17036 33212
rect 17092 33210 17116 33212
rect 17172 33210 17196 33212
rect 17252 33210 17258 33212
rect 17012 33158 17014 33210
rect 17194 33158 17196 33210
rect 16950 33156 16956 33158
rect 17012 33156 17036 33158
rect 17092 33156 17116 33158
rect 17172 33156 17196 33158
rect 17252 33156 17258 33158
rect 16950 33147 17258 33156
rect 16950 32124 17258 32133
rect 16950 32122 16956 32124
rect 17012 32122 17036 32124
rect 17092 32122 17116 32124
rect 17172 32122 17196 32124
rect 17252 32122 17258 32124
rect 17012 32070 17014 32122
rect 17194 32070 17196 32122
rect 16950 32068 16956 32070
rect 17012 32068 17036 32070
rect 17092 32068 17116 32070
rect 17172 32068 17196 32070
rect 17252 32068 17258 32070
rect 16950 32059 17258 32068
rect 16580 31136 16632 31142
rect 16580 31078 16632 31084
rect 16950 31036 17258 31045
rect 16950 31034 16956 31036
rect 17012 31034 17036 31036
rect 17092 31034 17116 31036
rect 17172 31034 17196 31036
rect 17252 31034 17258 31036
rect 17012 30982 17014 31034
rect 17194 30982 17196 31034
rect 16950 30980 16956 30982
rect 17012 30980 17036 30982
rect 17092 30980 17116 30982
rect 17172 30980 17196 30982
rect 17252 30980 17258 30982
rect 16950 30971 17258 30980
rect 16856 30048 16908 30054
rect 16856 29990 16908 29996
rect 16868 29170 16896 29990
rect 16950 29948 17258 29957
rect 16950 29946 16956 29948
rect 17012 29946 17036 29948
rect 17092 29946 17116 29948
rect 17172 29946 17196 29948
rect 17252 29946 17258 29948
rect 17012 29894 17014 29946
rect 17194 29894 17196 29946
rect 16950 29892 16956 29894
rect 17012 29892 17036 29894
rect 17092 29892 17116 29894
rect 17172 29892 17196 29894
rect 17252 29892 17258 29894
rect 16950 29883 17258 29892
rect 16856 29164 16908 29170
rect 16856 29106 16908 29112
rect 16950 28860 17258 28869
rect 16950 28858 16956 28860
rect 17012 28858 17036 28860
rect 17092 28858 17116 28860
rect 17172 28858 17196 28860
rect 17252 28858 17258 28860
rect 17012 28806 17014 28858
rect 17194 28806 17196 28858
rect 16950 28804 16956 28806
rect 17012 28804 17036 28806
rect 17092 28804 17116 28806
rect 17172 28804 17196 28806
rect 17252 28804 17258 28806
rect 16950 28795 17258 28804
rect 16950 27772 17258 27781
rect 16950 27770 16956 27772
rect 17012 27770 17036 27772
rect 17092 27770 17116 27772
rect 17172 27770 17196 27772
rect 17252 27770 17258 27772
rect 17012 27718 17014 27770
rect 17194 27718 17196 27770
rect 16950 27716 16956 27718
rect 17012 27716 17036 27718
rect 17092 27716 17116 27718
rect 17172 27716 17196 27718
rect 17252 27716 17258 27718
rect 16950 27707 17258 27716
rect 15844 27396 15896 27402
rect 15844 27338 15896 27344
rect 15856 25362 15884 27338
rect 16950 26684 17258 26693
rect 16950 26682 16956 26684
rect 17012 26682 17036 26684
rect 17092 26682 17116 26684
rect 17172 26682 17196 26684
rect 17252 26682 17258 26684
rect 17012 26630 17014 26682
rect 17194 26630 17196 26682
rect 16950 26628 16956 26630
rect 17012 26628 17036 26630
rect 17092 26628 17116 26630
rect 17172 26628 17196 26630
rect 17252 26628 17258 26630
rect 16950 26619 17258 26628
rect 16950 25596 17258 25605
rect 16950 25594 16956 25596
rect 17012 25594 17036 25596
rect 17092 25594 17116 25596
rect 17172 25594 17196 25596
rect 17252 25594 17258 25596
rect 17012 25542 17014 25594
rect 17194 25542 17196 25594
rect 16950 25540 16956 25542
rect 17012 25540 17036 25542
rect 17092 25540 17116 25542
rect 17172 25540 17196 25542
rect 17252 25540 17258 25542
rect 16950 25531 17258 25540
rect 15844 25356 15896 25362
rect 15844 25298 15896 25304
rect 16950 24508 17258 24517
rect 16950 24506 16956 24508
rect 17012 24506 17036 24508
rect 17092 24506 17116 24508
rect 17172 24506 17196 24508
rect 17252 24506 17258 24508
rect 17012 24454 17014 24506
rect 17194 24454 17196 24506
rect 16950 24452 16956 24454
rect 17012 24452 17036 24454
rect 17092 24452 17116 24454
rect 17172 24452 17196 24454
rect 17252 24452 17258 24454
rect 16950 24443 17258 24452
rect 16950 23420 17258 23429
rect 16950 23418 16956 23420
rect 17012 23418 17036 23420
rect 17092 23418 17116 23420
rect 17172 23418 17196 23420
rect 17252 23418 17258 23420
rect 17012 23366 17014 23418
rect 17194 23366 17196 23418
rect 16950 23364 16956 23366
rect 17012 23364 17036 23366
rect 17092 23364 17116 23366
rect 17172 23364 17196 23366
rect 17252 23364 17258 23366
rect 16950 23355 17258 23364
rect 16488 23112 16540 23118
rect 16488 23054 16540 23060
rect 15660 17060 15712 17066
rect 15660 17002 15712 17008
rect 15476 16584 15528 16590
rect 15476 16526 15528 16532
rect 16500 13326 16528 23054
rect 16950 22332 17258 22341
rect 16950 22330 16956 22332
rect 17012 22330 17036 22332
rect 17092 22330 17116 22332
rect 17172 22330 17196 22332
rect 17252 22330 17258 22332
rect 17012 22278 17014 22330
rect 17194 22278 17196 22330
rect 16950 22276 16956 22278
rect 17012 22276 17036 22278
rect 17092 22276 17116 22278
rect 17172 22276 17196 22278
rect 17252 22276 17258 22278
rect 16950 22267 17258 22276
rect 16950 21244 17258 21253
rect 16950 21242 16956 21244
rect 17012 21242 17036 21244
rect 17092 21242 17116 21244
rect 17172 21242 17196 21244
rect 17252 21242 17258 21244
rect 17012 21190 17014 21242
rect 17194 21190 17196 21242
rect 16950 21188 16956 21190
rect 17012 21188 17036 21190
rect 17092 21188 17116 21190
rect 17172 21188 17196 21190
rect 17252 21188 17258 21190
rect 16950 21179 17258 21188
rect 16950 20156 17258 20165
rect 16950 20154 16956 20156
rect 17012 20154 17036 20156
rect 17092 20154 17116 20156
rect 17172 20154 17196 20156
rect 17252 20154 17258 20156
rect 17012 20102 17014 20154
rect 17194 20102 17196 20154
rect 16950 20100 16956 20102
rect 17012 20100 17036 20102
rect 17092 20100 17116 20102
rect 17172 20100 17196 20102
rect 17252 20100 17258 20102
rect 16950 20091 17258 20100
rect 16950 19068 17258 19077
rect 16950 19066 16956 19068
rect 17012 19066 17036 19068
rect 17092 19066 17116 19068
rect 17172 19066 17196 19068
rect 17252 19066 17258 19068
rect 17012 19014 17014 19066
rect 17194 19014 17196 19066
rect 16950 19012 16956 19014
rect 17012 19012 17036 19014
rect 17092 19012 17116 19014
rect 17172 19012 17196 19014
rect 17252 19012 17258 19014
rect 16950 19003 17258 19012
rect 17328 18698 17356 44134
rect 17420 34678 17448 53994
rect 17512 51950 17540 64466
rect 17610 64220 17918 64229
rect 17610 64218 17616 64220
rect 17672 64218 17696 64220
rect 17752 64218 17776 64220
rect 17832 64218 17856 64220
rect 17912 64218 17918 64220
rect 17672 64166 17674 64218
rect 17854 64166 17856 64218
rect 17610 64164 17616 64166
rect 17672 64164 17696 64166
rect 17752 64164 17776 64166
rect 17832 64164 17856 64166
rect 17912 64164 17918 64166
rect 17610 64155 17918 64164
rect 18708 63986 18736 68342
rect 19892 64320 19944 64326
rect 19892 64262 19944 64268
rect 18972 64048 19024 64054
rect 18972 63990 19024 63996
rect 18604 63980 18656 63986
rect 18604 63922 18656 63928
rect 18696 63980 18748 63986
rect 18696 63922 18748 63928
rect 18512 63776 18564 63782
rect 18512 63718 18564 63724
rect 17610 63132 17918 63141
rect 17610 63130 17616 63132
rect 17672 63130 17696 63132
rect 17752 63130 17776 63132
rect 17832 63130 17856 63132
rect 17912 63130 17918 63132
rect 17672 63078 17674 63130
rect 17854 63078 17856 63130
rect 17610 63076 17616 63078
rect 17672 63076 17696 63078
rect 17752 63076 17776 63078
rect 17832 63076 17856 63078
rect 17912 63076 17918 63078
rect 17610 63067 17918 63076
rect 17610 62044 17918 62053
rect 17610 62042 17616 62044
rect 17672 62042 17696 62044
rect 17752 62042 17776 62044
rect 17832 62042 17856 62044
rect 17912 62042 17918 62044
rect 17672 61990 17674 62042
rect 17854 61990 17856 62042
rect 17610 61988 17616 61990
rect 17672 61988 17696 61990
rect 17752 61988 17776 61990
rect 17832 61988 17856 61990
rect 17912 61988 17918 61990
rect 17610 61979 17918 61988
rect 17610 60956 17918 60965
rect 17610 60954 17616 60956
rect 17672 60954 17696 60956
rect 17752 60954 17776 60956
rect 17832 60954 17856 60956
rect 17912 60954 17918 60956
rect 17672 60902 17674 60954
rect 17854 60902 17856 60954
rect 17610 60900 17616 60902
rect 17672 60900 17696 60902
rect 17752 60900 17776 60902
rect 17832 60900 17856 60902
rect 17912 60900 17918 60902
rect 17610 60891 17918 60900
rect 17610 59868 17918 59877
rect 17610 59866 17616 59868
rect 17672 59866 17696 59868
rect 17752 59866 17776 59868
rect 17832 59866 17856 59868
rect 17912 59866 17918 59868
rect 17672 59814 17674 59866
rect 17854 59814 17856 59866
rect 17610 59812 17616 59814
rect 17672 59812 17696 59814
rect 17752 59812 17776 59814
rect 17832 59812 17856 59814
rect 17912 59812 17918 59814
rect 17610 59803 17918 59812
rect 17610 58780 17918 58789
rect 17610 58778 17616 58780
rect 17672 58778 17696 58780
rect 17752 58778 17776 58780
rect 17832 58778 17856 58780
rect 17912 58778 17918 58780
rect 17672 58726 17674 58778
rect 17854 58726 17856 58778
rect 17610 58724 17616 58726
rect 17672 58724 17696 58726
rect 17752 58724 17776 58726
rect 17832 58724 17856 58726
rect 17912 58724 17918 58726
rect 17610 58715 17918 58724
rect 17610 57692 17918 57701
rect 17610 57690 17616 57692
rect 17672 57690 17696 57692
rect 17752 57690 17776 57692
rect 17832 57690 17856 57692
rect 17912 57690 17918 57692
rect 17672 57638 17674 57690
rect 17854 57638 17856 57690
rect 17610 57636 17616 57638
rect 17672 57636 17696 57638
rect 17752 57636 17776 57638
rect 17832 57636 17856 57638
rect 17912 57636 17918 57638
rect 17610 57627 17918 57636
rect 17610 56604 17918 56613
rect 17610 56602 17616 56604
rect 17672 56602 17696 56604
rect 17752 56602 17776 56604
rect 17832 56602 17856 56604
rect 17912 56602 17918 56604
rect 17672 56550 17674 56602
rect 17854 56550 17856 56602
rect 17610 56548 17616 56550
rect 17672 56548 17696 56550
rect 17752 56548 17776 56550
rect 17832 56548 17856 56550
rect 17912 56548 17918 56550
rect 17610 56539 17918 56548
rect 17610 55516 17918 55525
rect 17610 55514 17616 55516
rect 17672 55514 17696 55516
rect 17752 55514 17776 55516
rect 17832 55514 17856 55516
rect 17912 55514 17918 55516
rect 17672 55462 17674 55514
rect 17854 55462 17856 55514
rect 17610 55460 17616 55462
rect 17672 55460 17696 55462
rect 17752 55460 17776 55462
rect 17832 55460 17856 55462
rect 17912 55460 17918 55462
rect 17610 55451 17918 55460
rect 17610 54428 17918 54437
rect 17610 54426 17616 54428
rect 17672 54426 17696 54428
rect 17752 54426 17776 54428
rect 17832 54426 17856 54428
rect 17912 54426 17918 54428
rect 17672 54374 17674 54426
rect 17854 54374 17856 54426
rect 17610 54372 17616 54374
rect 17672 54372 17696 54374
rect 17752 54372 17776 54374
rect 17832 54372 17856 54374
rect 17912 54372 17918 54374
rect 17610 54363 17918 54372
rect 17610 53340 17918 53349
rect 17610 53338 17616 53340
rect 17672 53338 17696 53340
rect 17752 53338 17776 53340
rect 17832 53338 17856 53340
rect 17912 53338 17918 53340
rect 17672 53286 17674 53338
rect 17854 53286 17856 53338
rect 17610 53284 17616 53286
rect 17672 53284 17696 53286
rect 17752 53284 17776 53286
rect 17832 53284 17856 53286
rect 17912 53284 17918 53286
rect 17610 53275 17918 53284
rect 17610 52252 17918 52261
rect 17610 52250 17616 52252
rect 17672 52250 17696 52252
rect 17752 52250 17776 52252
rect 17832 52250 17856 52252
rect 17912 52250 17918 52252
rect 17672 52198 17674 52250
rect 17854 52198 17856 52250
rect 17610 52196 17616 52198
rect 17672 52196 17696 52198
rect 17752 52196 17776 52198
rect 17832 52196 17856 52198
rect 17912 52196 17918 52198
rect 17610 52187 17918 52196
rect 17500 51944 17552 51950
rect 17500 51886 17552 51892
rect 17512 51406 17540 51886
rect 17500 51400 17552 51406
rect 17500 51342 17552 51348
rect 17960 51400 18012 51406
rect 17960 51342 18012 51348
rect 17610 51164 17918 51173
rect 17610 51162 17616 51164
rect 17672 51162 17696 51164
rect 17752 51162 17776 51164
rect 17832 51162 17856 51164
rect 17912 51162 17918 51164
rect 17672 51110 17674 51162
rect 17854 51110 17856 51162
rect 17610 51108 17616 51110
rect 17672 51108 17696 51110
rect 17752 51108 17776 51110
rect 17832 51108 17856 51110
rect 17912 51108 17918 51110
rect 17610 51099 17918 51108
rect 17610 50076 17918 50085
rect 17610 50074 17616 50076
rect 17672 50074 17696 50076
rect 17752 50074 17776 50076
rect 17832 50074 17856 50076
rect 17912 50074 17918 50076
rect 17672 50022 17674 50074
rect 17854 50022 17856 50074
rect 17610 50020 17616 50022
rect 17672 50020 17696 50022
rect 17752 50020 17776 50022
rect 17832 50020 17856 50022
rect 17912 50020 17918 50022
rect 17610 50011 17918 50020
rect 17610 48988 17918 48997
rect 17610 48986 17616 48988
rect 17672 48986 17696 48988
rect 17752 48986 17776 48988
rect 17832 48986 17856 48988
rect 17912 48986 17918 48988
rect 17672 48934 17674 48986
rect 17854 48934 17856 48986
rect 17610 48932 17616 48934
rect 17672 48932 17696 48934
rect 17752 48932 17776 48934
rect 17832 48932 17856 48934
rect 17912 48932 17918 48934
rect 17610 48923 17918 48932
rect 17610 47900 17918 47909
rect 17610 47898 17616 47900
rect 17672 47898 17696 47900
rect 17752 47898 17776 47900
rect 17832 47898 17856 47900
rect 17912 47898 17918 47900
rect 17672 47846 17674 47898
rect 17854 47846 17856 47898
rect 17610 47844 17616 47846
rect 17672 47844 17696 47846
rect 17752 47844 17776 47846
rect 17832 47844 17856 47846
rect 17912 47844 17918 47846
rect 17610 47835 17918 47844
rect 17610 46812 17918 46821
rect 17610 46810 17616 46812
rect 17672 46810 17696 46812
rect 17752 46810 17776 46812
rect 17832 46810 17856 46812
rect 17912 46810 17918 46812
rect 17672 46758 17674 46810
rect 17854 46758 17856 46810
rect 17610 46756 17616 46758
rect 17672 46756 17696 46758
rect 17752 46756 17776 46758
rect 17832 46756 17856 46758
rect 17912 46756 17918 46758
rect 17610 46747 17918 46756
rect 17610 45724 17918 45733
rect 17610 45722 17616 45724
rect 17672 45722 17696 45724
rect 17752 45722 17776 45724
rect 17832 45722 17856 45724
rect 17912 45722 17918 45724
rect 17672 45670 17674 45722
rect 17854 45670 17856 45722
rect 17610 45668 17616 45670
rect 17672 45668 17696 45670
rect 17752 45668 17776 45670
rect 17832 45668 17856 45670
rect 17912 45668 17918 45670
rect 17610 45659 17918 45668
rect 17610 44636 17918 44645
rect 17610 44634 17616 44636
rect 17672 44634 17696 44636
rect 17752 44634 17776 44636
rect 17832 44634 17856 44636
rect 17912 44634 17918 44636
rect 17672 44582 17674 44634
rect 17854 44582 17856 44634
rect 17610 44580 17616 44582
rect 17672 44580 17696 44582
rect 17752 44580 17776 44582
rect 17832 44580 17856 44582
rect 17912 44580 17918 44582
rect 17610 44571 17918 44580
rect 17610 43548 17918 43557
rect 17610 43546 17616 43548
rect 17672 43546 17696 43548
rect 17752 43546 17776 43548
rect 17832 43546 17856 43548
rect 17912 43546 17918 43548
rect 17672 43494 17674 43546
rect 17854 43494 17856 43546
rect 17610 43492 17616 43494
rect 17672 43492 17696 43494
rect 17752 43492 17776 43494
rect 17832 43492 17856 43494
rect 17912 43492 17918 43494
rect 17610 43483 17918 43492
rect 17610 42460 17918 42469
rect 17610 42458 17616 42460
rect 17672 42458 17696 42460
rect 17752 42458 17776 42460
rect 17832 42458 17856 42460
rect 17912 42458 17918 42460
rect 17672 42406 17674 42458
rect 17854 42406 17856 42458
rect 17610 42404 17616 42406
rect 17672 42404 17696 42406
rect 17752 42404 17776 42406
rect 17832 42404 17856 42406
rect 17912 42404 17918 42406
rect 17610 42395 17918 42404
rect 17610 41372 17918 41381
rect 17610 41370 17616 41372
rect 17672 41370 17696 41372
rect 17752 41370 17776 41372
rect 17832 41370 17856 41372
rect 17912 41370 17918 41372
rect 17672 41318 17674 41370
rect 17854 41318 17856 41370
rect 17610 41316 17616 41318
rect 17672 41316 17696 41318
rect 17752 41316 17776 41318
rect 17832 41316 17856 41318
rect 17912 41316 17918 41318
rect 17610 41307 17918 41316
rect 17500 40520 17552 40526
rect 17500 40462 17552 40468
rect 17408 34672 17460 34678
rect 17408 34614 17460 34620
rect 17512 31906 17540 40462
rect 17610 40284 17918 40293
rect 17610 40282 17616 40284
rect 17672 40282 17696 40284
rect 17752 40282 17776 40284
rect 17832 40282 17856 40284
rect 17912 40282 17918 40284
rect 17672 40230 17674 40282
rect 17854 40230 17856 40282
rect 17610 40228 17616 40230
rect 17672 40228 17696 40230
rect 17752 40228 17776 40230
rect 17832 40228 17856 40230
rect 17912 40228 17918 40230
rect 17610 40219 17918 40228
rect 17610 39196 17918 39205
rect 17610 39194 17616 39196
rect 17672 39194 17696 39196
rect 17752 39194 17776 39196
rect 17832 39194 17856 39196
rect 17912 39194 17918 39196
rect 17672 39142 17674 39194
rect 17854 39142 17856 39194
rect 17610 39140 17616 39142
rect 17672 39140 17696 39142
rect 17752 39140 17776 39142
rect 17832 39140 17856 39142
rect 17912 39140 17918 39142
rect 17610 39131 17918 39140
rect 17610 38108 17918 38117
rect 17610 38106 17616 38108
rect 17672 38106 17696 38108
rect 17752 38106 17776 38108
rect 17832 38106 17856 38108
rect 17912 38106 17918 38108
rect 17672 38054 17674 38106
rect 17854 38054 17856 38106
rect 17610 38052 17616 38054
rect 17672 38052 17696 38054
rect 17752 38052 17776 38054
rect 17832 38052 17856 38054
rect 17912 38052 17918 38054
rect 17610 38043 17918 38052
rect 17610 37020 17918 37029
rect 17610 37018 17616 37020
rect 17672 37018 17696 37020
rect 17752 37018 17776 37020
rect 17832 37018 17856 37020
rect 17912 37018 17918 37020
rect 17672 36966 17674 37018
rect 17854 36966 17856 37018
rect 17610 36964 17616 36966
rect 17672 36964 17696 36966
rect 17752 36964 17776 36966
rect 17832 36964 17856 36966
rect 17912 36964 17918 36966
rect 17610 36955 17918 36964
rect 17610 35932 17918 35941
rect 17610 35930 17616 35932
rect 17672 35930 17696 35932
rect 17752 35930 17776 35932
rect 17832 35930 17856 35932
rect 17912 35930 17918 35932
rect 17672 35878 17674 35930
rect 17854 35878 17856 35930
rect 17610 35876 17616 35878
rect 17672 35876 17696 35878
rect 17752 35876 17776 35878
rect 17832 35876 17856 35878
rect 17912 35876 17918 35878
rect 17610 35867 17918 35876
rect 17610 34844 17918 34853
rect 17610 34842 17616 34844
rect 17672 34842 17696 34844
rect 17752 34842 17776 34844
rect 17832 34842 17856 34844
rect 17912 34842 17918 34844
rect 17672 34790 17674 34842
rect 17854 34790 17856 34842
rect 17610 34788 17616 34790
rect 17672 34788 17696 34790
rect 17752 34788 17776 34790
rect 17832 34788 17856 34790
rect 17912 34788 17918 34790
rect 17610 34779 17918 34788
rect 17610 33756 17918 33765
rect 17610 33754 17616 33756
rect 17672 33754 17696 33756
rect 17752 33754 17776 33756
rect 17832 33754 17856 33756
rect 17912 33754 17918 33756
rect 17672 33702 17674 33754
rect 17854 33702 17856 33754
rect 17610 33700 17616 33702
rect 17672 33700 17696 33702
rect 17752 33700 17776 33702
rect 17832 33700 17856 33702
rect 17912 33700 17918 33702
rect 17610 33691 17918 33700
rect 17610 32668 17918 32677
rect 17610 32666 17616 32668
rect 17672 32666 17696 32668
rect 17752 32666 17776 32668
rect 17832 32666 17856 32668
rect 17912 32666 17918 32668
rect 17672 32614 17674 32666
rect 17854 32614 17856 32666
rect 17610 32612 17616 32614
rect 17672 32612 17696 32614
rect 17752 32612 17776 32614
rect 17832 32612 17856 32614
rect 17912 32612 17918 32614
rect 17610 32603 17918 32612
rect 17420 31878 17540 31906
rect 17420 31754 17448 31878
rect 17420 31726 17540 31754
rect 17408 31476 17460 31482
rect 17408 31418 17460 31424
rect 17420 29850 17448 31418
rect 17408 29844 17460 29850
rect 17408 29786 17460 29792
rect 17512 28150 17540 31726
rect 17610 31580 17918 31589
rect 17610 31578 17616 31580
rect 17672 31578 17696 31580
rect 17752 31578 17776 31580
rect 17832 31578 17856 31580
rect 17912 31578 17918 31580
rect 17672 31526 17674 31578
rect 17854 31526 17856 31578
rect 17610 31524 17616 31526
rect 17672 31524 17696 31526
rect 17752 31524 17776 31526
rect 17832 31524 17856 31526
rect 17912 31524 17918 31526
rect 17610 31515 17918 31524
rect 17610 30492 17918 30501
rect 17610 30490 17616 30492
rect 17672 30490 17696 30492
rect 17752 30490 17776 30492
rect 17832 30490 17856 30492
rect 17912 30490 17918 30492
rect 17672 30438 17674 30490
rect 17854 30438 17856 30490
rect 17610 30436 17616 30438
rect 17672 30436 17696 30438
rect 17752 30436 17776 30438
rect 17832 30436 17856 30438
rect 17912 30436 17918 30438
rect 17610 30427 17918 30436
rect 17610 29404 17918 29413
rect 17610 29402 17616 29404
rect 17672 29402 17696 29404
rect 17752 29402 17776 29404
rect 17832 29402 17856 29404
rect 17912 29402 17918 29404
rect 17672 29350 17674 29402
rect 17854 29350 17856 29402
rect 17610 29348 17616 29350
rect 17672 29348 17696 29350
rect 17752 29348 17776 29350
rect 17832 29348 17856 29350
rect 17912 29348 17918 29350
rect 17610 29339 17918 29348
rect 17972 29238 18000 51342
rect 18052 32360 18104 32366
rect 18052 32302 18104 32308
rect 17960 29232 18012 29238
rect 17960 29174 18012 29180
rect 17960 28688 18012 28694
rect 17960 28630 18012 28636
rect 17972 28422 18000 28630
rect 17960 28416 18012 28422
rect 17960 28358 18012 28364
rect 17610 28316 17918 28325
rect 17610 28314 17616 28316
rect 17672 28314 17696 28316
rect 17752 28314 17776 28316
rect 17832 28314 17856 28316
rect 17912 28314 17918 28316
rect 17672 28262 17674 28314
rect 17854 28262 17856 28314
rect 17610 28260 17616 28262
rect 17672 28260 17696 28262
rect 17752 28260 17776 28262
rect 17832 28260 17856 28262
rect 17912 28260 17918 28262
rect 17610 28251 17918 28260
rect 17500 28144 17552 28150
rect 17500 28086 17552 28092
rect 17610 27228 17918 27237
rect 17610 27226 17616 27228
rect 17672 27226 17696 27228
rect 17752 27226 17776 27228
rect 17832 27226 17856 27228
rect 17912 27226 17918 27228
rect 17672 27174 17674 27226
rect 17854 27174 17856 27226
rect 17610 27172 17616 27174
rect 17672 27172 17696 27174
rect 17752 27172 17776 27174
rect 17832 27172 17856 27174
rect 17912 27172 17918 27174
rect 17610 27163 17918 27172
rect 18064 27062 18092 32302
rect 18144 31272 18196 31278
rect 18144 31214 18196 31220
rect 18156 29102 18184 31214
rect 18420 30048 18472 30054
rect 18420 29990 18472 29996
rect 18432 29850 18460 29990
rect 18420 29844 18472 29850
rect 18420 29786 18472 29792
rect 18524 29238 18552 63718
rect 18616 36038 18644 63922
rect 18708 52426 18736 63922
rect 18696 52420 18748 52426
rect 18696 52362 18748 52368
rect 18708 51474 18736 52362
rect 18696 51468 18748 51474
rect 18696 51410 18748 51416
rect 18696 45824 18748 45830
rect 18696 45766 18748 45772
rect 18604 36032 18656 36038
rect 18604 35974 18656 35980
rect 18604 33312 18656 33318
rect 18604 33254 18656 33260
rect 18616 30190 18644 33254
rect 18604 30184 18656 30190
rect 18604 30126 18656 30132
rect 18420 29232 18472 29238
rect 18420 29174 18472 29180
rect 18512 29232 18564 29238
rect 18512 29174 18564 29180
rect 18144 29096 18196 29102
rect 18144 29038 18196 29044
rect 18156 27470 18184 29038
rect 18144 27464 18196 27470
rect 18144 27406 18196 27412
rect 18052 27056 18104 27062
rect 18052 26998 18104 27004
rect 17610 26140 17918 26149
rect 17610 26138 17616 26140
rect 17672 26138 17696 26140
rect 17752 26138 17776 26140
rect 17832 26138 17856 26140
rect 17912 26138 17918 26140
rect 17672 26086 17674 26138
rect 17854 26086 17856 26138
rect 17610 26084 17616 26086
rect 17672 26084 17696 26086
rect 17752 26084 17776 26086
rect 17832 26084 17856 26086
rect 17912 26084 17918 26086
rect 17610 26075 17918 26084
rect 17610 25052 17918 25061
rect 17610 25050 17616 25052
rect 17672 25050 17696 25052
rect 17752 25050 17776 25052
rect 17832 25050 17856 25052
rect 17912 25050 17918 25052
rect 17672 24998 17674 25050
rect 17854 24998 17856 25050
rect 17610 24996 17616 24998
rect 17672 24996 17696 24998
rect 17752 24996 17776 24998
rect 17832 24996 17856 24998
rect 17912 24996 17918 24998
rect 17610 24987 17918 24996
rect 17610 23964 17918 23973
rect 17610 23962 17616 23964
rect 17672 23962 17696 23964
rect 17752 23962 17776 23964
rect 17832 23962 17856 23964
rect 17912 23962 17918 23964
rect 17672 23910 17674 23962
rect 17854 23910 17856 23962
rect 17610 23908 17616 23910
rect 17672 23908 17696 23910
rect 17752 23908 17776 23910
rect 17832 23908 17856 23910
rect 17912 23908 17918 23910
rect 17610 23899 17918 23908
rect 17610 22876 17918 22885
rect 17610 22874 17616 22876
rect 17672 22874 17696 22876
rect 17752 22874 17776 22876
rect 17832 22874 17856 22876
rect 17912 22874 17918 22876
rect 17672 22822 17674 22874
rect 17854 22822 17856 22874
rect 17610 22820 17616 22822
rect 17672 22820 17696 22822
rect 17752 22820 17776 22822
rect 17832 22820 17856 22822
rect 17912 22820 17918 22822
rect 17610 22811 17918 22820
rect 17610 21788 17918 21797
rect 17610 21786 17616 21788
rect 17672 21786 17696 21788
rect 17752 21786 17776 21788
rect 17832 21786 17856 21788
rect 17912 21786 17918 21788
rect 17672 21734 17674 21786
rect 17854 21734 17856 21786
rect 17610 21732 17616 21734
rect 17672 21732 17696 21734
rect 17752 21732 17776 21734
rect 17832 21732 17856 21734
rect 17912 21732 17918 21734
rect 17610 21723 17918 21732
rect 17610 20700 17918 20709
rect 17610 20698 17616 20700
rect 17672 20698 17696 20700
rect 17752 20698 17776 20700
rect 17832 20698 17856 20700
rect 17912 20698 17918 20700
rect 17672 20646 17674 20698
rect 17854 20646 17856 20698
rect 17610 20644 17616 20646
rect 17672 20644 17696 20646
rect 17752 20644 17776 20646
rect 17832 20644 17856 20646
rect 17912 20644 17918 20646
rect 17610 20635 17918 20644
rect 17610 19612 17918 19621
rect 17610 19610 17616 19612
rect 17672 19610 17696 19612
rect 17752 19610 17776 19612
rect 17832 19610 17856 19612
rect 17912 19610 17918 19612
rect 17672 19558 17674 19610
rect 17854 19558 17856 19610
rect 17610 19556 17616 19558
rect 17672 19556 17696 19558
rect 17752 19556 17776 19558
rect 17832 19556 17856 19558
rect 17912 19556 17918 19558
rect 17610 19547 17918 19556
rect 17316 18692 17368 18698
rect 17316 18634 17368 18640
rect 17610 18524 17918 18533
rect 17610 18522 17616 18524
rect 17672 18522 17696 18524
rect 17752 18522 17776 18524
rect 17832 18522 17856 18524
rect 17912 18522 17918 18524
rect 17672 18470 17674 18522
rect 17854 18470 17856 18522
rect 17610 18468 17616 18470
rect 17672 18468 17696 18470
rect 17752 18468 17776 18470
rect 17832 18468 17856 18470
rect 17912 18468 17918 18470
rect 17610 18459 17918 18468
rect 16950 17980 17258 17989
rect 16950 17978 16956 17980
rect 17012 17978 17036 17980
rect 17092 17978 17116 17980
rect 17172 17978 17196 17980
rect 17252 17978 17258 17980
rect 17012 17926 17014 17978
rect 17194 17926 17196 17978
rect 16950 17924 16956 17926
rect 17012 17924 17036 17926
rect 17092 17924 17116 17926
rect 17172 17924 17196 17926
rect 17252 17924 17258 17926
rect 16950 17915 17258 17924
rect 17610 17436 17918 17445
rect 17610 17434 17616 17436
rect 17672 17434 17696 17436
rect 17752 17434 17776 17436
rect 17832 17434 17856 17436
rect 17912 17434 17918 17436
rect 17672 17382 17674 17434
rect 17854 17382 17856 17434
rect 17610 17380 17616 17382
rect 17672 17380 17696 17382
rect 17752 17380 17776 17382
rect 17832 17380 17856 17382
rect 17912 17380 17918 17382
rect 17610 17371 17918 17380
rect 17316 16992 17368 16998
rect 17316 16934 17368 16940
rect 16950 16892 17258 16901
rect 16950 16890 16956 16892
rect 17012 16890 17036 16892
rect 17092 16890 17116 16892
rect 17172 16890 17196 16892
rect 17252 16890 17258 16892
rect 17012 16838 17014 16890
rect 17194 16838 17196 16890
rect 16950 16836 16956 16838
rect 17012 16836 17036 16838
rect 17092 16836 17116 16838
rect 17172 16836 17196 16838
rect 17252 16836 17258 16838
rect 16950 16827 17258 16836
rect 16950 15804 17258 15813
rect 16950 15802 16956 15804
rect 17012 15802 17036 15804
rect 17092 15802 17116 15804
rect 17172 15802 17196 15804
rect 17252 15802 17258 15804
rect 17012 15750 17014 15802
rect 17194 15750 17196 15802
rect 16950 15748 16956 15750
rect 17012 15748 17036 15750
rect 17092 15748 17116 15750
rect 17172 15748 17196 15750
rect 17252 15748 17258 15750
rect 16950 15739 17258 15748
rect 16950 14716 17258 14725
rect 16950 14714 16956 14716
rect 17012 14714 17036 14716
rect 17092 14714 17116 14716
rect 17172 14714 17196 14716
rect 17252 14714 17258 14716
rect 17012 14662 17014 14714
rect 17194 14662 17196 14714
rect 16950 14660 16956 14662
rect 17012 14660 17036 14662
rect 17092 14660 17116 14662
rect 17172 14660 17196 14662
rect 17252 14660 17258 14662
rect 16950 14651 17258 14660
rect 16950 13628 17258 13637
rect 16950 13626 16956 13628
rect 17012 13626 17036 13628
rect 17092 13626 17116 13628
rect 17172 13626 17196 13628
rect 17252 13626 17258 13628
rect 17012 13574 17014 13626
rect 17194 13574 17196 13626
rect 16950 13572 16956 13574
rect 17012 13572 17036 13574
rect 17092 13572 17116 13574
rect 17172 13572 17196 13574
rect 17252 13572 17258 13574
rect 16950 13563 17258 13572
rect 15844 13320 15896 13326
rect 15844 13262 15896 13268
rect 16488 13320 16540 13326
rect 16488 13262 16540 13268
rect 15856 4690 15884 13262
rect 16950 12540 17258 12549
rect 16950 12538 16956 12540
rect 17012 12538 17036 12540
rect 17092 12538 17116 12540
rect 17172 12538 17196 12540
rect 17252 12538 17258 12540
rect 17012 12486 17014 12538
rect 17194 12486 17196 12538
rect 16950 12484 16956 12486
rect 17012 12484 17036 12486
rect 17092 12484 17116 12486
rect 17172 12484 17196 12486
rect 17252 12484 17258 12486
rect 16950 12475 17258 12484
rect 16950 11452 17258 11461
rect 16950 11450 16956 11452
rect 17012 11450 17036 11452
rect 17092 11450 17116 11452
rect 17172 11450 17196 11452
rect 17252 11450 17258 11452
rect 17012 11398 17014 11450
rect 17194 11398 17196 11450
rect 16950 11396 16956 11398
rect 17012 11396 17036 11398
rect 17092 11396 17116 11398
rect 17172 11396 17196 11398
rect 17252 11396 17258 11398
rect 16950 11387 17258 11396
rect 16950 10364 17258 10373
rect 16950 10362 16956 10364
rect 17012 10362 17036 10364
rect 17092 10362 17116 10364
rect 17172 10362 17196 10364
rect 17252 10362 17258 10364
rect 17012 10310 17014 10362
rect 17194 10310 17196 10362
rect 16950 10308 16956 10310
rect 17012 10308 17036 10310
rect 17092 10308 17116 10310
rect 17172 10308 17196 10310
rect 17252 10308 17258 10310
rect 16950 10299 17258 10308
rect 17328 9654 17356 16934
rect 17610 16348 17918 16357
rect 17610 16346 17616 16348
rect 17672 16346 17696 16348
rect 17752 16346 17776 16348
rect 17832 16346 17856 16348
rect 17912 16346 17918 16348
rect 17672 16294 17674 16346
rect 17854 16294 17856 16346
rect 17610 16292 17616 16294
rect 17672 16292 17696 16294
rect 17752 16292 17776 16294
rect 17832 16292 17856 16294
rect 17912 16292 17918 16294
rect 17610 16283 17918 16292
rect 17610 15260 17918 15269
rect 17610 15258 17616 15260
rect 17672 15258 17696 15260
rect 17752 15258 17776 15260
rect 17832 15258 17856 15260
rect 17912 15258 17918 15260
rect 17672 15206 17674 15258
rect 17854 15206 17856 15258
rect 17610 15204 17616 15206
rect 17672 15204 17696 15206
rect 17752 15204 17776 15206
rect 17832 15204 17856 15206
rect 17912 15204 17918 15206
rect 17610 15195 17918 15204
rect 17610 14172 17918 14181
rect 17610 14170 17616 14172
rect 17672 14170 17696 14172
rect 17752 14170 17776 14172
rect 17832 14170 17856 14172
rect 17912 14170 17918 14172
rect 17672 14118 17674 14170
rect 17854 14118 17856 14170
rect 17610 14116 17616 14118
rect 17672 14116 17696 14118
rect 17752 14116 17776 14118
rect 17832 14116 17856 14118
rect 17912 14116 17918 14118
rect 17610 14107 17918 14116
rect 17610 13084 17918 13093
rect 17610 13082 17616 13084
rect 17672 13082 17696 13084
rect 17752 13082 17776 13084
rect 17832 13082 17856 13084
rect 17912 13082 17918 13084
rect 17672 13030 17674 13082
rect 17854 13030 17856 13082
rect 17610 13028 17616 13030
rect 17672 13028 17696 13030
rect 17752 13028 17776 13030
rect 17832 13028 17856 13030
rect 17912 13028 17918 13030
rect 17610 13019 17918 13028
rect 18064 12238 18092 26998
rect 18156 24818 18184 27406
rect 18144 24812 18196 24818
rect 18144 24754 18196 24760
rect 18432 17338 18460 29174
rect 18512 17604 18564 17610
rect 18512 17546 18564 17552
rect 18420 17332 18472 17338
rect 18420 17274 18472 17280
rect 18524 17270 18552 17546
rect 18604 17332 18656 17338
rect 18604 17274 18656 17280
rect 18512 17264 18564 17270
rect 18512 17206 18564 17212
rect 18616 14346 18644 17274
rect 18708 16522 18736 45766
rect 18880 38956 18932 38962
rect 18880 38898 18932 38904
rect 18892 34202 18920 38898
rect 18984 37738 19012 63990
rect 19616 62212 19668 62218
rect 19616 62154 19668 62160
rect 19628 51338 19656 62154
rect 19904 62150 19932 64262
rect 20720 63776 20772 63782
rect 20720 63718 20772 63724
rect 20352 63368 20404 63374
rect 20352 63310 20404 63316
rect 19892 62144 19944 62150
rect 19892 62086 19944 62092
rect 19616 51332 19668 51338
rect 19616 51274 19668 51280
rect 19904 46986 19932 62086
rect 19984 51332 20036 51338
rect 19984 51274 20036 51280
rect 19892 46980 19944 46986
rect 19892 46922 19944 46928
rect 19432 45008 19484 45014
rect 19432 44950 19484 44956
rect 19444 44878 19472 44950
rect 19432 44872 19484 44878
rect 19432 44814 19484 44820
rect 18972 37732 19024 37738
rect 18972 37674 19024 37680
rect 18984 36242 19012 37674
rect 18972 36236 19024 36242
rect 18972 36178 19024 36184
rect 18880 34196 18932 34202
rect 18880 34138 18932 34144
rect 18892 33318 18920 34138
rect 18880 33312 18932 33318
rect 18880 33254 18932 33260
rect 19156 32360 19208 32366
rect 19156 32302 19208 32308
rect 18880 30252 18932 30258
rect 18880 30194 18932 30200
rect 18788 30184 18840 30190
rect 18788 30126 18840 30132
rect 18800 17338 18828 30126
rect 18788 17332 18840 17338
rect 18788 17274 18840 17280
rect 18696 16516 18748 16522
rect 18696 16458 18748 16464
rect 18604 14340 18656 14346
rect 18604 14282 18656 14288
rect 18616 14006 18644 14282
rect 18604 14000 18656 14006
rect 18604 13942 18656 13948
rect 18800 12238 18828 17274
rect 18892 17270 18920 30194
rect 19168 28694 19196 32302
rect 19156 28688 19208 28694
rect 19156 28630 19208 28636
rect 19340 28416 19392 28422
rect 19340 28358 19392 28364
rect 19352 22778 19380 28358
rect 19340 22772 19392 22778
rect 19340 22714 19392 22720
rect 19444 19922 19472 44814
rect 19996 41478 20024 51274
rect 19984 41472 20036 41478
rect 19984 41414 20036 41420
rect 19614 34504 19670 34513
rect 19614 34439 19670 34448
rect 19628 33998 19656 34439
rect 19616 33992 19668 33998
rect 19616 33934 19668 33940
rect 19616 31408 19668 31414
rect 19616 31350 19668 31356
rect 19524 29028 19576 29034
rect 19524 28970 19576 28976
rect 19432 19916 19484 19922
rect 19432 19858 19484 19864
rect 18880 17264 18932 17270
rect 18880 17206 18932 17212
rect 19536 17202 19564 28970
rect 19628 23254 19656 31350
rect 19996 28626 20024 41414
rect 20364 35562 20392 63310
rect 20536 55684 20588 55690
rect 20536 55626 20588 55632
rect 20548 55282 20576 55626
rect 20536 55276 20588 55282
rect 20536 55218 20588 55224
rect 20352 35556 20404 35562
rect 20352 35498 20404 35504
rect 20732 29238 20760 63718
rect 20996 48544 21048 48550
rect 20996 48486 21048 48492
rect 20904 44940 20956 44946
rect 20904 44882 20956 44888
rect 20916 38962 20944 44882
rect 20904 38956 20956 38962
rect 20904 38898 20956 38904
rect 20916 35894 20944 38898
rect 20824 35866 20944 35894
rect 20720 29232 20772 29238
rect 20720 29174 20772 29180
rect 19984 28620 20036 28626
rect 19984 28562 20036 28568
rect 19800 28552 19852 28558
rect 19800 28494 19852 28500
rect 19812 28422 19840 28494
rect 19800 28416 19852 28422
rect 19800 28358 19852 28364
rect 20444 28416 20496 28422
rect 20444 28358 20496 28364
rect 20456 28082 20484 28358
rect 20444 28076 20496 28082
rect 20444 28018 20496 28024
rect 19984 27600 20036 27606
rect 19984 27542 20036 27548
rect 19996 27470 20024 27542
rect 20456 27538 20484 28018
rect 20444 27532 20496 27538
rect 20444 27474 20496 27480
rect 19984 27464 20036 27470
rect 19984 27406 20036 27412
rect 19996 27130 20024 27406
rect 19984 27124 20036 27130
rect 19984 27066 20036 27072
rect 19616 23248 19668 23254
rect 19616 23190 19668 23196
rect 20456 17270 20484 27474
rect 20824 17882 20852 35866
rect 20904 31816 20956 31822
rect 20904 31758 20956 31764
rect 20916 31278 20944 31758
rect 20904 31272 20956 31278
rect 20904 31214 20956 31220
rect 20812 17876 20864 17882
rect 20812 17818 20864 17824
rect 20444 17264 20496 17270
rect 20444 17206 20496 17212
rect 19524 17196 19576 17202
rect 19524 17138 19576 17144
rect 18052 12232 18104 12238
rect 18052 12174 18104 12180
rect 18604 12232 18656 12238
rect 18604 12174 18656 12180
rect 18788 12232 18840 12238
rect 18788 12174 18840 12180
rect 17610 11996 17918 12005
rect 17610 11994 17616 11996
rect 17672 11994 17696 11996
rect 17752 11994 17776 11996
rect 17832 11994 17856 11996
rect 17912 11994 17918 11996
rect 17672 11942 17674 11994
rect 17854 11942 17856 11994
rect 17610 11940 17616 11942
rect 17672 11940 17696 11942
rect 17752 11940 17776 11942
rect 17832 11940 17856 11942
rect 17912 11940 17918 11942
rect 17610 11931 17918 11940
rect 17610 10908 17918 10917
rect 17610 10906 17616 10908
rect 17672 10906 17696 10908
rect 17752 10906 17776 10908
rect 17832 10906 17856 10908
rect 17912 10906 17918 10908
rect 17672 10854 17674 10906
rect 17854 10854 17856 10906
rect 17610 10852 17616 10854
rect 17672 10852 17696 10854
rect 17752 10852 17776 10854
rect 17832 10852 17856 10854
rect 17912 10852 17918 10854
rect 17610 10843 17918 10852
rect 17610 9820 17918 9829
rect 17610 9818 17616 9820
rect 17672 9818 17696 9820
rect 17752 9818 17776 9820
rect 17832 9818 17856 9820
rect 17912 9818 17918 9820
rect 17672 9766 17674 9818
rect 17854 9766 17856 9818
rect 17610 9764 17616 9766
rect 17672 9764 17696 9766
rect 17752 9764 17776 9766
rect 17832 9764 17856 9766
rect 17912 9764 17918 9766
rect 17610 9755 17918 9764
rect 17316 9648 17368 9654
rect 17316 9590 17368 9596
rect 16950 9276 17258 9285
rect 16950 9274 16956 9276
rect 17012 9274 17036 9276
rect 17092 9274 17116 9276
rect 17172 9274 17196 9276
rect 17252 9274 17258 9276
rect 17012 9222 17014 9274
rect 17194 9222 17196 9274
rect 16950 9220 16956 9222
rect 17012 9220 17036 9222
rect 17092 9220 17116 9222
rect 17172 9220 17196 9222
rect 17252 9220 17258 9222
rect 16950 9211 17258 9220
rect 17610 8732 17918 8741
rect 17610 8730 17616 8732
rect 17672 8730 17696 8732
rect 17752 8730 17776 8732
rect 17832 8730 17856 8732
rect 17912 8730 17918 8732
rect 17672 8678 17674 8730
rect 17854 8678 17856 8730
rect 17610 8676 17616 8678
rect 17672 8676 17696 8678
rect 17752 8676 17776 8678
rect 17832 8676 17856 8678
rect 17912 8676 17918 8678
rect 17610 8667 17918 8676
rect 16950 8188 17258 8197
rect 16950 8186 16956 8188
rect 17012 8186 17036 8188
rect 17092 8186 17116 8188
rect 17172 8186 17196 8188
rect 17252 8186 17258 8188
rect 17012 8134 17014 8186
rect 17194 8134 17196 8186
rect 16950 8132 16956 8134
rect 17012 8132 17036 8134
rect 17092 8132 17116 8134
rect 17172 8132 17196 8134
rect 17252 8132 17258 8134
rect 16950 8123 17258 8132
rect 17610 7644 17918 7653
rect 17610 7642 17616 7644
rect 17672 7642 17696 7644
rect 17752 7642 17776 7644
rect 17832 7642 17856 7644
rect 17912 7642 17918 7644
rect 17672 7590 17674 7642
rect 17854 7590 17856 7642
rect 17610 7588 17616 7590
rect 17672 7588 17696 7590
rect 17752 7588 17776 7590
rect 17832 7588 17856 7590
rect 17912 7588 17918 7590
rect 17610 7579 17918 7588
rect 16950 7100 17258 7109
rect 16950 7098 16956 7100
rect 17012 7098 17036 7100
rect 17092 7098 17116 7100
rect 17172 7098 17196 7100
rect 17252 7098 17258 7100
rect 17012 7046 17014 7098
rect 17194 7046 17196 7098
rect 16950 7044 16956 7046
rect 17012 7044 17036 7046
rect 17092 7044 17116 7046
rect 17172 7044 17196 7046
rect 17252 7044 17258 7046
rect 16950 7035 17258 7044
rect 17610 6556 17918 6565
rect 17610 6554 17616 6556
rect 17672 6554 17696 6556
rect 17752 6554 17776 6556
rect 17832 6554 17856 6556
rect 17912 6554 17918 6556
rect 17672 6502 17674 6554
rect 17854 6502 17856 6554
rect 17610 6500 17616 6502
rect 17672 6500 17696 6502
rect 17752 6500 17776 6502
rect 17832 6500 17856 6502
rect 17912 6500 17918 6502
rect 17610 6491 17918 6500
rect 16950 6012 17258 6021
rect 16950 6010 16956 6012
rect 17012 6010 17036 6012
rect 17092 6010 17116 6012
rect 17172 6010 17196 6012
rect 17252 6010 17258 6012
rect 17012 5958 17014 6010
rect 17194 5958 17196 6010
rect 16950 5956 16956 5958
rect 17012 5956 17036 5958
rect 17092 5956 17116 5958
rect 17172 5956 17196 5958
rect 17252 5956 17258 5958
rect 16950 5947 17258 5956
rect 17610 5468 17918 5477
rect 17610 5466 17616 5468
rect 17672 5466 17696 5468
rect 17752 5466 17776 5468
rect 17832 5466 17856 5468
rect 17912 5466 17918 5468
rect 17672 5414 17674 5466
rect 17854 5414 17856 5466
rect 17610 5412 17616 5414
rect 17672 5412 17696 5414
rect 17752 5412 17776 5414
rect 17832 5412 17856 5414
rect 17912 5412 17918 5414
rect 17610 5403 17918 5412
rect 16950 4924 17258 4933
rect 16950 4922 16956 4924
rect 17012 4922 17036 4924
rect 17092 4922 17116 4924
rect 17172 4922 17196 4924
rect 17252 4922 17258 4924
rect 17012 4870 17014 4922
rect 17194 4870 17196 4922
rect 16950 4868 16956 4870
rect 17012 4868 17036 4870
rect 17092 4868 17116 4870
rect 17172 4868 17196 4870
rect 17252 4868 17258 4870
rect 16950 4859 17258 4868
rect 15844 4684 15896 4690
rect 15844 4626 15896 4632
rect 17610 4380 17918 4389
rect 17610 4378 17616 4380
rect 17672 4378 17696 4380
rect 17752 4378 17776 4380
rect 17832 4378 17856 4380
rect 17912 4378 17918 4380
rect 17672 4326 17674 4378
rect 17854 4326 17856 4378
rect 17610 4324 17616 4326
rect 17672 4324 17696 4326
rect 17752 4324 17776 4326
rect 17832 4324 17856 4326
rect 17912 4324 17918 4326
rect 17610 4315 17918 4324
rect 16950 3836 17258 3845
rect 16950 3834 16956 3836
rect 17012 3834 17036 3836
rect 17092 3834 17116 3836
rect 17172 3834 17196 3836
rect 17252 3834 17258 3836
rect 17012 3782 17014 3834
rect 17194 3782 17196 3834
rect 16950 3780 16956 3782
rect 17012 3780 17036 3782
rect 17092 3780 17116 3782
rect 17172 3780 17196 3782
rect 17252 3780 17258 3782
rect 16950 3771 17258 3780
rect 17610 3292 17918 3301
rect 17610 3290 17616 3292
rect 17672 3290 17696 3292
rect 17752 3290 17776 3292
rect 17832 3290 17856 3292
rect 17912 3290 17918 3292
rect 17672 3238 17674 3290
rect 17854 3238 17856 3290
rect 17610 3236 17616 3238
rect 17672 3236 17696 3238
rect 17752 3236 17776 3238
rect 17832 3236 17856 3238
rect 17912 3236 17918 3238
rect 17610 3227 17918 3236
rect 16950 2748 17258 2757
rect 16950 2746 16956 2748
rect 17012 2746 17036 2748
rect 17092 2746 17116 2748
rect 17172 2746 17196 2748
rect 17252 2746 17258 2748
rect 17012 2694 17014 2746
rect 17194 2694 17196 2746
rect 16950 2692 16956 2694
rect 17012 2692 17036 2694
rect 17092 2692 17116 2694
rect 17172 2692 17196 2694
rect 17252 2692 17258 2694
rect 16950 2683 17258 2692
rect 15200 2576 15252 2582
rect 15200 2518 15252 2524
rect 18616 2514 18644 12174
rect 19536 9654 19564 17138
rect 20916 16250 20944 31214
rect 21008 19922 21036 48486
rect 21088 33856 21140 33862
rect 21086 33824 21088 33833
rect 21140 33824 21142 33833
rect 21086 33759 21142 33768
rect 21192 30870 21220 69362
rect 21950 69116 22258 69125
rect 21950 69114 21956 69116
rect 22012 69114 22036 69116
rect 22092 69114 22116 69116
rect 22172 69114 22196 69116
rect 22252 69114 22258 69116
rect 22012 69062 22014 69114
rect 22194 69062 22196 69114
rect 21950 69060 21956 69062
rect 22012 69060 22036 69062
rect 22092 69060 22116 69062
rect 22172 69060 22196 69062
rect 22252 69060 22258 69062
rect 21950 69051 22258 69060
rect 26950 69116 27258 69125
rect 26950 69114 26956 69116
rect 27012 69114 27036 69116
rect 27092 69114 27116 69116
rect 27172 69114 27196 69116
rect 27252 69114 27258 69116
rect 27012 69062 27014 69114
rect 27194 69062 27196 69114
rect 26950 69060 26956 69062
rect 27012 69060 27036 69062
rect 27092 69060 27116 69062
rect 27172 69060 27196 69062
rect 27252 69060 27258 69062
rect 26950 69051 27258 69060
rect 22610 68572 22918 68581
rect 22610 68570 22616 68572
rect 22672 68570 22696 68572
rect 22752 68570 22776 68572
rect 22832 68570 22856 68572
rect 22912 68570 22918 68572
rect 22672 68518 22674 68570
rect 22854 68518 22856 68570
rect 22610 68516 22616 68518
rect 22672 68516 22696 68518
rect 22752 68516 22776 68518
rect 22832 68516 22856 68518
rect 22912 68516 22918 68518
rect 22610 68507 22918 68516
rect 21950 68028 22258 68037
rect 21950 68026 21956 68028
rect 22012 68026 22036 68028
rect 22092 68026 22116 68028
rect 22172 68026 22196 68028
rect 22252 68026 22258 68028
rect 22012 67974 22014 68026
rect 22194 67974 22196 68026
rect 21950 67972 21956 67974
rect 22012 67972 22036 67974
rect 22092 67972 22116 67974
rect 22172 67972 22196 67974
rect 22252 67972 22258 67974
rect 21950 67963 22258 67972
rect 26950 68028 27258 68037
rect 26950 68026 26956 68028
rect 27012 68026 27036 68028
rect 27092 68026 27116 68028
rect 27172 68026 27196 68028
rect 27252 68026 27258 68028
rect 27012 67974 27014 68026
rect 27194 67974 27196 68026
rect 26950 67972 26956 67974
rect 27012 67972 27036 67974
rect 27092 67972 27116 67974
rect 27172 67972 27196 67974
rect 27252 67972 27258 67974
rect 26950 67963 27258 67972
rect 24860 67652 24912 67658
rect 24860 67594 24912 67600
rect 25044 67652 25096 67658
rect 25044 67594 25096 67600
rect 22610 67484 22918 67493
rect 22610 67482 22616 67484
rect 22672 67482 22696 67484
rect 22752 67482 22776 67484
rect 22832 67482 22856 67484
rect 22912 67482 22918 67484
rect 22672 67430 22674 67482
rect 22854 67430 22856 67482
rect 22610 67428 22616 67430
rect 22672 67428 22696 67430
rect 22752 67428 22776 67430
rect 22832 67428 22856 67430
rect 22912 67428 22918 67430
rect 22610 67419 22918 67428
rect 21950 66940 22258 66949
rect 21950 66938 21956 66940
rect 22012 66938 22036 66940
rect 22092 66938 22116 66940
rect 22172 66938 22196 66940
rect 22252 66938 22258 66940
rect 22012 66886 22014 66938
rect 22194 66886 22196 66938
rect 21950 66884 21956 66886
rect 22012 66884 22036 66886
rect 22092 66884 22116 66886
rect 22172 66884 22196 66886
rect 22252 66884 22258 66886
rect 21950 66875 22258 66884
rect 22610 66396 22918 66405
rect 22610 66394 22616 66396
rect 22672 66394 22696 66396
rect 22752 66394 22776 66396
rect 22832 66394 22856 66396
rect 22912 66394 22918 66396
rect 22672 66342 22674 66394
rect 22854 66342 22856 66394
rect 22610 66340 22616 66342
rect 22672 66340 22696 66342
rect 22752 66340 22776 66342
rect 22832 66340 22856 66342
rect 22912 66340 22918 66342
rect 22610 66331 22918 66340
rect 24216 66156 24268 66162
rect 24216 66098 24268 66104
rect 21950 65852 22258 65861
rect 21950 65850 21956 65852
rect 22012 65850 22036 65852
rect 22092 65850 22116 65852
rect 22172 65850 22196 65852
rect 22252 65850 22258 65852
rect 22012 65798 22014 65850
rect 22194 65798 22196 65850
rect 21950 65796 21956 65798
rect 22012 65796 22036 65798
rect 22092 65796 22116 65798
rect 22172 65796 22196 65798
rect 22252 65796 22258 65798
rect 21950 65787 22258 65796
rect 22610 65308 22918 65317
rect 22610 65306 22616 65308
rect 22672 65306 22696 65308
rect 22752 65306 22776 65308
rect 22832 65306 22856 65308
rect 22912 65306 22918 65308
rect 22672 65254 22674 65306
rect 22854 65254 22856 65306
rect 22610 65252 22616 65254
rect 22672 65252 22696 65254
rect 22752 65252 22776 65254
rect 22832 65252 22856 65254
rect 22912 65252 22918 65254
rect 22610 65243 22918 65252
rect 23112 65136 23164 65142
rect 23112 65078 23164 65084
rect 23020 65068 23072 65074
rect 23020 65010 23072 65016
rect 22376 64932 22428 64938
rect 22376 64874 22428 64880
rect 21950 64764 22258 64773
rect 21950 64762 21956 64764
rect 22012 64762 22036 64764
rect 22092 64762 22116 64764
rect 22172 64762 22196 64764
rect 22252 64762 22258 64764
rect 22012 64710 22014 64762
rect 22194 64710 22196 64762
rect 21950 64708 21956 64710
rect 22012 64708 22036 64710
rect 22092 64708 22116 64710
rect 22172 64708 22196 64710
rect 22252 64708 22258 64710
rect 21950 64699 22258 64708
rect 21824 63980 21876 63986
rect 21824 63922 21876 63928
rect 21836 55826 21864 63922
rect 21950 63676 22258 63685
rect 21950 63674 21956 63676
rect 22012 63674 22036 63676
rect 22092 63674 22116 63676
rect 22172 63674 22196 63676
rect 22252 63674 22258 63676
rect 22012 63622 22014 63674
rect 22194 63622 22196 63674
rect 21950 63620 21956 63622
rect 22012 63620 22036 63622
rect 22092 63620 22116 63622
rect 22172 63620 22196 63622
rect 22252 63620 22258 63622
rect 21950 63611 22258 63620
rect 21950 62588 22258 62597
rect 21950 62586 21956 62588
rect 22012 62586 22036 62588
rect 22092 62586 22116 62588
rect 22172 62586 22196 62588
rect 22252 62586 22258 62588
rect 22012 62534 22014 62586
rect 22194 62534 22196 62586
rect 21950 62532 21956 62534
rect 22012 62532 22036 62534
rect 22092 62532 22116 62534
rect 22172 62532 22196 62534
rect 22252 62532 22258 62534
rect 21950 62523 22258 62532
rect 21950 61500 22258 61509
rect 21950 61498 21956 61500
rect 22012 61498 22036 61500
rect 22092 61498 22116 61500
rect 22172 61498 22196 61500
rect 22252 61498 22258 61500
rect 22012 61446 22014 61498
rect 22194 61446 22196 61498
rect 21950 61444 21956 61446
rect 22012 61444 22036 61446
rect 22092 61444 22116 61446
rect 22172 61444 22196 61446
rect 22252 61444 22258 61446
rect 21950 61435 22258 61444
rect 21950 60412 22258 60421
rect 21950 60410 21956 60412
rect 22012 60410 22036 60412
rect 22092 60410 22116 60412
rect 22172 60410 22196 60412
rect 22252 60410 22258 60412
rect 22012 60358 22014 60410
rect 22194 60358 22196 60410
rect 21950 60356 21956 60358
rect 22012 60356 22036 60358
rect 22092 60356 22116 60358
rect 22172 60356 22196 60358
rect 22252 60356 22258 60358
rect 21950 60347 22258 60356
rect 21950 59324 22258 59333
rect 21950 59322 21956 59324
rect 22012 59322 22036 59324
rect 22092 59322 22116 59324
rect 22172 59322 22196 59324
rect 22252 59322 22258 59324
rect 22012 59270 22014 59322
rect 22194 59270 22196 59322
rect 21950 59268 21956 59270
rect 22012 59268 22036 59270
rect 22092 59268 22116 59270
rect 22172 59268 22196 59270
rect 22252 59268 22258 59270
rect 21950 59259 22258 59268
rect 21950 58236 22258 58245
rect 21950 58234 21956 58236
rect 22012 58234 22036 58236
rect 22092 58234 22116 58236
rect 22172 58234 22196 58236
rect 22252 58234 22258 58236
rect 22012 58182 22014 58234
rect 22194 58182 22196 58234
rect 21950 58180 21956 58182
rect 22012 58180 22036 58182
rect 22092 58180 22116 58182
rect 22172 58180 22196 58182
rect 22252 58180 22258 58182
rect 21950 58171 22258 58180
rect 21950 57148 22258 57157
rect 21950 57146 21956 57148
rect 22012 57146 22036 57148
rect 22092 57146 22116 57148
rect 22172 57146 22196 57148
rect 22252 57146 22258 57148
rect 22012 57094 22014 57146
rect 22194 57094 22196 57146
rect 21950 57092 21956 57094
rect 22012 57092 22036 57094
rect 22092 57092 22116 57094
rect 22172 57092 22196 57094
rect 22252 57092 22258 57094
rect 21950 57083 22258 57092
rect 21950 56060 22258 56069
rect 21950 56058 21956 56060
rect 22012 56058 22036 56060
rect 22092 56058 22116 56060
rect 22172 56058 22196 56060
rect 22252 56058 22258 56060
rect 22012 56006 22014 56058
rect 22194 56006 22196 56058
rect 21950 56004 21956 56006
rect 22012 56004 22036 56006
rect 22092 56004 22116 56006
rect 22172 56004 22196 56006
rect 22252 56004 22258 56006
rect 21950 55995 22258 56004
rect 21456 55820 21508 55826
rect 21456 55762 21508 55768
rect 21824 55820 21876 55826
rect 21824 55762 21876 55768
rect 21364 51876 21416 51882
rect 21364 51818 21416 51824
rect 21376 38962 21404 51818
rect 21468 47598 21496 55762
rect 22284 55344 22336 55350
rect 22284 55286 22336 55292
rect 21950 54972 22258 54981
rect 21950 54970 21956 54972
rect 22012 54970 22036 54972
rect 22092 54970 22116 54972
rect 22172 54970 22196 54972
rect 22252 54970 22258 54972
rect 22012 54918 22014 54970
rect 22194 54918 22196 54970
rect 21950 54916 21956 54918
rect 22012 54916 22036 54918
rect 22092 54916 22116 54918
rect 22172 54916 22196 54918
rect 22252 54916 22258 54918
rect 21950 54907 22258 54916
rect 21950 53884 22258 53893
rect 21950 53882 21956 53884
rect 22012 53882 22036 53884
rect 22092 53882 22116 53884
rect 22172 53882 22196 53884
rect 22252 53882 22258 53884
rect 22012 53830 22014 53882
rect 22194 53830 22196 53882
rect 21950 53828 21956 53830
rect 22012 53828 22036 53830
rect 22092 53828 22116 53830
rect 22172 53828 22196 53830
rect 22252 53828 22258 53830
rect 21950 53819 22258 53828
rect 21950 52796 22258 52805
rect 21950 52794 21956 52796
rect 22012 52794 22036 52796
rect 22092 52794 22116 52796
rect 22172 52794 22196 52796
rect 22252 52794 22258 52796
rect 22012 52742 22014 52794
rect 22194 52742 22196 52794
rect 21950 52740 21956 52742
rect 22012 52740 22036 52742
rect 22092 52740 22116 52742
rect 22172 52740 22196 52742
rect 22252 52740 22258 52742
rect 21950 52731 22258 52740
rect 21950 51708 22258 51717
rect 21950 51706 21956 51708
rect 22012 51706 22036 51708
rect 22092 51706 22116 51708
rect 22172 51706 22196 51708
rect 22252 51706 22258 51708
rect 22012 51654 22014 51706
rect 22194 51654 22196 51706
rect 21950 51652 21956 51654
rect 22012 51652 22036 51654
rect 22092 51652 22116 51654
rect 22172 51652 22196 51654
rect 22252 51652 22258 51654
rect 21950 51643 22258 51652
rect 21950 50620 22258 50629
rect 21950 50618 21956 50620
rect 22012 50618 22036 50620
rect 22092 50618 22116 50620
rect 22172 50618 22196 50620
rect 22252 50618 22258 50620
rect 22012 50566 22014 50618
rect 22194 50566 22196 50618
rect 21950 50564 21956 50566
rect 22012 50564 22036 50566
rect 22092 50564 22116 50566
rect 22172 50564 22196 50566
rect 22252 50564 22258 50566
rect 21950 50555 22258 50564
rect 21950 49532 22258 49541
rect 21950 49530 21956 49532
rect 22012 49530 22036 49532
rect 22092 49530 22116 49532
rect 22172 49530 22196 49532
rect 22252 49530 22258 49532
rect 22012 49478 22014 49530
rect 22194 49478 22196 49530
rect 21950 49476 21956 49478
rect 22012 49476 22036 49478
rect 22092 49476 22116 49478
rect 22172 49476 22196 49478
rect 22252 49476 22258 49478
rect 21950 49467 22258 49476
rect 21640 48748 21692 48754
rect 21640 48690 21692 48696
rect 21456 47592 21508 47598
rect 21456 47534 21508 47540
rect 21364 38956 21416 38962
rect 21364 38898 21416 38904
rect 21376 31822 21404 38898
rect 21364 31816 21416 31822
rect 21364 31758 21416 31764
rect 21180 30864 21232 30870
rect 21180 30806 21232 30812
rect 20996 19916 21048 19922
rect 20996 19858 21048 19864
rect 21180 17876 21232 17882
rect 21180 17818 21232 17824
rect 21192 16658 21220 17818
rect 21180 16652 21232 16658
rect 21180 16594 21232 16600
rect 20904 16244 20956 16250
rect 20904 16186 20956 16192
rect 19524 9648 19576 9654
rect 19524 9590 19576 9596
rect 19984 9648 20036 9654
rect 19984 9590 20036 9596
rect 18880 7880 18932 7886
rect 18878 7848 18880 7857
rect 18932 7848 18934 7857
rect 18878 7783 18934 7792
rect 19996 5234 20024 9590
rect 19984 5228 20036 5234
rect 19984 5170 20036 5176
rect 21652 2854 21680 48690
rect 21950 48444 22258 48453
rect 21950 48442 21956 48444
rect 22012 48442 22036 48444
rect 22092 48442 22116 48444
rect 22172 48442 22196 48444
rect 22252 48442 22258 48444
rect 22012 48390 22014 48442
rect 22194 48390 22196 48442
rect 21950 48388 21956 48390
rect 22012 48388 22036 48390
rect 22092 48388 22116 48390
rect 22172 48388 22196 48390
rect 22252 48388 22258 48390
rect 21950 48379 22258 48388
rect 21950 47356 22258 47365
rect 21950 47354 21956 47356
rect 22012 47354 22036 47356
rect 22092 47354 22116 47356
rect 22172 47354 22196 47356
rect 22252 47354 22258 47356
rect 22012 47302 22014 47354
rect 22194 47302 22196 47354
rect 21950 47300 21956 47302
rect 22012 47300 22036 47302
rect 22092 47300 22116 47302
rect 22172 47300 22196 47302
rect 22252 47300 22258 47302
rect 21950 47291 22258 47300
rect 21950 46268 22258 46277
rect 21950 46266 21956 46268
rect 22012 46266 22036 46268
rect 22092 46266 22116 46268
rect 22172 46266 22196 46268
rect 22252 46266 22258 46268
rect 22012 46214 22014 46266
rect 22194 46214 22196 46266
rect 21950 46212 21956 46214
rect 22012 46212 22036 46214
rect 22092 46212 22116 46214
rect 22172 46212 22196 46214
rect 22252 46212 22258 46214
rect 21950 46203 22258 46212
rect 21950 45180 22258 45189
rect 21950 45178 21956 45180
rect 22012 45178 22036 45180
rect 22092 45178 22116 45180
rect 22172 45178 22196 45180
rect 22252 45178 22258 45180
rect 22012 45126 22014 45178
rect 22194 45126 22196 45178
rect 21950 45124 21956 45126
rect 22012 45124 22036 45126
rect 22092 45124 22116 45126
rect 22172 45124 22196 45126
rect 22252 45124 22258 45126
rect 21950 45115 22258 45124
rect 22296 44810 22324 55286
rect 22388 54534 22416 64874
rect 22610 64220 22918 64229
rect 22610 64218 22616 64220
rect 22672 64218 22696 64220
rect 22752 64218 22776 64220
rect 22832 64218 22856 64220
rect 22912 64218 22918 64220
rect 22672 64166 22674 64218
rect 22854 64166 22856 64218
rect 22610 64164 22616 64166
rect 22672 64164 22696 64166
rect 22752 64164 22776 64166
rect 22832 64164 22856 64166
rect 22912 64164 22918 64166
rect 22610 64155 22918 64164
rect 22610 63132 22918 63141
rect 22610 63130 22616 63132
rect 22672 63130 22696 63132
rect 22752 63130 22776 63132
rect 22832 63130 22856 63132
rect 22912 63130 22918 63132
rect 22672 63078 22674 63130
rect 22854 63078 22856 63130
rect 22610 63076 22616 63078
rect 22672 63076 22696 63078
rect 22752 63076 22776 63078
rect 22832 63076 22856 63078
rect 22912 63076 22918 63078
rect 22610 63067 22918 63076
rect 22610 62044 22918 62053
rect 22610 62042 22616 62044
rect 22672 62042 22696 62044
rect 22752 62042 22776 62044
rect 22832 62042 22856 62044
rect 22912 62042 22918 62044
rect 22672 61990 22674 62042
rect 22854 61990 22856 62042
rect 22610 61988 22616 61990
rect 22672 61988 22696 61990
rect 22752 61988 22776 61990
rect 22832 61988 22856 61990
rect 22912 61988 22918 61990
rect 22610 61979 22918 61988
rect 22610 60956 22918 60965
rect 22610 60954 22616 60956
rect 22672 60954 22696 60956
rect 22752 60954 22776 60956
rect 22832 60954 22856 60956
rect 22912 60954 22918 60956
rect 22672 60902 22674 60954
rect 22854 60902 22856 60954
rect 22610 60900 22616 60902
rect 22672 60900 22696 60902
rect 22752 60900 22776 60902
rect 22832 60900 22856 60902
rect 22912 60900 22918 60902
rect 22610 60891 22918 60900
rect 23032 60042 23060 65010
rect 23020 60036 23072 60042
rect 23020 59978 23072 59984
rect 22610 59868 22918 59877
rect 22610 59866 22616 59868
rect 22672 59866 22696 59868
rect 22752 59866 22776 59868
rect 22832 59866 22856 59868
rect 22912 59866 22918 59868
rect 22672 59814 22674 59866
rect 22854 59814 22856 59866
rect 22610 59812 22616 59814
rect 22672 59812 22696 59814
rect 22752 59812 22776 59814
rect 22832 59812 22856 59814
rect 22912 59812 22918 59814
rect 22610 59803 22918 59812
rect 22610 58780 22918 58789
rect 22610 58778 22616 58780
rect 22672 58778 22696 58780
rect 22752 58778 22776 58780
rect 22832 58778 22856 58780
rect 22912 58778 22918 58780
rect 22672 58726 22674 58778
rect 22854 58726 22856 58778
rect 22610 58724 22616 58726
rect 22672 58724 22696 58726
rect 22752 58724 22776 58726
rect 22832 58724 22856 58726
rect 22912 58724 22918 58726
rect 22610 58715 22918 58724
rect 22610 57692 22918 57701
rect 22610 57690 22616 57692
rect 22672 57690 22696 57692
rect 22752 57690 22776 57692
rect 22832 57690 22856 57692
rect 22912 57690 22918 57692
rect 22672 57638 22674 57690
rect 22854 57638 22856 57690
rect 22610 57636 22616 57638
rect 22672 57636 22696 57638
rect 22752 57636 22776 57638
rect 22832 57636 22856 57638
rect 22912 57636 22918 57638
rect 22610 57627 22918 57636
rect 23124 57458 23152 65078
rect 23296 65000 23348 65006
rect 23296 64942 23348 64948
rect 23204 59968 23256 59974
rect 23204 59910 23256 59916
rect 23112 57452 23164 57458
rect 23112 57394 23164 57400
rect 22610 56604 22918 56613
rect 22610 56602 22616 56604
rect 22672 56602 22696 56604
rect 22752 56602 22776 56604
rect 22832 56602 22856 56604
rect 22912 56602 22918 56604
rect 22672 56550 22674 56602
rect 22854 56550 22856 56602
rect 22610 56548 22616 56550
rect 22672 56548 22696 56550
rect 22752 56548 22776 56550
rect 22832 56548 22856 56550
rect 22912 56548 22918 56550
rect 22610 56539 22918 56548
rect 22610 55516 22918 55525
rect 22610 55514 22616 55516
rect 22672 55514 22696 55516
rect 22752 55514 22776 55516
rect 22832 55514 22856 55516
rect 22912 55514 22918 55516
rect 22672 55462 22674 55514
rect 22854 55462 22856 55514
rect 22610 55460 22616 55462
rect 22672 55460 22696 55462
rect 22752 55460 22776 55462
rect 22832 55460 22856 55462
rect 22912 55460 22918 55462
rect 22610 55451 22918 55460
rect 23020 55072 23072 55078
rect 23020 55014 23072 55020
rect 22376 54528 22428 54534
rect 22376 54470 22428 54476
rect 22388 54194 22416 54470
rect 22610 54428 22918 54437
rect 22610 54426 22616 54428
rect 22672 54426 22696 54428
rect 22752 54426 22776 54428
rect 22832 54426 22856 54428
rect 22912 54426 22918 54428
rect 22672 54374 22674 54426
rect 22854 54374 22856 54426
rect 22610 54372 22616 54374
rect 22672 54372 22696 54374
rect 22752 54372 22776 54374
rect 22832 54372 22856 54374
rect 22912 54372 22918 54374
rect 22610 54363 22918 54372
rect 22376 54188 22428 54194
rect 22376 54130 22428 54136
rect 22610 53340 22918 53349
rect 22610 53338 22616 53340
rect 22672 53338 22696 53340
rect 22752 53338 22776 53340
rect 22832 53338 22856 53340
rect 22912 53338 22918 53340
rect 22672 53286 22674 53338
rect 22854 53286 22856 53338
rect 22610 53284 22616 53286
rect 22672 53284 22696 53286
rect 22752 53284 22776 53286
rect 22832 53284 22856 53286
rect 22912 53284 22918 53286
rect 22610 53275 22918 53284
rect 22376 53236 22428 53242
rect 22376 53178 22428 53184
rect 22388 50726 22416 53178
rect 22610 52252 22918 52261
rect 22610 52250 22616 52252
rect 22672 52250 22696 52252
rect 22752 52250 22776 52252
rect 22832 52250 22856 52252
rect 22912 52250 22918 52252
rect 22672 52198 22674 52250
rect 22854 52198 22856 52250
rect 22610 52196 22616 52198
rect 22672 52196 22696 52198
rect 22752 52196 22776 52198
rect 22832 52196 22856 52198
rect 22912 52196 22918 52198
rect 22610 52187 22918 52196
rect 22610 51164 22918 51173
rect 22610 51162 22616 51164
rect 22672 51162 22696 51164
rect 22752 51162 22776 51164
rect 22832 51162 22856 51164
rect 22912 51162 22918 51164
rect 22672 51110 22674 51162
rect 22854 51110 22856 51162
rect 22610 51108 22616 51110
rect 22672 51108 22696 51110
rect 22752 51108 22776 51110
rect 22832 51108 22856 51110
rect 22912 51108 22918 51110
rect 22610 51099 22918 51108
rect 22376 50720 22428 50726
rect 22376 50662 22428 50668
rect 22610 50076 22918 50085
rect 22610 50074 22616 50076
rect 22672 50074 22696 50076
rect 22752 50074 22776 50076
rect 22832 50074 22856 50076
rect 22912 50074 22918 50076
rect 22672 50022 22674 50074
rect 22854 50022 22856 50074
rect 22610 50020 22616 50022
rect 22672 50020 22696 50022
rect 22752 50020 22776 50022
rect 22832 50020 22856 50022
rect 22912 50020 22918 50022
rect 22610 50011 22918 50020
rect 22610 48988 22918 48997
rect 22610 48986 22616 48988
rect 22672 48986 22696 48988
rect 22752 48986 22776 48988
rect 22832 48986 22856 48988
rect 22912 48986 22918 48988
rect 22672 48934 22674 48986
rect 22854 48934 22856 48986
rect 22610 48932 22616 48934
rect 22672 48932 22696 48934
rect 22752 48932 22776 48934
rect 22832 48932 22856 48934
rect 22912 48932 22918 48934
rect 22610 48923 22918 48932
rect 22610 47900 22918 47909
rect 22610 47898 22616 47900
rect 22672 47898 22696 47900
rect 22752 47898 22776 47900
rect 22832 47898 22856 47900
rect 22912 47898 22918 47900
rect 22672 47846 22674 47898
rect 22854 47846 22856 47898
rect 22610 47844 22616 47846
rect 22672 47844 22696 47846
rect 22752 47844 22776 47846
rect 22832 47844 22856 47846
rect 22912 47844 22918 47846
rect 22610 47835 22918 47844
rect 22610 46812 22918 46821
rect 22610 46810 22616 46812
rect 22672 46810 22696 46812
rect 22752 46810 22776 46812
rect 22832 46810 22856 46812
rect 22912 46810 22918 46812
rect 22672 46758 22674 46810
rect 22854 46758 22856 46810
rect 22610 46756 22616 46758
rect 22672 46756 22696 46758
rect 22752 46756 22776 46758
rect 22832 46756 22856 46758
rect 22912 46756 22918 46758
rect 22610 46747 22918 46756
rect 23032 45898 23060 55014
rect 23124 54262 23152 57394
rect 23112 54256 23164 54262
rect 23112 54198 23164 54204
rect 23020 45892 23072 45898
rect 23020 45834 23072 45840
rect 22610 45724 22918 45733
rect 22610 45722 22616 45724
rect 22672 45722 22696 45724
rect 22752 45722 22776 45724
rect 22832 45722 22856 45724
rect 22912 45722 22918 45724
rect 22672 45670 22674 45722
rect 22854 45670 22856 45722
rect 22610 45668 22616 45670
rect 22672 45668 22696 45670
rect 22752 45668 22776 45670
rect 22832 45668 22856 45670
rect 22912 45668 22918 45670
rect 22610 45659 22918 45668
rect 22284 44804 22336 44810
rect 22284 44746 22336 44752
rect 22468 44804 22520 44810
rect 22468 44746 22520 44752
rect 22376 44736 22428 44742
rect 22376 44678 22428 44684
rect 21950 44092 22258 44101
rect 21950 44090 21956 44092
rect 22012 44090 22036 44092
rect 22092 44090 22116 44092
rect 22172 44090 22196 44092
rect 22252 44090 22258 44092
rect 22012 44038 22014 44090
rect 22194 44038 22196 44090
rect 21950 44036 21956 44038
rect 22012 44036 22036 44038
rect 22092 44036 22116 44038
rect 22172 44036 22196 44038
rect 22252 44036 22258 44038
rect 21950 44027 22258 44036
rect 21950 43004 22258 43013
rect 21950 43002 21956 43004
rect 22012 43002 22036 43004
rect 22092 43002 22116 43004
rect 22172 43002 22196 43004
rect 22252 43002 22258 43004
rect 22012 42950 22014 43002
rect 22194 42950 22196 43002
rect 21950 42948 21956 42950
rect 22012 42948 22036 42950
rect 22092 42948 22116 42950
rect 22172 42948 22196 42950
rect 22252 42948 22258 42950
rect 21950 42939 22258 42948
rect 21950 41916 22258 41925
rect 21950 41914 21956 41916
rect 22012 41914 22036 41916
rect 22092 41914 22116 41916
rect 22172 41914 22196 41916
rect 22252 41914 22258 41916
rect 22012 41862 22014 41914
rect 22194 41862 22196 41914
rect 21950 41860 21956 41862
rect 22012 41860 22036 41862
rect 22092 41860 22116 41862
rect 22172 41860 22196 41862
rect 22252 41860 22258 41862
rect 21950 41851 22258 41860
rect 22388 41206 22416 44678
rect 22376 41200 22428 41206
rect 22376 41142 22428 41148
rect 21950 40828 22258 40837
rect 21950 40826 21956 40828
rect 22012 40826 22036 40828
rect 22092 40826 22116 40828
rect 22172 40826 22196 40828
rect 22252 40826 22258 40828
rect 22012 40774 22014 40826
rect 22194 40774 22196 40826
rect 21950 40772 21956 40774
rect 22012 40772 22036 40774
rect 22092 40772 22116 40774
rect 22172 40772 22196 40774
rect 22252 40772 22258 40774
rect 21950 40763 22258 40772
rect 21950 39740 22258 39749
rect 21950 39738 21956 39740
rect 22012 39738 22036 39740
rect 22092 39738 22116 39740
rect 22172 39738 22196 39740
rect 22252 39738 22258 39740
rect 22012 39686 22014 39738
rect 22194 39686 22196 39738
rect 21950 39684 21956 39686
rect 22012 39684 22036 39686
rect 22092 39684 22116 39686
rect 22172 39684 22196 39686
rect 22252 39684 22258 39686
rect 21950 39675 22258 39684
rect 22008 39500 22060 39506
rect 22008 39442 22060 39448
rect 22020 39030 22048 39442
rect 22192 39364 22244 39370
rect 22192 39306 22244 39312
rect 22204 39098 22232 39306
rect 22192 39092 22244 39098
rect 22192 39034 22244 39040
rect 22008 39024 22060 39030
rect 22008 38966 22060 38972
rect 21732 38752 21784 38758
rect 21732 38694 21784 38700
rect 21744 23730 21772 38694
rect 21950 38652 22258 38661
rect 21950 38650 21956 38652
rect 22012 38650 22036 38652
rect 22092 38650 22116 38652
rect 22172 38650 22196 38652
rect 22252 38650 22258 38652
rect 22012 38598 22014 38650
rect 22194 38598 22196 38650
rect 21950 38596 21956 38598
rect 22012 38596 22036 38598
rect 22092 38596 22116 38598
rect 22172 38596 22196 38598
rect 22252 38596 22258 38598
rect 21950 38587 22258 38596
rect 21950 37564 22258 37573
rect 21950 37562 21956 37564
rect 22012 37562 22036 37564
rect 22092 37562 22116 37564
rect 22172 37562 22196 37564
rect 22252 37562 22258 37564
rect 22012 37510 22014 37562
rect 22194 37510 22196 37562
rect 21950 37508 21956 37510
rect 22012 37508 22036 37510
rect 22092 37508 22116 37510
rect 22172 37508 22196 37510
rect 22252 37508 22258 37510
rect 21950 37499 22258 37508
rect 21950 36476 22258 36485
rect 21950 36474 21956 36476
rect 22012 36474 22036 36476
rect 22092 36474 22116 36476
rect 22172 36474 22196 36476
rect 22252 36474 22258 36476
rect 22012 36422 22014 36474
rect 22194 36422 22196 36474
rect 21950 36420 21956 36422
rect 22012 36420 22036 36422
rect 22092 36420 22116 36422
rect 22172 36420 22196 36422
rect 22252 36420 22258 36422
rect 21950 36411 22258 36420
rect 21950 35388 22258 35397
rect 21950 35386 21956 35388
rect 22012 35386 22036 35388
rect 22092 35386 22116 35388
rect 22172 35386 22196 35388
rect 22252 35386 22258 35388
rect 22012 35334 22014 35386
rect 22194 35334 22196 35386
rect 21950 35332 21956 35334
rect 22012 35332 22036 35334
rect 22092 35332 22116 35334
rect 22172 35332 22196 35334
rect 22252 35332 22258 35334
rect 21950 35323 22258 35332
rect 21950 34300 22258 34309
rect 21950 34298 21956 34300
rect 22012 34298 22036 34300
rect 22092 34298 22116 34300
rect 22172 34298 22196 34300
rect 22252 34298 22258 34300
rect 22012 34246 22014 34298
rect 22194 34246 22196 34298
rect 21950 34244 21956 34246
rect 22012 34244 22036 34246
rect 22092 34244 22116 34246
rect 22172 34244 22196 34246
rect 22252 34244 22258 34246
rect 21950 34235 22258 34244
rect 21950 33212 22258 33221
rect 21950 33210 21956 33212
rect 22012 33210 22036 33212
rect 22092 33210 22116 33212
rect 22172 33210 22196 33212
rect 22252 33210 22258 33212
rect 22012 33158 22014 33210
rect 22194 33158 22196 33210
rect 21950 33156 21956 33158
rect 22012 33156 22036 33158
rect 22092 33156 22116 33158
rect 22172 33156 22196 33158
rect 22252 33156 22258 33158
rect 21950 33147 22258 33156
rect 21950 32124 22258 32133
rect 21950 32122 21956 32124
rect 22012 32122 22036 32124
rect 22092 32122 22116 32124
rect 22172 32122 22196 32124
rect 22252 32122 22258 32124
rect 22012 32070 22014 32122
rect 22194 32070 22196 32122
rect 21950 32068 21956 32070
rect 22012 32068 22036 32070
rect 22092 32068 22116 32070
rect 22172 32068 22196 32070
rect 22252 32068 22258 32070
rect 21950 32059 22258 32068
rect 21950 31036 22258 31045
rect 21950 31034 21956 31036
rect 22012 31034 22036 31036
rect 22092 31034 22116 31036
rect 22172 31034 22196 31036
rect 22252 31034 22258 31036
rect 22012 30982 22014 31034
rect 22194 30982 22196 31034
rect 21950 30980 21956 30982
rect 22012 30980 22036 30982
rect 22092 30980 22116 30982
rect 22172 30980 22196 30982
rect 22252 30980 22258 30982
rect 21950 30971 22258 30980
rect 22480 30326 22508 44746
rect 22610 44636 22918 44645
rect 22610 44634 22616 44636
rect 22672 44634 22696 44636
rect 22752 44634 22776 44636
rect 22832 44634 22856 44636
rect 22912 44634 22918 44636
rect 22672 44582 22674 44634
rect 22854 44582 22856 44634
rect 22610 44580 22616 44582
rect 22672 44580 22696 44582
rect 22752 44580 22776 44582
rect 22832 44580 22856 44582
rect 22912 44580 22918 44582
rect 22610 44571 22918 44580
rect 22610 43548 22918 43557
rect 22610 43546 22616 43548
rect 22672 43546 22696 43548
rect 22752 43546 22776 43548
rect 22832 43546 22856 43548
rect 22912 43546 22918 43548
rect 22672 43494 22674 43546
rect 22854 43494 22856 43546
rect 22610 43492 22616 43494
rect 22672 43492 22696 43494
rect 22752 43492 22776 43494
rect 22832 43492 22856 43494
rect 22912 43492 22918 43494
rect 22610 43483 22918 43492
rect 22610 42460 22918 42469
rect 22610 42458 22616 42460
rect 22672 42458 22696 42460
rect 22752 42458 22776 42460
rect 22832 42458 22856 42460
rect 22912 42458 22918 42460
rect 22672 42406 22674 42458
rect 22854 42406 22856 42458
rect 22610 42404 22616 42406
rect 22672 42404 22696 42406
rect 22752 42404 22776 42406
rect 22832 42404 22856 42406
rect 22912 42404 22918 42406
rect 22610 42395 22918 42404
rect 22610 41372 22918 41381
rect 22610 41370 22616 41372
rect 22672 41370 22696 41372
rect 22752 41370 22776 41372
rect 22832 41370 22856 41372
rect 22912 41370 22918 41372
rect 22672 41318 22674 41370
rect 22854 41318 22856 41370
rect 22610 41316 22616 41318
rect 22672 41316 22696 41318
rect 22752 41316 22776 41318
rect 22832 41316 22856 41318
rect 22912 41316 22918 41318
rect 22610 41307 22918 41316
rect 22610 40284 22918 40293
rect 22610 40282 22616 40284
rect 22672 40282 22696 40284
rect 22752 40282 22776 40284
rect 22832 40282 22856 40284
rect 22912 40282 22918 40284
rect 22672 40230 22674 40282
rect 22854 40230 22856 40282
rect 22610 40228 22616 40230
rect 22672 40228 22696 40230
rect 22752 40228 22776 40230
rect 22832 40228 22856 40230
rect 22912 40228 22918 40230
rect 22610 40219 22918 40228
rect 22610 39196 22918 39205
rect 22610 39194 22616 39196
rect 22672 39194 22696 39196
rect 22752 39194 22776 39196
rect 22832 39194 22856 39196
rect 22912 39194 22918 39196
rect 22672 39142 22674 39194
rect 22854 39142 22856 39194
rect 22610 39140 22616 39142
rect 22672 39140 22696 39142
rect 22752 39140 22776 39142
rect 22832 39140 22856 39142
rect 22912 39140 22918 39142
rect 22610 39131 22918 39140
rect 23216 38962 23244 59910
rect 23308 53038 23336 64942
rect 24228 63238 24256 66098
rect 24872 64326 24900 67594
rect 24860 64320 24912 64326
rect 24860 64262 24912 64268
rect 24872 63578 24900 64262
rect 24860 63572 24912 63578
rect 24860 63514 24912 63520
rect 24216 63232 24268 63238
rect 24216 63174 24268 63180
rect 23388 60036 23440 60042
rect 23388 59978 23440 59984
rect 23400 54738 23428 59978
rect 24124 57384 24176 57390
rect 24124 57326 24176 57332
rect 23388 54732 23440 54738
rect 23388 54674 23440 54680
rect 23400 54126 23428 54674
rect 23388 54120 23440 54126
rect 23388 54062 23440 54068
rect 23296 53032 23348 53038
rect 23296 52974 23348 52980
rect 23204 38956 23256 38962
rect 23204 38898 23256 38904
rect 22610 38108 22918 38117
rect 22610 38106 22616 38108
rect 22672 38106 22696 38108
rect 22752 38106 22776 38108
rect 22832 38106 22856 38108
rect 22912 38106 22918 38108
rect 22672 38054 22674 38106
rect 22854 38054 22856 38106
rect 22610 38052 22616 38054
rect 22672 38052 22696 38054
rect 22752 38052 22776 38054
rect 22832 38052 22856 38054
rect 22912 38052 22918 38054
rect 22610 38043 22918 38052
rect 22610 37020 22918 37029
rect 22610 37018 22616 37020
rect 22672 37018 22696 37020
rect 22752 37018 22776 37020
rect 22832 37018 22856 37020
rect 22912 37018 22918 37020
rect 22672 36966 22674 37018
rect 22854 36966 22856 37018
rect 22610 36964 22616 36966
rect 22672 36964 22696 36966
rect 22752 36964 22776 36966
rect 22832 36964 22856 36966
rect 22912 36964 22918 36966
rect 22610 36955 22918 36964
rect 22610 35932 22918 35941
rect 22610 35930 22616 35932
rect 22672 35930 22696 35932
rect 22752 35930 22776 35932
rect 22832 35930 22856 35932
rect 22912 35930 22918 35932
rect 22672 35878 22674 35930
rect 22854 35878 22856 35930
rect 22610 35876 22616 35878
rect 22672 35876 22696 35878
rect 22752 35876 22776 35878
rect 22832 35876 22856 35878
rect 22912 35876 22918 35878
rect 22610 35867 22918 35876
rect 22610 34844 22918 34853
rect 22610 34842 22616 34844
rect 22672 34842 22696 34844
rect 22752 34842 22776 34844
rect 22832 34842 22856 34844
rect 22912 34842 22918 34844
rect 22672 34790 22674 34842
rect 22854 34790 22856 34842
rect 22610 34788 22616 34790
rect 22672 34788 22696 34790
rect 22752 34788 22776 34790
rect 22832 34788 22856 34790
rect 22912 34788 22918 34790
rect 22610 34779 22918 34788
rect 23308 34066 23336 52974
rect 24136 52494 24164 57326
rect 24124 52488 24176 52494
rect 24124 52430 24176 52436
rect 23756 39432 23808 39438
rect 23756 39374 23808 39380
rect 23296 34060 23348 34066
rect 23296 34002 23348 34008
rect 22610 33756 22918 33765
rect 22610 33754 22616 33756
rect 22672 33754 22696 33756
rect 22752 33754 22776 33756
rect 22832 33754 22856 33756
rect 22912 33754 22918 33756
rect 22672 33702 22674 33754
rect 22854 33702 22856 33754
rect 22610 33700 22616 33702
rect 22672 33700 22696 33702
rect 22752 33700 22776 33702
rect 22832 33700 22856 33702
rect 22912 33700 22918 33702
rect 22610 33691 22918 33700
rect 22610 32668 22918 32677
rect 22610 32666 22616 32668
rect 22672 32666 22696 32668
rect 22752 32666 22776 32668
rect 22832 32666 22856 32668
rect 22912 32666 22918 32668
rect 22672 32614 22674 32666
rect 22854 32614 22856 32666
rect 22610 32612 22616 32614
rect 22672 32612 22696 32614
rect 22752 32612 22776 32614
rect 22832 32612 22856 32614
rect 22912 32612 22918 32614
rect 22610 32603 22918 32612
rect 23308 31754 23336 34002
rect 23308 31726 23428 31754
rect 22610 31580 22918 31589
rect 22610 31578 22616 31580
rect 22672 31578 22696 31580
rect 22752 31578 22776 31580
rect 22832 31578 22856 31580
rect 22912 31578 22918 31580
rect 22672 31526 22674 31578
rect 22854 31526 22856 31578
rect 22610 31524 22616 31526
rect 22672 31524 22696 31526
rect 22752 31524 22776 31526
rect 22832 31524 22856 31526
rect 22912 31524 22918 31526
rect 22610 31515 22918 31524
rect 22610 30492 22918 30501
rect 22610 30490 22616 30492
rect 22672 30490 22696 30492
rect 22752 30490 22776 30492
rect 22832 30490 22856 30492
rect 22912 30490 22918 30492
rect 22672 30438 22674 30490
rect 22854 30438 22856 30490
rect 22610 30436 22616 30438
rect 22672 30436 22696 30438
rect 22752 30436 22776 30438
rect 22832 30436 22856 30438
rect 22912 30436 22918 30438
rect 22610 30427 22918 30436
rect 22468 30320 22520 30326
rect 22468 30262 22520 30268
rect 23020 30320 23072 30326
rect 23020 30262 23072 30268
rect 21950 29948 22258 29957
rect 21950 29946 21956 29948
rect 22012 29946 22036 29948
rect 22092 29946 22116 29948
rect 22172 29946 22196 29948
rect 22252 29946 22258 29948
rect 22012 29894 22014 29946
rect 22194 29894 22196 29946
rect 21950 29892 21956 29894
rect 22012 29892 22036 29894
rect 22092 29892 22116 29894
rect 22172 29892 22196 29894
rect 22252 29892 22258 29894
rect 21950 29883 22258 29892
rect 22610 29404 22918 29413
rect 22610 29402 22616 29404
rect 22672 29402 22696 29404
rect 22752 29402 22776 29404
rect 22832 29402 22856 29404
rect 22912 29402 22918 29404
rect 22672 29350 22674 29402
rect 22854 29350 22856 29402
rect 22610 29348 22616 29350
rect 22672 29348 22696 29350
rect 22752 29348 22776 29350
rect 22832 29348 22856 29350
rect 22912 29348 22918 29350
rect 22610 29339 22918 29348
rect 23032 29170 23060 30262
rect 23020 29164 23072 29170
rect 23020 29106 23072 29112
rect 21950 28860 22258 28869
rect 21950 28858 21956 28860
rect 22012 28858 22036 28860
rect 22092 28858 22116 28860
rect 22172 28858 22196 28860
rect 22252 28858 22258 28860
rect 22012 28806 22014 28858
rect 22194 28806 22196 28858
rect 21950 28804 21956 28806
rect 22012 28804 22036 28806
rect 22092 28804 22116 28806
rect 22172 28804 22196 28806
rect 22252 28804 22258 28806
rect 21950 28795 22258 28804
rect 22008 28484 22060 28490
rect 22008 28426 22060 28432
rect 22020 28082 22048 28426
rect 22610 28316 22918 28325
rect 22610 28314 22616 28316
rect 22672 28314 22696 28316
rect 22752 28314 22776 28316
rect 22832 28314 22856 28316
rect 22912 28314 22918 28316
rect 22672 28262 22674 28314
rect 22854 28262 22856 28314
rect 22610 28260 22616 28262
rect 22672 28260 22696 28262
rect 22752 28260 22776 28262
rect 22832 28260 22856 28262
rect 22912 28260 22918 28262
rect 22610 28251 22918 28260
rect 22008 28076 22060 28082
rect 22008 28018 22060 28024
rect 21950 27772 22258 27781
rect 21950 27770 21956 27772
rect 22012 27770 22036 27772
rect 22092 27770 22116 27772
rect 22172 27770 22196 27772
rect 22252 27770 22258 27772
rect 22012 27718 22014 27770
rect 22194 27718 22196 27770
rect 21950 27716 21956 27718
rect 22012 27716 22036 27718
rect 22092 27716 22116 27718
rect 22172 27716 22196 27718
rect 22252 27716 22258 27718
rect 21950 27707 22258 27716
rect 22468 27668 22520 27674
rect 22468 27610 22520 27616
rect 21950 26684 22258 26693
rect 21950 26682 21956 26684
rect 22012 26682 22036 26684
rect 22092 26682 22116 26684
rect 22172 26682 22196 26684
rect 22252 26682 22258 26684
rect 22012 26630 22014 26682
rect 22194 26630 22196 26682
rect 21950 26628 21956 26630
rect 22012 26628 22036 26630
rect 22092 26628 22116 26630
rect 22172 26628 22196 26630
rect 22252 26628 22258 26630
rect 21950 26619 22258 26628
rect 21950 25596 22258 25605
rect 21950 25594 21956 25596
rect 22012 25594 22036 25596
rect 22092 25594 22116 25596
rect 22172 25594 22196 25596
rect 22252 25594 22258 25596
rect 22012 25542 22014 25594
rect 22194 25542 22196 25594
rect 21950 25540 21956 25542
rect 22012 25540 22036 25542
rect 22092 25540 22116 25542
rect 22172 25540 22196 25542
rect 22252 25540 22258 25542
rect 21950 25531 22258 25540
rect 21950 24508 22258 24517
rect 21950 24506 21956 24508
rect 22012 24506 22036 24508
rect 22092 24506 22116 24508
rect 22172 24506 22196 24508
rect 22252 24506 22258 24508
rect 22012 24454 22014 24506
rect 22194 24454 22196 24506
rect 21950 24452 21956 24454
rect 22012 24452 22036 24454
rect 22092 24452 22116 24454
rect 22172 24452 22196 24454
rect 22252 24452 22258 24454
rect 21950 24443 22258 24452
rect 21732 23724 21784 23730
rect 21732 23666 21784 23672
rect 21744 17134 21772 23666
rect 21824 23520 21876 23526
rect 21824 23462 21876 23468
rect 21732 17128 21784 17134
rect 21732 17070 21784 17076
rect 21836 3058 21864 23462
rect 21950 23420 22258 23429
rect 21950 23418 21956 23420
rect 22012 23418 22036 23420
rect 22092 23418 22116 23420
rect 22172 23418 22196 23420
rect 22252 23418 22258 23420
rect 22012 23366 22014 23418
rect 22194 23366 22196 23418
rect 21950 23364 21956 23366
rect 22012 23364 22036 23366
rect 22092 23364 22116 23366
rect 22172 23364 22196 23366
rect 22252 23364 22258 23366
rect 21950 23355 22258 23364
rect 21950 22332 22258 22341
rect 21950 22330 21956 22332
rect 22012 22330 22036 22332
rect 22092 22330 22116 22332
rect 22172 22330 22196 22332
rect 22252 22330 22258 22332
rect 22012 22278 22014 22330
rect 22194 22278 22196 22330
rect 21950 22276 21956 22278
rect 22012 22276 22036 22278
rect 22092 22276 22116 22278
rect 22172 22276 22196 22278
rect 22252 22276 22258 22278
rect 21950 22267 22258 22276
rect 22376 21616 22428 21622
rect 22376 21558 22428 21564
rect 21950 21244 22258 21253
rect 21950 21242 21956 21244
rect 22012 21242 22036 21244
rect 22092 21242 22116 21244
rect 22172 21242 22196 21244
rect 22252 21242 22258 21244
rect 22012 21190 22014 21242
rect 22194 21190 22196 21242
rect 21950 21188 21956 21190
rect 22012 21188 22036 21190
rect 22092 21188 22116 21190
rect 22172 21188 22196 21190
rect 22252 21188 22258 21190
rect 21950 21179 22258 21188
rect 21950 20156 22258 20165
rect 21950 20154 21956 20156
rect 22012 20154 22036 20156
rect 22092 20154 22116 20156
rect 22172 20154 22196 20156
rect 22252 20154 22258 20156
rect 22012 20102 22014 20154
rect 22194 20102 22196 20154
rect 21950 20100 21956 20102
rect 22012 20100 22036 20102
rect 22092 20100 22116 20102
rect 22172 20100 22196 20102
rect 22252 20100 22258 20102
rect 21950 20091 22258 20100
rect 21950 19068 22258 19077
rect 21950 19066 21956 19068
rect 22012 19066 22036 19068
rect 22092 19066 22116 19068
rect 22172 19066 22196 19068
rect 22252 19066 22258 19068
rect 22012 19014 22014 19066
rect 22194 19014 22196 19066
rect 21950 19012 21956 19014
rect 22012 19012 22036 19014
rect 22092 19012 22116 19014
rect 22172 19012 22196 19014
rect 22252 19012 22258 19014
rect 21950 19003 22258 19012
rect 21950 17980 22258 17989
rect 21950 17978 21956 17980
rect 22012 17978 22036 17980
rect 22092 17978 22116 17980
rect 22172 17978 22196 17980
rect 22252 17978 22258 17980
rect 22012 17926 22014 17978
rect 22194 17926 22196 17978
rect 21950 17924 21956 17926
rect 22012 17924 22036 17926
rect 22092 17924 22116 17926
rect 22172 17924 22196 17926
rect 22252 17924 22258 17926
rect 21950 17915 22258 17924
rect 21950 16892 22258 16901
rect 21950 16890 21956 16892
rect 22012 16890 22036 16892
rect 22092 16890 22116 16892
rect 22172 16890 22196 16892
rect 22252 16890 22258 16892
rect 22012 16838 22014 16890
rect 22194 16838 22196 16890
rect 21950 16836 21956 16838
rect 22012 16836 22036 16838
rect 22092 16836 22116 16838
rect 22172 16836 22196 16838
rect 22252 16836 22258 16838
rect 21950 16827 22258 16836
rect 21950 15804 22258 15813
rect 21950 15802 21956 15804
rect 22012 15802 22036 15804
rect 22092 15802 22116 15804
rect 22172 15802 22196 15804
rect 22252 15802 22258 15804
rect 22012 15750 22014 15802
rect 22194 15750 22196 15802
rect 21950 15748 21956 15750
rect 22012 15748 22036 15750
rect 22092 15748 22116 15750
rect 22172 15748 22196 15750
rect 22252 15748 22258 15750
rect 21950 15739 22258 15748
rect 21950 14716 22258 14725
rect 21950 14714 21956 14716
rect 22012 14714 22036 14716
rect 22092 14714 22116 14716
rect 22172 14714 22196 14716
rect 22252 14714 22258 14716
rect 22012 14662 22014 14714
rect 22194 14662 22196 14714
rect 21950 14660 21956 14662
rect 22012 14660 22036 14662
rect 22092 14660 22116 14662
rect 22172 14660 22196 14662
rect 22252 14660 22258 14662
rect 21950 14651 22258 14660
rect 21950 13628 22258 13637
rect 21950 13626 21956 13628
rect 22012 13626 22036 13628
rect 22092 13626 22116 13628
rect 22172 13626 22196 13628
rect 22252 13626 22258 13628
rect 22012 13574 22014 13626
rect 22194 13574 22196 13626
rect 21950 13572 21956 13574
rect 22012 13572 22036 13574
rect 22092 13572 22116 13574
rect 22172 13572 22196 13574
rect 22252 13572 22258 13574
rect 21950 13563 22258 13572
rect 21950 12540 22258 12549
rect 21950 12538 21956 12540
rect 22012 12538 22036 12540
rect 22092 12538 22116 12540
rect 22172 12538 22196 12540
rect 22252 12538 22258 12540
rect 22012 12486 22014 12538
rect 22194 12486 22196 12538
rect 21950 12484 21956 12486
rect 22012 12484 22036 12486
rect 22092 12484 22116 12486
rect 22172 12484 22196 12486
rect 22252 12484 22258 12486
rect 21950 12475 22258 12484
rect 21950 11452 22258 11461
rect 21950 11450 21956 11452
rect 22012 11450 22036 11452
rect 22092 11450 22116 11452
rect 22172 11450 22196 11452
rect 22252 11450 22258 11452
rect 22012 11398 22014 11450
rect 22194 11398 22196 11450
rect 21950 11396 21956 11398
rect 22012 11396 22036 11398
rect 22092 11396 22116 11398
rect 22172 11396 22196 11398
rect 22252 11396 22258 11398
rect 21950 11387 22258 11396
rect 22388 10538 22416 21558
rect 22376 10532 22428 10538
rect 22376 10474 22428 10480
rect 21950 10364 22258 10373
rect 21950 10362 21956 10364
rect 22012 10362 22036 10364
rect 22092 10362 22116 10364
rect 22172 10362 22196 10364
rect 22252 10362 22258 10364
rect 22012 10310 22014 10362
rect 22194 10310 22196 10362
rect 21950 10308 21956 10310
rect 22012 10308 22036 10310
rect 22092 10308 22116 10310
rect 22172 10308 22196 10310
rect 22252 10308 22258 10310
rect 21950 10299 22258 10308
rect 21950 9276 22258 9285
rect 21950 9274 21956 9276
rect 22012 9274 22036 9276
rect 22092 9274 22116 9276
rect 22172 9274 22196 9276
rect 22252 9274 22258 9276
rect 22012 9222 22014 9274
rect 22194 9222 22196 9274
rect 21950 9220 21956 9222
rect 22012 9220 22036 9222
rect 22092 9220 22116 9222
rect 22172 9220 22196 9222
rect 22252 9220 22258 9222
rect 21950 9211 22258 9220
rect 22480 9178 22508 27610
rect 22610 27228 22918 27237
rect 22610 27226 22616 27228
rect 22672 27226 22696 27228
rect 22752 27226 22776 27228
rect 22832 27226 22856 27228
rect 22912 27226 22918 27228
rect 22672 27174 22674 27226
rect 22854 27174 22856 27226
rect 22610 27172 22616 27174
rect 22672 27172 22696 27174
rect 22752 27172 22776 27174
rect 22832 27172 22856 27174
rect 22912 27172 22918 27174
rect 22610 27163 22918 27172
rect 22610 26140 22918 26149
rect 22610 26138 22616 26140
rect 22672 26138 22696 26140
rect 22752 26138 22776 26140
rect 22832 26138 22856 26140
rect 22912 26138 22918 26140
rect 22672 26086 22674 26138
rect 22854 26086 22856 26138
rect 22610 26084 22616 26086
rect 22672 26084 22696 26086
rect 22752 26084 22776 26086
rect 22832 26084 22856 26086
rect 22912 26084 22918 26086
rect 22610 26075 22918 26084
rect 22610 25052 22918 25061
rect 22610 25050 22616 25052
rect 22672 25050 22696 25052
rect 22752 25050 22776 25052
rect 22832 25050 22856 25052
rect 22912 25050 22918 25052
rect 22672 24998 22674 25050
rect 22854 24998 22856 25050
rect 22610 24996 22616 24998
rect 22672 24996 22696 24998
rect 22752 24996 22776 24998
rect 22832 24996 22856 24998
rect 22912 24996 22918 24998
rect 22610 24987 22918 24996
rect 23020 24744 23072 24750
rect 23020 24686 23072 24692
rect 22610 23964 22918 23973
rect 22610 23962 22616 23964
rect 22672 23962 22696 23964
rect 22752 23962 22776 23964
rect 22832 23962 22856 23964
rect 22912 23962 22918 23964
rect 22672 23910 22674 23962
rect 22854 23910 22856 23962
rect 22610 23908 22616 23910
rect 22672 23908 22696 23910
rect 22752 23908 22776 23910
rect 22832 23908 22856 23910
rect 22912 23908 22918 23910
rect 22610 23899 22918 23908
rect 22610 22876 22918 22885
rect 22610 22874 22616 22876
rect 22672 22874 22696 22876
rect 22752 22874 22776 22876
rect 22832 22874 22856 22876
rect 22912 22874 22918 22876
rect 22672 22822 22674 22874
rect 22854 22822 22856 22874
rect 22610 22820 22616 22822
rect 22672 22820 22696 22822
rect 22752 22820 22776 22822
rect 22832 22820 22856 22822
rect 22912 22820 22918 22822
rect 22610 22811 22918 22820
rect 22610 21788 22918 21797
rect 22610 21786 22616 21788
rect 22672 21786 22696 21788
rect 22752 21786 22776 21788
rect 22832 21786 22856 21788
rect 22912 21786 22918 21788
rect 22672 21734 22674 21786
rect 22854 21734 22856 21786
rect 22610 21732 22616 21734
rect 22672 21732 22696 21734
rect 22752 21732 22776 21734
rect 22832 21732 22856 21734
rect 22912 21732 22918 21734
rect 22610 21723 22918 21732
rect 22560 21548 22612 21554
rect 22560 21490 22612 21496
rect 22572 21350 22600 21490
rect 22560 21344 22612 21350
rect 22560 21286 22612 21292
rect 22610 20700 22918 20709
rect 22610 20698 22616 20700
rect 22672 20698 22696 20700
rect 22752 20698 22776 20700
rect 22832 20698 22856 20700
rect 22912 20698 22918 20700
rect 22672 20646 22674 20698
rect 22854 20646 22856 20698
rect 22610 20644 22616 20646
rect 22672 20644 22696 20646
rect 22752 20644 22776 20646
rect 22832 20644 22856 20646
rect 22912 20644 22918 20646
rect 22610 20635 22918 20644
rect 23032 20058 23060 24686
rect 23400 22094 23428 31726
rect 23480 24812 23532 24818
rect 23480 24754 23532 24760
rect 23308 22066 23428 22094
rect 23020 20052 23072 20058
rect 23020 19994 23072 20000
rect 22610 19612 22918 19621
rect 22610 19610 22616 19612
rect 22672 19610 22696 19612
rect 22752 19610 22776 19612
rect 22832 19610 22856 19612
rect 22912 19610 22918 19612
rect 22672 19558 22674 19610
rect 22854 19558 22856 19610
rect 22610 19556 22616 19558
rect 22672 19556 22696 19558
rect 22752 19556 22776 19558
rect 22832 19556 22856 19558
rect 22912 19556 22918 19558
rect 22610 19547 22918 19556
rect 22610 18524 22918 18533
rect 22610 18522 22616 18524
rect 22672 18522 22696 18524
rect 22752 18522 22776 18524
rect 22832 18522 22856 18524
rect 22912 18522 22918 18524
rect 22672 18470 22674 18522
rect 22854 18470 22856 18522
rect 22610 18468 22616 18470
rect 22672 18468 22696 18470
rect 22752 18468 22776 18470
rect 22832 18468 22856 18470
rect 22912 18468 22918 18470
rect 22610 18459 22918 18468
rect 22610 17436 22918 17445
rect 22610 17434 22616 17436
rect 22672 17434 22696 17436
rect 22752 17434 22776 17436
rect 22832 17434 22856 17436
rect 22912 17434 22918 17436
rect 22672 17382 22674 17434
rect 22854 17382 22856 17434
rect 22610 17380 22616 17382
rect 22672 17380 22696 17382
rect 22752 17380 22776 17382
rect 22832 17380 22856 17382
rect 22912 17380 22918 17382
rect 22610 17371 22918 17380
rect 22610 16348 22918 16357
rect 22610 16346 22616 16348
rect 22672 16346 22696 16348
rect 22752 16346 22776 16348
rect 22832 16346 22856 16348
rect 22912 16346 22918 16348
rect 22672 16294 22674 16346
rect 22854 16294 22856 16346
rect 22610 16292 22616 16294
rect 22672 16292 22696 16294
rect 22752 16292 22776 16294
rect 22832 16292 22856 16294
rect 22912 16292 22918 16294
rect 22610 16283 22918 16292
rect 23308 15910 23336 22066
rect 23492 21978 23520 24754
rect 23400 21962 23520 21978
rect 23388 21956 23520 21962
rect 23440 21950 23520 21956
rect 23388 21898 23440 21904
rect 23400 21350 23428 21898
rect 23388 21344 23440 21350
rect 23388 21286 23440 21292
rect 23400 19922 23428 21286
rect 23388 19916 23440 19922
rect 23388 19858 23440 19864
rect 23400 16658 23428 19858
rect 23388 16652 23440 16658
rect 23388 16594 23440 16600
rect 22744 15904 22796 15910
rect 22744 15846 22796 15852
rect 23296 15904 23348 15910
rect 23296 15846 23348 15852
rect 22756 15434 22784 15846
rect 22744 15428 22796 15434
rect 22744 15370 22796 15376
rect 22610 15260 22918 15269
rect 22610 15258 22616 15260
rect 22672 15258 22696 15260
rect 22752 15258 22776 15260
rect 22832 15258 22856 15260
rect 22912 15258 22918 15260
rect 22672 15206 22674 15258
rect 22854 15206 22856 15258
rect 22610 15204 22616 15206
rect 22672 15204 22696 15206
rect 22752 15204 22776 15206
rect 22832 15204 22856 15206
rect 22912 15204 22918 15206
rect 22610 15195 22918 15204
rect 22610 14172 22918 14181
rect 22610 14170 22616 14172
rect 22672 14170 22696 14172
rect 22752 14170 22776 14172
rect 22832 14170 22856 14172
rect 22912 14170 22918 14172
rect 22672 14118 22674 14170
rect 22854 14118 22856 14170
rect 22610 14116 22616 14118
rect 22672 14116 22696 14118
rect 22752 14116 22776 14118
rect 22832 14116 22856 14118
rect 22912 14116 22918 14118
rect 22610 14107 22918 14116
rect 22610 13084 22918 13093
rect 22610 13082 22616 13084
rect 22672 13082 22696 13084
rect 22752 13082 22776 13084
rect 22832 13082 22856 13084
rect 22912 13082 22918 13084
rect 22672 13030 22674 13082
rect 22854 13030 22856 13082
rect 22610 13028 22616 13030
rect 22672 13028 22696 13030
rect 22752 13028 22776 13030
rect 22832 13028 22856 13030
rect 22912 13028 22918 13030
rect 22610 13019 22918 13028
rect 23768 12238 23796 39374
rect 24136 38962 24164 52430
rect 24124 38956 24176 38962
rect 24124 38898 24176 38904
rect 24136 24274 24164 38898
rect 24228 32026 24256 63174
rect 24860 62892 24912 62898
rect 24860 62834 24912 62840
rect 24872 60110 24900 62834
rect 24952 62144 25004 62150
rect 24952 62086 25004 62092
rect 24860 60104 24912 60110
rect 24860 60046 24912 60052
rect 24676 53032 24728 53038
rect 24676 52974 24728 52980
rect 24400 49088 24452 49094
rect 24400 49030 24452 49036
rect 24216 32020 24268 32026
rect 24216 31962 24268 31968
rect 24216 24880 24268 24886
rect 24216 24822 24268 24828
rect 24228 24410 24256 24822
rect 24216 24404 24268 24410
rect 24216 24346 24268 24352
rect 24124 24268 24176 24274
rect 24124 24210 24176 24216
rect 24412 19854 24440 49030
rect 24584 33856 24636 33862
rect 24584 33798 24636 33804
rect 24596 33658 24624 33798
rect 24584 33652 24636 33658
rect 24584 33594 24636 33600
rect 24688 33318 24716 52974
rect 24964 50318 24992 62086
rect 25056 52902 25084 67594
rect 26950 66940 27258 66949
rect 26950 66938 26956 66940
rect 27012 66938 27036 66940
rect 27092 66938 27116 66940
rect 27172 66938 27196 66940
rect 27252 66938 27258 66940
rect 27012 66886 27014 66938
rect 27194 66886 27196 66938
rect 26950 66884 26956 66886
rect 27012 66884 27036 66886
rect 27092 66884 27116 66886
rect 27172 66884 27196 66886
rect 27252 66884 27258 66886
rect 26950 66875 27258 66884
rect 25504 66020 25556 66026
rect 25504 65962 25556 65968
rect 25136 63572 25188 63578
rect 25136 63514 25188 63520
rect 25044 52896 25096 52902
rect 25044 52838 25096 52844
rect 25056 52494 25084 52838
rect 25044 52488 25096 52494
rect 25044 52430 25096 52436
rect 24952 50312 25004 50318
rect 24952 50254 25004 50260
rect 24860 50244 24912 50250
rect 24860 50186 24912 50192
rect 24768 49428 24820 49434
rect 24768 49370 24820 49376
rect 24676 33312 24728 33318
rect 24676 33254 24728 33260
rect 24584 22704 24636 22710
rect 24582 22672 24584 22681
rect 24636 22672 24638 22681
rect 24582 22607 24638 22616
rect 24676 22432 24728 22438
rect 24676 22374 24728 22380
rect 24688 21962 24716 22374
rect 24676 21956 24728 21962
rect 24676 21898 24728 21904
rect 24400 19848 24452 19854
rect 24400 19790 24452 19796
rect 24124 18216 24176 18222
rect 24124 18158 24176 18164
rect 24136 18086 24164 18158
rect 24124 18080 24176 18086
rect 24124 18022 24176 18028
rect 24780 14822 24808 49370
rect 24872 43858 24900 50186
rect 24860 43852 24912 43858
rect 24860 43794 24912 43800
rect 24872 41414 24900 43794
rect 25044 41540 25096 41546
rect 25044 41482 25096 41488
rect 24872 41386 24992 41414
rect 24964 37874 24992 41386
rect 24952 37868 25004 37874
rect 24952 37810 25004 37816
rect 25056 23050 25084 41482
rect 25148 34202 25176 63514
rect 25228 61804 25280 61810
rect 25228 61746 25280 61752
rect 25240 59022 25268 61746
rect 25228 59016 25280 59022
rect 25228 58958 25280 58964
rect 25320 53508 25372 53514
rect 25320 53450 25372 53456
rect 25332 52562 25360 53450
rect 25320 52556 25372 52562
rect 25320 52498 25372 52504
rect 25332 41414 25360 52498
rect 25516 52358 25544 65962
rect 26950 65852 27258 65861
rect 26950 65850 26956 65852
rect 27012 65850 27036 65852
rect 27092 65850 27116 65852
rect 27172 65850 27196 65852
rect 27252 65850 27258 65852
rect 27012 65798 27014 65850
rect 27194 65798 27196 65850
rect 26950 65796 26956 65798
rect 27012 65796 27036 65798
rect 27092 65796 27116 65798
rect 27172 65796 27196 65798
rect 27252 65796 27258 65798
rect 26950 65787 27258 65796
rect 26700 64932 26752 64938
rect 26700 64874 26752 64880
rect 26712 64394 26740 64874
rect 26950 64764 27258 64773
rect 26950 64762 26956 64764
rect 27012 64762 27036 64764
rect 27092 64762 27116 64764
rect 27172 64762 27196 64764
rect 27252 64762 27258 64764
rect 27012 64710 27014 64762
rect 27194 64710 27196 64762
rect 26950 64708 26956 64710
rect 27012 64708 27036 64710
rect 27092 64708 27116 64710
rect 27172 64708 27196 64710
rect 27252 64708 27258 64710
rect 26950 64699 27258 64708
rect 26700 64388 26752 64394
rect 26700 64330 26752 64336
rect 26950 63676 27258 63685
rect 26950 63674 26956 63676
rect 27012 63674 27036 63676
rect 27092 63674 27116 63676
rect 27172 63674 27196 63676
rect 27252 63674 27258 63676
rect 27012 63622 27014 63674
rect 27194 63622 27196 63674
rect 26950 63620 26956 63622
rect 27012 63620 27036 63622
rect 27092 63620 27116 63622
rect 27172 63620 27196 63622
rect 27252 63620 27258 63622
rect 26950 63611 27258 63620
rect 26950 62588 27258 62597
rect 26950 62586 26956 62588
rect 27012 62586 27036 62588
rect 27092 62586 27116 62588
rect 27172 62586 27196 62588
rect 27252 62586 27258 62588
rect 27012 62534 27014 62586
rect 27194 62534 27196 62586
rect 26950 62532 26956 62534
rect 27012 62532 27036 62534
rect 27092 62532 27116 62534
rect 27172 62532 27196 62534
rect 27252 62532 27258 62534
rect 26950 62523 27258 62532
rect 26148 61600 26200 61606
rect 26148 61542 26200 61548
rect 25596 59016 25648 59022
rect 25596 58958 25648 58964
rect 25504 52352 25556 52358
rect 25504 52294 25556 52300
rect 25412 47116 25464 47122
rect 25412 47058 25464 47064
rect 25240 41386 25360 41414
rect 25240 39506 25268 41386
rect 25228 39500 25280 39506
rect 25228 39442 25280 39448
rect 25240 38758 25268 39442
rect 25228 38752 25280 38758
rect 25228 38694 25280 38700
rect 25136 34196 25188 34202
rect 25136 34138 25188 34144
rect 25148 34066 25176 34138
rect 25136 34060 25188 34066
rect 25136 34002 25188 34008
rect 25228 32292 25280 32298
rect 25228 32234 25280 32240
rect 25240 31822 25268 32234
rect 25424 31890 25452 47058
rect 25516 43858 25544 52294
rect 25504 43852 25556 43858
rect 25504 43794 25556 43800
rect 25608 41138 25636 58958
rect 25780 57248 25832 57254
rect 25780 57190 25832 57196
rect 25792 48278 25820 57190
rect 26056 52488 26108 52494
rect 26056 52430 26108 52436
rect 25780 48272 25832 48278
rect 25780 48214 25832 48220
rect 25792 47122 25820 48214
rect 25780 47116 25832 47122
rect 25780 47058 25832 47064
rect 25964 45824 26016 45830
rect 25964 45766 26016 45772
rect 25596 41132 25648 41138
rect 25596 41074 25648 41080
rect 25608 38554 25636 41074
rect 25596 38548 25648 38554
rect 25596 38490 25648 38496
rect 25608 37942 25636 38490
rect 25596 37936 25648 37942
rect 25596 37878 25648 37884
rect 25412 31884 25464 31890
rect 25412 31826 25464 31832
rect 25228 31816 25280 31822
rect 25228 31758 25280 31764
rect 25044 23044 25096 23050
rect 25044 22986 25096 22992
rect 25976 18834 26004 45766
rect 26068 41750 26096 52430
rect 26056 41744 26108 41750
rect 26056 41686 26108 41692
rect 26068 39438 26096 41686
rect 26056 39432 26108 39438
rect 26056 39374 26108 39380
rect 26056 38752 26108 38758
rect 26056 38694 26108 38700
rect 25964 18828 26016 18834
rect 25964 18770 26016 18776
rect 24768 14816 24820 14822
rect 24768 14758 24820 14764
rect 23756 12232 23808 12238
rect 23756 12174 23808 12180
rect 22610 11996 22918 12005
rect 22610 11994 22616 11996
rect 22672 11994 22696 11996
rect 22752 11994 22776 11996
rect 22832 11994 22856 11996
rect 22912 11994 22918 11996
rect 22672 11942 22674 11994
rect 22854 11942 22856 11994
rect 22610 11940 22616 11942
rect 22672 11940 22696 11942
rect 22752 11940 22776 11942
rect 22832 11940 22856 11942
rect 22912 11940 22918 11942
rect 22610 11931 22918 11940
rect 22610 10908 22918 10917
rect 22610 10906 22616 10908
rect 22672 10906 22696 10908
rect 22752 10906 22776 10908
rect 22832 10906 22856 10908
rect 22912 10906 22918 10908
rect 22672 10854 22674 10906
rect 22854 10854 22856 10906
rect 22610 10852 22616 10854
rect 22672 10852 22696 10854
rect 22752 10852 22776 10854
rect 22832 10852 22856 10854
rect 22912 10852 22918 10854
rect 22610 10843 22918 10852
rect 22610 9820 22918 9829
rect 22610 9818 22616 9820
rect 22672 9818 22696 9820
rect 22752 9818 22776 9820
rect 22832 9818 22856 9820
rect 22912 9818 22918 9820
rect 22672 9766 22674 9818
rect 22854 9766 22856 9818
rect 22610 9764 22616 9766
rect 22672 9764 22696 9766
rect 22752 9764 22776 9766
rect 22832 9764 22856 9766
rect 22912 9764 22918 9766
rect 22610 9755 22918 9764
rect 22468 9172 22520 9178
rect 22468 9114 22520 9120
rect 22610 8732 22918 8741
rect 22610 8730 22616 8732
rect 22672 8730 22696 8732
rect 22752 8730 22776 8732
rect 22832 8730 22856 8732
rect 22912 8730 22918 8732
rect 22672 8678 22674 8730
rect 22854 8678 22856 8730
rect 22610 8676 22616 8678
rect 22672 8676 22696 8678
rect 22752 8676 22776 8678
rect 22832 8676 22856 8678
rect 22912 8676 22918 8678
rect 22610 8667 22918 8676
rect 21950 8188 22258 8197
rect 21950 8186 21956 8188
rect 22012 8186 22036 8188
rect 22092 8186 22116 8188
rect 22172 8186 22196 8188
rect 22252 8186 22258 8188
rect 22012 8134 22014 8186
rect 22194 8134 22196 8186
rect 21950 8132 21956 8134
rect 22012 8132 22036 8134
rect 22092 8132 22116 8134
rect 22172 8132 22196 8134
rect 22252 8132 22258 8134
rect 21950 8123 22258 8132
rect 22610 7644 22918 7653
rect 22610 7642 22616 7644
rect 22672 7642 22696 7644
rect 22752 7642 22776 7644
rect 22832 7642 22856 7644
rect 22912 7642 22918 7644
rect 22672 7590 22674 7642
rect 22854 7590 22856 7642
rect 22610 7588 22616 7590
rect 22672 7588 22696 7590
rect 22752 7588 22776 7590
rect 22832 7588 22856 7590
rect 22912 7588 22918 7590
rect 22610 7579 22918 7588
rect 21950 7100 22258 7109
rect 21950 7098 21956 7100
rect 22012 7098 22036 7100
rect 22092 7098 22116 7100
rect 22172 7098 22196 7100
rect 22252 7098 22258 7100
rect 22012 7046 22014 7098
rect 22194 7046 22196 7098
rect 21950 7044 21956 7046
rect 22012 7044 22036 7046
rect 22092 7044 22116 7046
rect 22172 7044 22196 7046
rect 22252 7044 22258 7046
rect 21950 7035 22258 7044
rect 22610 6556 22918 6565
rect 22610 6554 22616 6556
rect 22672 6554 22696 6556
rect 22752 6554 22776 6556
rect 22832 6554 22856 6556
rect 22912 6554 22918 6556
rect 22672 6502 22674 6554
rect 22854 6502 22856 6554
rect 22610 6500 22616 6502
rect 22672 6500 22696 6502
rect 22752 6500 22776 6502
rect 22832 6500 22856 6502
rect 22912 6500 22918 6502
rect 22610 6491 22918 6500
rect 21950 6012 22258 6021
rect 21950 6010 21956 6012
rect 22012 6010 22036 6012
rect 22092 6010 22116 6012
rect 22172 6010 22196 6012
rect 22252 6010 22258 6012
rect 22012 5958 22014 6010
rect 22194 5958 22196 6010
rect 21950 5956 21956 5958
rect 22012 5956 22036 5958
rect 22092 5956 22116 5958
rect 22172 5956 22196 5958
rect 22252 5956 22258 5958
rect 21950 5947 22258 5956
rect 22610 5468 22918 5477
rect 22610 5466 22616 5468
rect 22672 5466 22696 5468
rect 22752 5466 22776 5468
rect 22832 5466 22856 5468
rect 22912 5466 22918 5468
rect 22672 5414 22674 5466
rect 22854 5414 22856 5466
rect 22610 5412 22616 5414
rect 22672 5412 22696 5414
rect 22752 5412 22776 5414
rect 22832 5412 22856 5414
rect 22912 5412 22918 5414
rect 22610 5403 22918 5412
rect 21950 4924 22258 4933
rect 21950 4922 21956 4924
rect 22012 4922 22036 4924
rect 22092 4922 22116 4924
rect 22172 4922 22196 4924
rect 22252 4922 22258 4924
rect 22012 4870 22014 4922
rect 22194 4870 22196 4922
rect 21950 4868 21956 4870
rect 22012 4868 22036 4870
rect 22092 4868 22116 4870
rect 22172 4868 22196 4870
rect 22252 4868 22258 4870
rect 21950 4859 22258 4868
rect 23768 4554 23796 12174
rect 25780 12096 25832 12102
rect 25780 12038 25832 12044
rect 25792 4622 25820 12038
rect 26068 4826 26096 38694
rect 26160 25226 26188 61542
rect 26950 61500 27258 61509
rect 26950 61498 26956 61500
rect 27012 61498 27036 61500
rect 27092 61498 27116 61500
rect 27172 61498 27196 61500
rect 27252 61498 27258 61500
rect 27012 61446 27014 61498
rect 27194 61446 27196 61498
rect 26950 61444 26956 61446
rect 27012 61444 27036 61446
rect 27092 61444 27116 61446
rect 27172 61444 27196 61446
rect 27252 61444 27258 61446
rect 26950 61435 27258 61444
rect 26950 60412 27258 60421
rect 26950 60410 26956 60412
rect 27012 60410 27036 60412
rect 27092 60410 27116 60412
rect 27172 60410 27196 60412
rect 27252 60410 27258 60412
rect 27012 60358 27014 60410
rect 27194 60358 27196 60410
rect 26950 60356 26956 60358
rect 27012 60356 27036 60358
rect 27092 60356 27116 60358
rect 27172 60356 27196 60358
rect 27252 60356 27258 60358
rect 26950 60347 27258 60356
rect 26950 59324 27258 59333
rect 26950 59322 26956 59324
rect 27012 59322 27036 59324
rect 27092 59322 27116 59324
rect 27172 59322 27196 59324
rect 27252 59322 27258 59324
rect 27012 59270 27014 59322
rect 27194 59270 27196 59322
rect 26950 59268 26956 59270
rect 27012 59268 27036 59270
rect 27092 59268 27116 59270
rect 27172 59268 27196 59270
rect 27252 59268 27258 59270
rect 26950 59259 27258 59268
rect 26950 58236 27258 58245
rect 26950 58234 26956 58236
rect 27012 58234 27036 58236
rect 27092 58234 27116 58236
rect 27172 58234 27196 58236
rect 27252 58234 27258 58236
rect 27012 58182 27014 58234
rect 27194 58182 27196 58234
rect 26950 58180 26956 58182
rect 27012 58180 27036 58182
rect 27092 58180 27116 58182
rect 27172 58180 27196 58182
rect 27252 58180 27258 58182
rect 26950 58171 27258 58180
rect 26950 57148 27258 57157
rect 26950 57146 26956 57148
rect 27012 57146 27036 57148
rect 27092 57146 27116 57148
rect 27172 57146 27196 57148
rect 27252 57146 27258 57148
rect 27012 57094 27014 57146
rect 27194 57094 27196 57146
rect 26950 57092 26956 57094
rect 27012 57092 27036 57094
rect 27092 57092 27116 57094
rect 27172 57092 27196 57094
rect 27252 57092 27258 57094
rect 26950 57083 27258 57092
rect 26950 56060 27258 56069
rect 26950 56058 26956 56060
rect 27012 56058 27036 56060
rect 27092 56058 27116 56060
rect 27172 56058 27196 56060
rect 27252 56058 27258 56060
rect 27012 56006 27014 56058
rect 27194 56006 27196 56058
rect 26950 56004 26956 56006
rect 27012 56004 27036 56006
rect 27092 56004 27116 56006
rect 27172 56004 27196 56006
rect 27252 56004 27258 56006
rect 26950 55995 27258 56004
rect 26950 54972 27258 54981
rect 26950 54970 26956 54972
rect 27012 54970 27036 54972
rect 27092 54970 27116 54972
rect 27172 54970 27196 54972
rect 27252 54970 27258 54972
rect 27012 54918 27014 54970
rect 27194 54918 27196 54970
rect 26950 54916 26956 54918
rect 27012 54916 27036 54918
rect 27092 54916 27116 54918
rect 27172 54916 27196 54918
rect 27252 54916 27258 54918
rect 26950 54907 27258 54916
rect 26950 53884 27258 53893
rect 26950 53882 26956 53884
rect 27012 53882 27036 53884
rect 27092 53882 27116 53884
rect 27172 53882 27196 53884
rect 27252 53882 27258 53884
rect 27012 53830 27014 53882
rect 27194 53830 27196 53882
rect 26950 53828 26956 53830
rect 27012 53828 27036 53830
rect 27092 53828 27116 53830
rect 27172 53828 27196 53830
rect 27252 53828 27258 53830
rect 26950 53819 27258 53828
rect 26950 52796 27258 52805
rect 26950 52794 26956 52796
rect 27012 52794 27036 52796
rect 27092 52794 27116 52796
rect 27172 52794 27196 52796
rect 27252 52794 27258 52796
rect 27012 52742 27014 52794
rect 27194 52742 27196 52794
rect 26950 52740 26956 52742
rect 27012 52740 27036 52742
rect 27092 52740 27116 52742
rect 27172 52740 27196 52742
rect 27252 52740 27258 52742
rect 26950 52731 27258 52740
rect 26950 51708 27258 51717
rect 26950 51706 26956 51708
rect 27012 51706 27036 51708
rect 27092 51706 27116 51708
rect 27172 51706 27196 51708
rect 27252 51706 27258 51708
rect 27012 51654 27014 51706
rect 27194 51654 27196 51706
rect 26950 51652 26956 51654
rect 27012 51652 27036 51654
rect 27092 51652 27116 51654
rect 27172 51652 27196 51654
rect 27252 51652 27258 51654
rect 26950 51643 27258 51652
rect 26950 50620 27258 50629
rect 26950 50618 26956 50620
rect 27012 50618 27036 50620
rect 27092 50618 27116 50620
rect 27172 50618 27196 50620
rect 27252 50618 27258 50620
rect 27012 50566 27014 50618
rect 27194 50566 27196 50618
rect 26950 50564 26956 50566
rect 27012 50564 27036 50566
rect 27092 50564 27116 50566
rect 27172 50564 27196 50566
rect 27252 50564 27258 50566
rect 26950 50555 27258 50564
rect 26950 49532 27258 49541
rect 26950 49530 26956 49532
rect 27012 49530 27036 49532
rect 27092 49530 27116 49532
rect 27172 49530 27196 49532
rect 27252 49530 27258 49532
rect 27012 49478 27014 49530
rect 27194 49478 27196 49530
rect 26950 49476 26956 49478
rect 27012 49476 27036 49478
rect 27092 49476 27116 49478
rect 27172 49476 27196 49478
rect 27252 49476 27258 49478
rect 26950 49467 27258 49476
rect 26516 49156 26568 49162
rect 26516 49098 26568 49104
rect 26528 48346 26556 49098
rect 26950 48444 27258 48453
rect 26950 48442 26956 48444
rect 27012 48442 27036 48444
rect 27092 48442 27116 48444
rect 27172 48442 27196 48444
rect 27252 48442 27258 48444
rect 27012 48390 27014 48442
rect 27194 48390 27196 48442
rect 26950 48388 26956 48390
rect 27012 48388 27036 48390
rect 27092 48388 27116 48390
rect 27172 48388 27196 48390
rect 27252 48388 27258 48390
rect 26950 48379 27258 48388
rect 26516 48340 26568 48346
rect 26516 48282 26568 48288
rect 26528 45898 26556 48282
rect 26950 47356 27258 47365
rect 26950 47354 26956 47356
rect 27012 47354 27036 47356
rect 27092 47354 27116 47356
rect 27172 47354 27196 47356
rect 27252 47354 27258 47356
rect 27012 47302 27014 47354
rect 27194 47302 27196 47354
rect 26950 47300 26956 47302
rect 27012 47300 27036 47302
rect 27092 47300 27116 47302
rect 27172 47300 27196 47302
rect 27252 47300 27258 47302
rect 26950 47291 27258 47300
rect 26950 46268 27258 46277
rect 26950 46266 26956 46268
rect 27012 46266 27036 46268
rect 27092 46266 27116 46268
rect 27172 46266 27196 46268
rect 27252 46266 27258 46268
rect 27012 46214 27014 46266
rect 27194 46214 27196 46266
rect 26950 46212 26956 46214
rect 27012 46212 27036 46214
rect 27092 46212 27116 46214
rect 27172 46212 27196 46214
rect 27252 46212 27258 46214
rect 26950 46203 27258 46212
rect 26516 45892 26568 45898
rect 26516 45834 26568 45840
rect 26950 45180 27258 45189
rect 26950 45178 26956 45180
rect 27012 45178 27036 45180
rect 27092 45178 27116 45180
rect 27172 45178 27196 45180
rect 27252 45178 27258 45180
rect 27012 45126 27014 45178
rect 27194 45126 27196 45178
rect 26950 45124 26956 45126
rect 27012 45124 27036 45126
rect 27092 45124 27116 45126
rect 27172 45124 27196 45126
rect 27252 45124 27258 45126
rect 26950 45115 27258 45124
rect 26950 44092 27258 44101
rect 26950 44090 26956 44092
rect 27012 44090 27036 44092
rect 27092 44090 27116 44092
rect 27172 44090 27196 44092
rect 27252 44090 27258 44092
rect 27012 44038 27014 44090
rect 27194 44038 27196 44090
rect 26950 44036 26956 44038
rect 27012 44036 27036 44038
rect 27092 44036 27116 44038
rect 27172 44036 27196 44038
rect 27252 44036 27258 44038
rect 26950 44027 27258 44036
rect 26950 43004 27258 43013
rect 26950 43002 26956 43004
rect 27012 43002 27036 43004
rect 27092 43002 27116 43004
rect 27172 43002 27196 43004
rect 27252 43002 27258 43004
rect 27012 42950 27014 43002
rect 27194 42950 27196 43002
rect 26950 42948 26956 42950
rect 27012 42948 27036 42950
rect 27092 42948 27116 42950
rect 27172 42948 27196 42950
rect 27252 42948 27258 42950
rect 26950 42939 27258 42948
rect 26950 41916 27258 41925
rect 26950 41914 26956 41916
rect 27012 41914 27036 41916
rect 27092 41914 27116 41916
rect 27172 41914 27196 41916
rect 27252 41914 27258 41916
rect 27012 41862 27014 41914
rect 27194 41862 27196 41914
rect 26950 41860 26956 41862
rect 27012 41860 27036 41862
rect 27092 41860 27116 41862
rect 27172 41860 27196 41862
rect 27252 41860 27258 41862
rect 26950 41851 27258 41860
rect 26344 41546 26740 41562
rect 26332 41540 26752 41546
rect 26384 41534 26700 41540
rect 26332 41482 26384 41488
rect 26700 41482 26752 41488
rect 26950 40828 27258 40837
rect 26950 40826 26956 40828
rect 27012 40826 27036 40828
rect 27092 40826 27116 40828
rect 27172 40826 27196 40828
rect 27252 40826 27258 40828
rect 27012 40774 27014 40826
rect 27194 40774 27196 40826
rect 26950 40772 26956 40774
rect 27012 40772 27036 40774
rect 27092 40772 27116 40774
rect 27172 40772 27196 40774
rect 27252 40772 27258 40774
rect 26950 40763 27258 40772
rect 26950 39740 27258 39749
rect 26950 39738 26956 39740
rect 27012 39738 27036 39740
rect 27092 39738 27116 39740
rect 27172 39738 27196 39740
rect 27252 39738 27258 39740
rect 27012 39686 27014 39738
rect 27194 39686 27196 39738
rect 26950 39684 26956 39686
rect 27012 39684 27036 39686
rect 27092 39684 27116 39686
rect 27172 39684 27196 39686
rect 27252 39684 27258 39686
rect 26950 39675 27258 39684
rect 26950 38652 27258 38661
rect 26950 38650 26956 38652
rect 27012 38650 27036 38652
rect 27092 38650 27116 38652
rect 27172 38650 27196 38652
rect 27252 38650 27258 38652
rect 27012 38598 27014 38650
rect 27194 38598 27196 38650
rect 26950 38596 26956 38598
rect 27012 38596 27036 38598
rect 27092 38596 27116 38598
rect 27172 38596 27196 38598
rect 27252 38596 27258 38598
rect 26950 38587 27258 38596
rect 26792 38548 26844 38554
rect 26792 38490 26844 38496
rect 26804 36786 26832 38490
rect 26950 37564 27258 37573
rect 26950 37562 26956 37564
rect 27012 37562 27036 37564
rect 27092 37562 27116 37564
rect 27172 37562 27196 37564
rect 27252 37562 27258 37564
rect 27012 37510 27014 37562
rect 27194 37510 27196 37562
rect 26950 37508 26956 37510
rect 27012 37508 27036 37510
rect 27092 37508 27116 37510
rect 27172 37508 27196 37510
rect 27252 37508 27258 37510
rect 26950 37499 27258 37508
rect 26792 36780 26844 36786
rect 26792 36722 26844 36728
rect 26804 29102 26832 36722
rect 26950 36476 27258 36485
rect 26950 36474 26956 36476
rect 27012 36474 27036 36476
rect 27092 36474 27116 36476
rect 27172 36474 27196 36476
rect 27252 36474 27258 36476
rect 27012 36422 27014 36474
rect 27194 36422 27196 36474
rect 26950 36420 26956 36422
rect 27012 36420 27036 36422
rect 27092 36420 27116 36422
rect 27172 36420 27196 36422
rect 27252 36420 27258 36422
rect 26950 36411 27258 36420
rect 26950 35388 27258 35397
rect 26950 35386 26956 35388
rect 27012 35386 27036 35388
rect 27092 35386 27116 35388
rect 27172 35386 27196 35388
rect 27252 35386 27258 35388
rect 27012 35334 27014 35386
rect 27194 35334 27196 35386
rect 26950 35332 26956 35334
rect 27012 35332 27036 35334
rect 27092 35332 27116 35334
rect 27172 35332 27196 35334
rect 27252 35332 27258 35334
rect 26950 35323 27258 35332
rect 26950 34300 27258 34309
rect 26950 34298 26956 34300
rect 27012 34298 27036 34300
rect 27092 34298 27116 34300
rect 27172 34298 27196 34300
rect 27252 34298 27258 34300
rect 27012 34246 27014 34298
rect 27194 34246 27196 34298
rect 26950 34244 26956 34246
rect 27012 34244 27036 34246
rect 27092 34244 27116 34246
rect 27172 34244 27196 34246
rect 27252 34244 27258 34246
rect 26950 34235 27258 34244
rect 26950 33212 27258 33221
rect 26950 33210 26956 33212
rect 27012 33210 27036 33212
rect 27092 33210 27116 33212
rect 27172 33210 27196 33212
rect 27252 33210 27258 33212
rect 27012 33158 27014 33210
rect 27194 33158 27196 33210
rect 26950 33156 26956 33158
rect 27012 33156 27036 33158
rect 27092 33156 27116 33158
rect 27172 33156 27196 33158
rect 27252 33156 27258 33158
rect 26950 33147 27258 33156
rect 26950 32124 27258 32133
rect 26950 32122 26956 32124
rect 27012 32122 27036 32124
rect 27092 32122 27116 32124
rect 27172 32122 27196 32124
rect 27252 32122 27258 32124
rect 27012 32070 27014 32122
rect 27194 32070 27196 32122
rect 26950 32068 26956 32070
rect 27012 32068 27036 32070
rect 27092 32068 27116 32070
rect 27172 32068 27196 32070
rect 27252 32068 27258 32070
rect 26950 32059 27258 32068
rect 26950 31036 27258 31045
rect 26950 31034 26956 31036
rect 27012 31034 27036 31036
rect 27092 31034 27116 31036
rect 27172 31034 27196 31036
rect 27252 31034 27258 31036
rect 27012 30982 27014 31034
rect 27194 30982 27196 31034
rect 26950 30980 26956 30982
rect 27012 30980 27036 30982
rect 27092 30980 27116 30982
rect 27172 30980 27196 30982
rect 27252 30980 27258 30982
rect 26950 30971 27258 30980
rect 26950 29948 27258 29957
rect 26950 29946 26956 29948
rect 27012 29946 27036 29948
rect 27092 29946 27116 29948
rect 27172 29946 27196 29948
rect 27252 29946 27258 29948
rect 27012 29894 27014 29946
rect 27194 29894 27196 29946
rect 26950 29892 26956 29894
rect 27012 29892 27036 29894
rect 27092 29892 27116 29894
rect 27172 29892 27196 29894
rect 27252 29892 27258 29894
rect 26950 29883 27258 29892
rect 26792 29096 26844 29102
rect 26792 29038 26844 29044
rect 26950 28860 27258 28869
rect 26950 28858 26956 28860
rect 27012 28858 27036 28860
rect 27092 28858 27116 28860
rect 27172 28858 27196 28860
rect 27252 28858 27258 28860
rect 27012 28806 27014 28858
rect 27194 28806 27196 28858
rect 26950 28804 26956 28806
rect 27012 28804 27036 28806
rect 27092 28804 27116 28806
rect 27172 28804 27196 28806
rect 27252 28804 27258 28806
rect 26950 28795 27258 28804
rect 26950 27772 27258 27781
rect 26950 27770 26956 27772
rect 27012 27770 27036 27772
rect 27092 27770 27116 27772
rect 27172 27770 27196 27772
rect 27252 27770 27258 27772
rect 27012 27718 27014 27770
rect 27194 27718 27196 27770
rect 26950 27716 26956 27718
rect 27012 27716 27036 27718
rect 27092 27716 27116 27718
rect 27172 27716 27196 27718
rect 27252 27716 27258 27718
rect 26950 27707 27258 27716
rect 26950 26684 27258 26693
rect 26950 26682 26956 26684
rect 27012 26682 27036 26684
rect 27092 26682 27116 26684
rect 27172 26682 27196 26684
rect 27252 26682 27258 26684
rect 27012 26630 27014 26682
rect 27194 26630 27196 26682
rect 26950 26628 26956 26630
rect 27012 26628 27036 26630
rect 27092 26628 27116 26630
rect 27172 26628 27196 26630
rect 27252 26628 27258 26630
rect 26950 26619 27258 26628
rect 26950 25596 27258 25605
rect 26950 25594 26956 25596
rect 27012 25594 27036 25596
rect 27092 25594 27116 25596
rect 27172 25594 27196 25596
rect 27252 25594 27258 25596
rect 27012 25542 27014 25594
rect 27194 25542 27196 25594
rect 26950 25540 26956 25542
rect 27012 25540 27036 25542
rect 27092 25540 27116 25542
rect 27172 25540 27196 25542
rect 27252 25540 27258 25542
rect 26950 25531 27258 25540
rect 26148 25220 26200 25226
rect 26148 25162 26200 25168
rect 26950 24508 27258 24517
rect 26950 24506 26956 24508
rect 27012 24506 27036 24508
rect 27092 24506 27116 24508
rect 27172 24506 27196 24508
rect 27252 24506 27258 24508
rect 27012 24454 27014 24506
rect 27194 24454 27196 24506
rect 26950 24452 26956 24454
rect 27012 24452 27036 24454
rect 27092 24452 27116 24454
rect 27172 24452 27196 24454
rect 27252 24452 27258 24454
rect 26950 24443 27258 24452
rect 27356 24342 27384 69362
rect 31950 69116 32258 69125
rect 31950 69114 31956 69116
rect 32012 69114 32036 69116
rect 32092 69114 32116 69116
rect 32172 69114 32196 69116
rect 32252 69114 32258 69116
rect 32012 69062 32014 69114
rect 32194 69062 32196 69114
rect 31950 69060 31956 69062
rect 32012 69060 32036 69062
rect 32092 69060 32116 69062
rect 32172 69060 32196 69062
rect 32252 69060 32258 69062
rect 31950 69051 32258 69060
rect 27610 68572 27918 68581
rect 27610 68570 27616 68572
rect 27672 68570 27696 68572
rect 27752 68570 27776 68572
rect 27832 68570 27856 68572
rect 27912 68570 27918 68572
rect 27672 68518 27674 68570
rect 27854 68518 27856 68570
rect 27610 68516 27616 68518
rect 27672 68516 27696 68518
rect 27752 68516 27776 68518
rect 27832 68516 27856 68518
rect 27912 68516 27918 68518
rect 27610 68507 27918 68516
rect 32610 68572 32918 68581
rect 32610 68570 32616 68572
rect 32672 68570 32696 68572
rect 32752 68570 32776 68572
rect 32832 68570 32856 68572
rect 32912 68570 32918 68572
rect 32672 68518 32674 68570
rect 32854 68518 32856 68570
rect 32610 68516 32616 68518
rect 32672 68516 32696 68518
rect 32752 68516 32776 68518
rect 32832 68516 32856 68518
rect 32912 68516 32918 68518
rect 32610 68507 32918 68516
rect 29092 68400 29144 68406
rect 29092 68342 29144 68348
rect 27610 67484 27918 67493
rect 27610 67482 27616 67484
rect 27672 67482 27696 67484
rect 27752 67482 27776 67484
rect 27832 67482 27856 67484
rect 27912 67482 27918 67484
rect 27672 67430 27674 67482
rect 27854 67430 27856 67482
rect 27610 67428 27616 67430
rect 27672 67428 27696 67430
rect 27752 67428 27776 67430
rect 27832 67428 27856 67430
rect 27912 67428 27918 67430
rect 27610 67419 27918 67428
rect 27610 66396 27918 66405
rect 27610 66394 27616 66396
rect 27672 66394 27696 66396
rect 27752 66394 27776 66396
rect 27832 66394 27856 66396
rect 27912 66394 27918 66396
rect 27672 66342 27674 66394
rect 27854 66342 27856 66394
rect 27610 66340 27616 66342
rect 27672 66340 27696 66342
rect 27752 66340 27776 66342
rect 27832 66340 27856 66342
rect 27912 66340 27918 66342
rect 27610 66331 27918 66340
rect 27610 65308 27918 65317
rect 27610 65306 27616 65308
rect 27672 65306 27696 65308
rect 27752 65306 27776 65308
rect 27832 65306 27856 65308
rect 27912 65306 27918 65308
rect 27672 65254 27674 65306
rect 27854 65254 27856 65306
rect 27610 65252 27616 65254
rect 27672 65252 27696 65254
rect 27752 65252 27776 65254
rect 27832 65252 27856 65254
rect 27912 65252 27918 65254
rect 27610 65243 27918 65252
rect 27528 64320 27580 64326
rect 27528 64262 27580 64268
rect 27436 63912 27488 63918
rect 27436 63854 27488 63860
rect 27448 55418 27476 63854
rect 27436 55412 27488 55418
rect 27436 55354 27488 55360
rect 27436 53576 27488 53582
rect 27436 53518 27488 53524
rect 27448 36922 27476 53518
rect 27540 51950 27568 64262
rect 27610 64220 27918 64229
rect 27610 64218 27616 64220
rect 27672 64218 27696 64220
rect 27752 64218 27776 64220
rect 27832 64218 27856 64220
rect 27912 64218 27918 64220
rect 27672 64166 27674 64218
rect 27854 64166 27856 64218
rect 27610 64164 27616 64166
rect 27672 64164 27696 64166
rect 27752 64164 27776 64166
rect 27832 64164 27856 64166
rect 27912 64164 27918 64166
rect 27610 64155 27918 64164
rect 27610 63132 27918 63141
rect 27610 63130 27616 63132
rect 27672 63130 27696 63132
rect 27752 63130 27776 63132
rect 27832 63130 27856 63132
rect 27912 63130 27918 63132
rect 27672 63078 27674 63130
rect 27854 63078 27856 63130
rect 27610 63076 27616 63078
rect 27672 63076 27696 63078
rect 27752 63076 27776 63078
rect 27832 63076 27856 63078
rect 27912 63076 27918 63078
rect 27610 63067 27918 63076
rect 27610 62044 27918 62053
rect 27610 62042 27616 62044
rect 27672 62042 27696 62044
rect 27752 62042 27776 62044
rect 27832 62042 27856 62044
rect 27912 62042 27918 62044
rect 27672 61990 27674 62042
rect 27854 61990 27856 62042
rect 27610 61988 27616 61990
rect 27672 61988 27696 61990
rect 27752 61988 27776 61990
rect 27832 61988 27856 61990
rect 27912 61988 27918 61990
rect 27610 61979 27918 61988
rect 27610 60956 27918 60965
rect 27610 60954 27616 60956
rect 27672 60954 27696 60956
rect 27752 60954 27776 60956
rect 27832 60954 27856 60956
rect 27912 60954 27918 60956
rect 27672 60902 27674 60954
rect 27854 60902 27856 60954
rect 27610 60900 27616 60902
rect 27672 60900 27696 60902
rect 27752 60900 27776 60902
rect 27832 60900 27856 60902
rect 27912 60900 27918 60902
rect 27610 60891 27918 60900
rect 27610 59868 27918 59877
rect 27610 59866 27616 59868
rect 27672 59866 27696 59868
rect 27752 59866 27776 59868
rect 27832 59866 27856 59868
rect 27912 59866 27918 59868
rect 27672 59814 27674 59866
rect 27854 59814 27856 59866
rect 27610 59812 27616 59814
rect 27672 59812 27696 59814
rect 27752 59812 27776 59814
rect 27832 59812 27856 59814
rect 27912 59812 27918 59814
rect 27610 59803 27918 59812
rect 27610 58780 27918 58789
rect 27610 58778 27616 58780
rect 27672 58778 27696 58780
rect 27752 58778 27776 58780
rect 27832 58778 27856 58780
rect 27912 58778 27918 58780
rect 27672 58726 27674 58778
rect 27854 58726 27856 58778
rect 27610 58724 27616 58726
rect 27672 58724 27696 58726
rect 27752 58724 27776 58726
rect 27832 58724 27856 58726
rect 27912 58724 27918 58726
rect 27610 58715 27918 58724
rect 27610 57692 27918 57701
rect 27610 57690 27616 57692
rect 27672 57690 27696 57692
rect 27752 57690 27776 57692
rect 27832 57690 27856 57692
rect 27912 57690 27918 57692
rect 27672 57638 27674 57690
rect 27854 57638 27856 57690
rect 27610 57636 27616 57638
rect 27672 57636 27696 57638
rect 27752 57636 27776 57638
rect 27832 57636 27856 57638
rect 27912 57636 27918 57638
rect 27610 57627 27918 57636
rect 27610 56604 27918 56613
rect 27610 56602 27616 56604
rect 27672 56602 27696 56604
rect 27752 56602 27776 56604
rect 27832 56602 27856 56604
rect 27912 56602 27918 56604
rect 27672 56550 27674 56602
rect 27854 56550 27856 56602
rect 27610 56548 27616 56550
rect 27672 56548 27696 56550
rect 27752 56548 27776 56550
rect 27832 56548 27856 56550
rect 27912 56548 27918 56550
rect 27610 56539 27918 56548
rect 28540 56432 28592 56438
rect 28540 56374 28592 56380
rect 29000 56432 29052 56438
rect 29000 56374 29052 56380
rect 28552 56166 28580 56374
rect 28540 56160 28592 56166
rect 28540 56102 28592 56108
rect 28632 56160 28684 56166
rect 28632 56102 28684 56108
rect 27610 55516 27918 55525
rect 27610 55514 27616 55516
rect 27672 55514 27696 55516
rect 27752 55514 27776 55516
rect 27832 55514 27856 55516
rect 27912 55514 27918 55516
rect 27672 55462 27674 55514
rect 27854 55462 27856 55514
rect 27610 55460 27616 55462
rect 27672 55460 27696 55462
rect 27752 55460 27776 55462
rect 27832 55460 27856 55462
rect 27912 55460 27918 55462
rect 27610 55451 27918 55460
rect 27610 54428 27918 54437
rect 27610 54426 27616 54428
rect 27672 54426 27696 54428
rect 27752 54426 27776 54428
rect 27832 54426 27856 54428
rect 27912 54426 27918 54428
rect 27672 54374 27674 54426
rect 27854 54374 27856 54426
rect 27610 54372 27616 54374
rect 27672 54372 27696 54374
rect 27752 54372 27776 54374
rect 27832 54372 27856 54374
rect 27912 54372 27918 54374
rect 27610 54363 27918 54372
rect 27610 53340 27918 53349
rect 27610 53338 27616 53340
rect 27672 53338 27696 53340
rect 27752 53338 27776 53340
rect 27832 53338 27856 53340
rect 27912 53338 27918 53340
rect 27672 53286 27674 53338
rect 27854 53286 27856 53338
rect 27610 53284 27616 53286
rect 27672 53284 27696 53286
rect 27752 53284 27776 53286
rect 27832 53284 27856 53286
rect 27912 53284 27918 53286
rect 27610 53275 27918 53284
rect 28552 52426 28580 56102
rect 28644 55622 28672 56102
rect 28632 55616 28684 55622
rect 28632 55558 28684 55564
rect 28540 52420 28592 52426
rect 28540 52362 28592 52368
rect 27610 52252 27918 52261
rect 27610 52250 27616 52252
rect 27672 52250 27696 52252
rect 27752 52250 27776 52252
rect 27832 52250 27856 52252
rect 27912 52250 27918 52252
rect 27672 52198 27674 52250
rect 27854 52198 27856 52250
rect 27610 52196 27616 52198
rect 27672 52196 27696 52198
rect 27752 52196 27776 52198
rect 27832 52196 27856 52198
rect 27912 52196 27918 52198
rect 27610 52187 27918 52196
rect 27528 51944 27580 51950
rect 27528 51886 27580 51892
rect 27610 51164 27918 51173
rect 27610 51162 27616 51164
rect 27672 51162 27696 51164
rect 27752 51162 27776 51164
rect 27832 51162 27856 51164
rect 27912 51162 27918 51164
rect 27672 51110 27674 51162
rect 27854 51110 27856 51162
rect 27610 51108 27616 51110
rect 27672 51108 27696 51110
rect 27752 51108 27776 51110
rect 27832 51108 27856 51110
rect 27912 51108 27918 51110
rect 27610 51099 27918 51108
rect 27610 50076 27918 50085
rect 27610 50074 27616 50076
rect 27672 50074 27696 50076
rect 27752 50074 27776 50076
rect 27832 50074 27856 50076
rect 27912 50074 27918 50076
rect 27672 50022 27674 50074
rect 27854 50022 27856 50074
rect 27610 50020 27616 50022
rect 27672 50020 27696 50022
rect 27752 50020 27776 50022
rect 27832 50020 27856 50022
rect 27912 50020 27918 50022
rect 27610 50011 27918 50020
rect 27610 48988 27918 48997
rect 27610 48986 27616 48988
rect 27672 48986 27696 48988
rect 27752 48986 27776 48988
rect 27832 48986 27856 48988
rect 27912 48986 27918 48988
rect 27672 48934 27674 48986
rect 27854 48934 27856 48986
rect 27610 48932 27616 48934
rect 27672 48932 27696 48934
rect 27752 48932 27776 48934
rect 27832 48932 27856 48934
rect 27912 48932 27918 48934
rect 27610 48923 27918 48932
rect 27610 47900 27918 47909
rect 27610 47898 27616 47900
rect 27672 47898 27696 47900
rect 27752 47898 27776 47900
rect 27832 47898 27856 47900
rect 27912 47898 27918 47900
rect 27672 47846 27674 47898
rect 27854 47846 27856 47898
rect 27610 47844 27616 47846
rect 27672 47844 27696 47846
rect 27752 47844 27776 47846
rect 27832 47844 27856 47846
rect 27912 47844 27918 47846
rect 27610 47835 27918 47844
rect 27610 46812 27918 46821
rect 27610 46810 27616 46812
rect 27672 46810 27696 46812
rect 27752 46810 27776 46812
rect 27832 46810 27856 46812
rect 27912 46810 27918 46812
rect 27672 46758 27674 46810
rect 27854 46758 27856 46810
rect 27610 46756 27616 46758
rect 27672 46756 27696 46758
rect 27752 46756 27776 46758
rect 27832 46756 27856 46758
rect 27912 46756 27918 46758
rect 27610 46747 27918 46756
rect 27610 45724 27918 45733
rect 27610 45722 27616 45724
rect 27672 45722 27696 45724
rect 27752 45722 27776 45724
rect 27832 45722 27856 45724
rect 27912 45722 27918 45724
rect 27672 45670 27674 45722
rect 27854 45670 27856 45722
rect 27610 45668 27616 45670
rect 27672 45668 27696 45670
rect 27752 45668 27776 45670
rect 27832 45668 27856 45670
rect 27912 45668 27918 45670
rect 27610 45659 27918 45668
rect 27610 44636 27918 44645
rect 27610 44634 27616 44636
rect 27672 44634 27696 44636
rect 27752 44634 27776 44636
rect 27832 44634 27856 44636
rect 27912 44634 27918 44636
rect 27672 44582 27674 44634
rect 27854 44582 27856 44634
rect 27610 44580 27616 44582
rect 27672 44580 27696 44582
rect 27752 44580 27776 44582
rect 27832 44580 27856 44582
rect 27912 44580 27918 44582
rect 27610 44571 27918 44580
rect 28264 43784 28316 43790
rect 28264 43726 28316 43732
rect 27610 43548 27918 43557
rect 27610 43546 27616 43548
rect 27672 43546 27696 43548
rect 27752 43546 27776 43548
rect 27832 43546 27856 43548
rect 27912 43546 27918 43548
rect 27672 43494 27674 43546
rect 27854 43494 27856 43546
rect 27610 43492 27616 43494
rect 27672 43492 27696 43494
rect 27752 43492 27776 43494
rect 27832 43492 27856 43494
rect 27912 43492 27918 43494
rect 27610 43483 27918 43492
rect 27610 42460 27918 42469
rect 27610 42458 27616 42460
rect 27672 42458 27696 42460
rect 27752 42458 27776 42460
rect 27832 42458 27856 42460
rect 27912 42458 27918 42460
rect 27672 42406 27674 42458
rect 27854 42406 27856 42458
rect 27610 42404 27616 42406
rect 27672 42404 27696 42406
rect 27752 42404 27776 42406
rect 27832 42404 27856 42406
rect 27912 42404 27918 42406
rect 27610 42395 27918 42404
rect 27988 41540 28040 41546
rect 27988 41482 28040 41488
rect 27610 41372 27918 41381
rect 27610 41370 27616 41372
rect 27672 41370 27696 41372
rect 27752 41370 27776 41372
rect 27832 41370 27856 41372
rect 27912 41370 27918 41372
rect 27672 41318 27674 41370
rect 27854 41318 27856 41370
rect 27610 41316 27616 41318
rect 27672 41316 27696 41318
rect 27752 41316 27776 41318
rect 27832 41316 27856 41318
rect 27912 41316 27918 41318
rect 27610 41307 27918 41316
rect 27610 40284 27918 40293
rect 27610 40282 27616 40284
rect 27672 40282 27696 40284
rect 27752 40282 27776 40284
rect 27832 40282 27856 40284
rect 27912 40282 27918 40284
rect 27672 40230 27674 40282
rect 27854 40230 27856 40282
rect 27610 40228 27616 40230
rect 27672 40228 27696 40230
rect 27752 40228 27776 40230
rect 27832 40228 27856 40230
rect 27912 40228 27918 40230
rect 27610 40219 27918 40228
rect 27610 39196 27918 39205
rect 27610 39194 27616 39196
rect 27672 39194 27696 39196
rect 27752 39194 27776 39196
rect 27832 39194 27856 39196
rect 27912 39194 27918 39196
rect 27672 39142 27674 39194
rect 27854 39142 27856 39194
rect 27610 39140 27616 39142
rect 27672 39140 27696 39142
rect 27752 39140 27776 39142
rect 27832 39140 27856 39142
rect 27912 39140 27918 39142
rect 27610 39131 27918 39140
rect 27610 38108 27918 38117
rect 27610 38106 27616 38108
rect 27672 38106 27696 38108
rect 27752 38106 27776 38108
rect 27832 38106 27856 38108
rect 27912 38106 27918 38108
rect 27672 38054 27674 38106
rect 27854 38054 27856 38106
rect 27610 38052 27616 38054
rect 27672 38052 27696 38054
rect 27752 38052 27776 38054
rect 27832 38052 27856 38054
rect 27912 38052 27918 38054
rect 27610 38043 27918 38052
rect 28000 37194 28028 41482
rect 27988 37188 28040 37194
rect 27988 37130 28040 37136
rect 27610 37020 27918 37029
rect 27610 37018 27616 37020
rect 27672 37018 27696 37020
rect 27752 37018 27776 37020
rect 27832 37018 27856 37020
rect 27912 37018 27918 37020
rect 27672 36966 27674 37018
rect 27854 36966 27856 37018
rect 27610 36964 27616 36966
rect 27672 36964 27696 36966
rect 27752 36964 27776 36966
rect 27832 36964 27856 36966
rect 27912 36964 27918 36966
rect 27610 36955 27918 36964
rect 27436 36916 27488 36922
rect 27436 36858 27488 36864
rect 27610 35932 27918 35941
rect 27610 35930 27616 35932
rect 27672 35930 27696 35932
rect 27752 35930 27776 35932
rect 27832 35930 27856 35932
rect 27912 35930 27918 35932
rect 27672 35878 27674 35930
rect 27854 35878 27856 35930
rect 27610 35876 27616 35878
rect 27672 35876 27696 35878
rect 27752 35876 27776 35878
rect 27832 35876 27856 35878
rect 27912 35876 27918 35878
rect 27610 35867 27918 35876
rect 27610 34844 27918 34853
rect 27610 34842 27616 34844
rect 27672 34842 27696 34844
rect 27752 34842 27776 34844
rect 27832 34842 27856 34844
rect 27912 34842 27918 34844
rect 27672 34790 27674 34842
rect 27854 34790 27856 34842
rect 27610 34788 27616 34790
rect 27672 34788 27696 34790
rect 27752 34788 27776 34790
rect 27832 34788 27856 34790
rect 27912 34788 27918 34790
rect 27610 34779 27918 34788
rect 27610 33756 27918 33765
rect 27610 33754 27616 33756
rect 27672 33754 27696 33756
rect 27752 33754 27776 33756
rect 27832 33754 27856 33756
rect 27912 33754 27918 33756
rect 27672 33702 27674 33754
rect 27854 33702 27856 33754
rect 27610 33700 27616 33702
rect 27672 33700 27696 33702
rect 27752 33700 27776 33702
rect 27832 33700 27856 33702
rect 27912 33700 27918 33702
rect 27610 33691 27918 33700
rect 27610 32668 27918 32677
rect 27610 32666 27616 32668
rect 27672 32666 27696 32668
rect 27752 32666 27776 32668
rect 27832 32666 27856 32668
rect 27912 32666 27918 32668
rect 27672 32614 27674 32666
rect 27854 32614 27856 32666
rect 27610 32612 27616 32614
rect 27672 32612 27696 32614
rect 27752 32612 27776 32614
rect 27832 32612 27856 32614
rect 27912 32612 27918 32614
rect 27610 32603 27918 32612
rect 28276 32502 28304 43726
rect 28264 32496 28316 32502
rect 28264 32438 28316 32444
rect 27610 31580 27918 31589
rect 27610 31578 27616 31580
rect 27672 31578 27696 31580
rect 27752 31578 27776 31580
rect 27832 31578 27856 31580
rect 27912 31578 27918 31580
rect 27672 31526 27674 31578
rect 27854 31526 27856 31578
rect 27610 31524 27616 31526
rect 27672 31524 27696 31526
rect 27752 31524 27776 31526
rect 27832 31524 27856 31526
rect 27912 31524 27918 31526
rect 27610 31515 27918 31524
rect 27610 30492 27918 30501
rect 27610 30490 27616 30492
rect 27672 30490 27696 30492
rect 27752 30490 27776 30492
rect 27832 30490 27856 30492
rect 27912 30490 27918 30492
rect 27672 30438 27674 30490
rect 27854 30438 27856 30490
rect 27610 30436 27616 30438
rect 27672 30436 27696 30438
rect 27752 30436 27776 30438
rect 27832 30436 27856 30438
rect 27912 30436 27918 30438
rect 27610 30427 27918 30436
rect 28644 30122 28672 55558
rect 28908 53644 28960 53650
rect 28908 53586 28960 53592
rect 28920 53038 28948 53586
rect 28908 53032 28960 53038
rect 28908 52974 28960 52980
rect 28816 52420 28868 52426
rect 28816 52362 28868 52368
rect 28828 51610 28856 52362
rect 28816 51604 28868 51610
rect 28816 51546 28868 51552
rect 28816 46572 28868 46578
rect 28816 46514 28868 46520
rect 28828 45937 28856 46514
rect 28920 46374 28948 52974
rect 28908 46368 28960 46374
rect 28908 46310 28960 46316
rect 28814 45928 28870 45937
rect 28920 45898 28948 46310
rect 28814 45863 28870 45872
rect 28908 45892 28960 45898
rect 28908 45834 28960 45840
rect 28920 41682 28948 45834
rect 28908 41676 28960 41682
rect 28908 41618 28960 41624
rect 28920 41546 28948 41618
rect 28908 41540 28960 41546
rect 28908 41482 28960 41488
rect 29012 41414 29040 56374
rect 29104 50862 29132 68342
rect 32404 68332 32456 68338
rect 32404 68274 32456 68280
rect 31852 68264 31904 68270
rect 31852 68206 31904 68212
rect 29920 67720 29972 67726
rect 29920 67662 29972 67668
rect 29644 60104 29696 60110
rect 29644 60046 29696 60052
rect 29656 56930 29684 60046
rect 29828 57860 29880 57866
rect 29828 57802 29880 57808
rect 29736 57792 29788 57798
rect 29736 57734 29788 57740
rect 29748 57390 29776 57734
rect 29840 57594 29868 57802
rect 29828 57588 29880 57594
rect 29828 57530 29880 57536
rect 29828 57452 29880 57458
rect 29828 57394 29880 57400
rect 29736 57384 29788 57390
rect 29736 57326 29788 57332
rect 29840 57050 29868 57394
rect 29828 57044 29880 57050
rect 29828 56986 29880 56992
rect 29656 56902 29868 56930
rect 29840 56778 29868 56902
rect 29828 56772 29880 56778
rect 29828 56714 29880 56720
rect 29184 56160 29236 56166
rect 29184 56102 29236 56108
rect 29092 50856 29144 50862
rect 29092 50798 29144 50804
rect 29104 49842 29132 50798
rect 29092 49836 29144 49842
rect 29092 49778 29144 49784
rect 29104 43722 29132 49778
rect 29092 43716 29144 43722
rect 29092 43658 29144 43664
rect 29012 41386 29132 41414
rect 29000 37800 29052 37806
rect 29000 37742 29052 37748
rect 29012 37466 29040 37742
rect 29000 37460 29052 37466
rect 29000 37402 29052 37408
rect 28908 32428 28960 32434
rect 28908 32370 28960 32376
rect 28724 31952 28776 31958
rect 28724 31894 28776 31900
rect 28632 30116 28684 30122
rect 28632 30058 28684 30064
rect 27610 29404 27918 29413
rect 27610 29402 27616 29404
rect 27672 29402 27696 29404
rect 27752 29402 27776 29404
rect 27832 29402 27856 29404
rect 27912 29402 27918 29404
rect 27672 29350 27674 29402
rect 27854 29350 27856 29402
rect 27610 29348 27616 29350
rect 27672 29348 27696 29350
rect 27752 29348 27776 29350
rect 27832 29348 27856 29350
rect 27912 29348 27918 29350
rect 27610 29339 27918 29348
rect 27610 28316 27918 28325
rect 27610 28314 27616 28316
rect 27672 28314 27696 28316
rect 27752 28314 27776 28316
rect 27832 28314 27856 28316
rect 27912 28314 27918 28316
rect 27672 28262 27674 28314
rect 27854 28262 27856 28314
rect 27610 28260 27616 28262
rect 27672 28260 27696 28262
rect 27752 28260 27776 28262
rect 27832 28260 27856 28262
rect 27912 28260 27918 28262
rect 27610 28251 27918 28260
rect 27610 27228 27918 27237
rect 27610 27226 27616 27228
rect 27672 27226 27696 27228
rect 27752 27226 27776 27228
rect 27832 27226 27856 27228
rect 27912 27226 27918 27228
rect 27672 27174 27674 27226
rect 27854 27174 27856 27226
rect 27610 27172 27616 27174
rect 27672 27172 27696 27174
rect 27752 27172 27776 27174
rect 27832 27172 27856 27174
rect 27912 27172 27918 27174
rect 27610 27163 27918 27172
rect 27610 26140 27918 26149
rect 27610 26138 27616 26140
rect 27672 26138 27696 26140
rect 27752 26138 27776 26140
rect 27832 26138 27856 26140
rect 27912 26138 27918 26140
rect 27672 26086 27674 26138
rect 27854 26086 27856 26138
rect 27610 26084 27616 26086
rect 27672 26084 27696 26086
rect 27752 26084 27776 26086
rect 27832 26084 27856 26086
rect 27912 26084 27918 26086
rect 27610 26075 27918 26084
rect 27610 25052 27918 25061
rect 27610 25050 27616 25052
rect 27672 25050 27696 25052
rect 27752 25050 27776 25052
rect 27832 25050 27856 25052
rect 27912 25050 27918 25052
rect 27672 24998 27674 25050
rect 27854 24998 27856 25050
rect 27610 24996 27616 24998
rect 27672 24996 27696 24998
rect 27752 24996 27776 24998
rect 27832 24996 27856 24998
rect 27912 24996 27918 24998
rect 27610 24987 27918 24996
rect 27344 24336 27396 24342
rect 27344 24278 27396 24284
rect 27610 23964 27918 23973
rect 27610 23962 27616 23964
rect 27672 23962 27696 23964
rect 27752 23962 27776 23964
rect 27832 23962 27856 23964
rect 27912 23962 27918 23964
rect 27672 23910 27674 23962
rect 27854 23910 27856 23962
rect 27610 23908 27616 23910
rect 27672 23908 27696 23910
rect 27752 23908 27776 23910
rect 27832 23908 27856 23910
rect 27912 23908 27918 23910
rect 27610 23899 27918 23908
rect 26950 23420 27258 23429
rect 26950 23418 26956 23420
rect 27012 23418 27036 23420
rect 27092 23418 27116 23420
rect 27172 23418 27196 23420
rect 27252 23418 27258 23420
rect 27012 23366 27014 23418
rect 27194 23366 27196 23418
rect 26950 23364 26956 23366
rect 27012 23364 27036 23366
rect 27092 23364 27116 23366
rect 27172 23364 27196 23366
rect 27252 23364 27258 23366
rect 26950 23355 27258 23364
rect 27610 22876 27918 22885
rect 27610 22874 27616 22876
rect 27672 22874 27696 22876
rect 27752 22874 27776 22876
rect 27832 22874 27856 22876
rect 27912 22874 27918 22876
rect 27672 22822 27674 22874
rect 27854 22822 27856 22874
rect 27610 22820 27616 22822
rect 27672 22820 27696 22822
rect 27752 22820 27776 22822
rect 27832 22820 27856 22822
rect 27912 22820 27918 22822
rect 27610 22811 27918 22820
rect 26950 22332 27258 22341
rect 26950 22330 26956 22332
rect 27012 22330 27036 22332
rect 27092 22330 27116 22332
rect 27172 22330 27196 22332
rect 27252 22330 27258 22332
rect 27012 22278 27014 22330
rect 27194 22278 27196 22330
rect 26950 22276 26956 22278
rect 27012 22276 27036 22278
rect 27092 22276 27116 22278
rect 27172 22276 27196 22278
rect 27252 22276 27258 22278
rect 26950 22267 27258 22276
rect 27610 21788 27918 21797
rect 27610 21786 27616 21788
rect 27672 21786 27696 21788
rect 27752 21786 27776 21788
rect 27832 21786 27856 21788
rect 27912 21786 27918 21788
rect 27672 21734 27674 21786
rect 27854 21734 27856 21786
rect 27610 21732 27616 21734
rect 27672 21732 27696 21734
rect 27752 21732 27776 21734
rect 27832 21732 27856 21734
rect 27912 21732 27918 21734
rect 27610 21723 27918 21732
rect 27528 21616 27580 21622
rect 27528 21558 27580 21564
rect 26950 21244 27258 21253
rect 26950 21242 26956 21244
rect 27012 21242 27036 21244
rect 27092 21242 27116 21244
rect 27172 21242 27196 21244
rect 27252 21242 27258 21244
rect 27012 21190 27014 21242
rect 27194 21190 27196 21242
rect 26950 21188 26956 21190
rect 27012 21188 27036 21190
rect 27092 21188 27116 21190
rect 27172 21188 27196 21190
rect 27252 21188 27258 21190
rect 26950 21179 27258 21188
rect 26950 20156 27258 20165
rect 26950 20154 26956 20156
rect 27012 20154 27036 20156
rect 27092 20154 27116 20156
rect 27172 20154 27196 20156
rect 27252 20154 27258 20156
rect 27012 20102 27014 20154
rect 27194 20102 27196 20154
rect 26950 20100 26956 20102
rect 27012 20100 27036 20102
rect 27092 20100 27116 20102
rect 27172 20100 27196 20102
rect 27252 20100 27258 20102
rect 26950 20091 27258 20100
rect 26950 19068 27258 19077
rect 26950 19066 26956 19068
rect 27012 19066 27036 19068
rect 27092 19066 27116 19068
rect 27172 19066 27196 19068
rect 27252 19066 27258 19068
rect 27012 19014 27014 19066
rect 27194 19014 27196 19066
rect 26950 19012 26956 19014
rect 27012 19012 27036 19014
rect 27092 19012 27116 19014
rect 27172 19012 27196 19014
rect 27252 19012 27258 19014
rect 26950 19003 27258 19012
rect 26804 18154 27016 18170
rect 26792 18148 27028 18154
rect 26844 18142 26976 18148
rect 26792 18090 26844 18096
rect 26976 18090 27028 18096
rect 26950 17980 27258 17989
rect 26950 17978 26956 17980
rect 27012 17978 27036 17980
rect 27092 17978 27116 17980
rect 27172 17978 27196 17980
rect 27252 17978 27258 17980
rect 27012 17926 27014 17978
rect 27194 17926 27196 17978
rect 26950 17924 26956 17926
rect 27012 17924 27036 17926
rect 27092 17924 27116 17926
rect 27172 17924 27196 17926
rect 27252 17924 27258 17926
rect 26950 17915 27258 17924
rect 26950 16892 27258 16901
rect 26950 16890 26956 16892
rect 27012 16890 27036 16892
rect 27092 16890 27116 16892
rect 27172 16890 27196 16892
rect 27252 16890 27258 16892
rect 27012 16838 27014 16890
rect 27194 16838 27196 16890
rect 26950 16836 26956 16838
rect 27012 16836 27036 16838
rect 27092 16836 27116 16838
rect 27172 16836 27196 16838
rect 27252 16836 27258 16838
rect 26950 16827 27258 16836
rect 26950 15804 27258 15813
rect 26950 15802 26956 15804
rect 27012 15802 27036 15804
rect 27092 15802 27116 15804
rect 27172 15802 27196 15804
rect 27252 15802 27258 15804
rect 27012 15750 27014 15802
rect 27194 15750 27196 15802
rect 26950 15748 26956 15750
rect 27012 15748 27036 15750
rect 27092 15748 27116 15750
rect 27172 15748 27196 15750
rect 27252 15748 27258 15750
rect 26950 15739 27258 15748
rect 26950 14716 27258 14725
rect 26950 14714 26956 14716
rect 27012 14714 27036 14716
rect 27092 14714 27116 14716
rect 27172 14714 27196 14716
rect 27252 14714 27258 14716
rect 27012 14662 27014 14714
rect 27194 14662 27196 14714
rect 26950 14660 26956 14662
rect 27012 14660 27036 14662
rect 27092 14660 27116 14662
rect 27172 14660 27196 14662
rect 27252 14660 27258 14662
rect 26950 14651 27258 14660
rect 26950 13628 27258 13637
rect 26950 13626 26956 13628
rect 27012 13626 27036 13628
rect 27092 13626 27116 13628
rect 27172 13626 27196 13628
rect 27252 13626 27258 13628
rect 27012 13574 27014 13626
rect 27194 13574 27196 13626
rect 26950 13572 26956 13574
rect 27012 13572 27036 13574
rect 27092 13572 27116 13574
rect 27172 13572 27196 13574
rect 27252 13572 27258 13574
rect 26950 13563 27258 13572
rect 27540 13530 27568 21558
rect 27610 20700 27918 20709
rect 27610 20698 27616 20700
rect 27672 20698 27696 20700
rect 27752 20698 27776 20700
rect 27832 20698 27856 20700
rect 27912 20698 27918 20700
rect 27672 20646 27674 20698
rect 27854 20646 27856 20698
rect 27610 20644 27616 20646
rect 27672 20644 27696 20646
rect 27752 20644 27776 20646
rect 27832 20644 27856 20646
rect 27912 20644 27918 20646
rect 27610 20635 27918 20644
rect 27610 19612 27918 19621
rect 27610 19610 27616 19612
rect 27672 19610 27696 19612
rect 27752 19610 27776 19612
rect 27832 19610 27856 19612
rect 27912 19610 27918 19612
rect 27672 19558 27674 19610
rect 27854 19558 27856 19610
rect 27610 19556 27616 19558
rect 27672 19556 27696 19558
rect 27752 19556 27776 19558
rect 27832 19556 27856 19558
rect 27912 19556 27918 19558
rect 27610 19547 27918 19556
rect 27610 18524 27918 18533
rect 27610 18522 27616 18524
rect 27672 18522 27696 18524
rect 27752 18522 27776 18524
rect 27832 18522 27856 18524
rect 27912 18522 27918 18524
rect 27672 18470 27674 18522
rect 27854 18470 27856 18522
rect 27610 18468 27616 18470
rect 27672 18468 27696 18470
rect 27752 18468 27776 18470
rect 27832 18468 27856 18470
rect 27912 18468 27918 18470
rect 27610 18459 27918 18468
rect 27610 17436 27918 17445
rect 27610 17434 27616 17436
rect 27672 17434 27696 17436
rect 27752 17434 27776 17436
rect 27832 17434 27856 17436
rect 27912 17434 27918 17436
rect 27672 17382 27674 17434
rect 27854 17382 27856 17434
rect 27610 17380 27616 17382
rect 27672 17380 27696 17382
rect 27752 17380 27776 17382
rect 27832 17380 27856 17382
rect 27912 17380 27918 17382
rect 27610 17371 27918 17380
rect 28736 17270 28764 31894
rect 28920 17270 28948 32370
rect 29000 30048 29052 30054
rect 29000 29990 29052 29996
rect 29012 27606 29040 29990
rect 29104 28218 29132 41386
rect 29092 28212 29144 28218
rect 29092 28154 29144 28160
rect 29092 28076 29144 28082
rect 29092 28018 29144 28024
rect 29104 27878 29132 28018
rect 29092 27872 29144 27878
rect 29092 27814 29144 27820
rect 29000 27600 29052 27606
rect 29000 27542 29052 27548
rect 29104 25226 29132 27814
rect 29092 25220 29144 25226
rect 29092 25162 29144 25168
rect 29000 25152 29052 25158
rect 29000 25094 29052 25100
rect 29012 21486 29040 25094
rect 29000 21480 29052 21486
rect 29000 21422 29052 21428
rect 29012 17270 29040 21422
rect 28724 17264 28776 17270
rect 28724 17206 28776 17212
rect 28908 17264 28960 17270
rect 28908 17206 28960 17212
rect 29000 17264 29052 17270
rect 29000 17206 29052 17212
rect 28540 16992 28592 16998
rect 28540 16934 28592 16940
rect 28552 16794 28580 16934
rect 28540 16788 28592 16794
rect 28540 16730 28592 16736
rect 27610 16348 27918 16357
rect 27610 16346 27616 16348
rect 27672 16346 27696 16348
rect 27752 16346 27776 16348
rect 27832 16346 27856 16348
rect 27912 16346 27918 16348
rect 27672 16294 27674 16346
rect 27854 16294 27856 16346
rect 27610 16292 27616 16294
rect 27672 16292 27696 16294
rect 27752 16292 27776 16294
rect 27832 16292 27856 16294
rect 27912 16292 27918 16294
rect 27610 16283 27918 16292
rect 27610 15260 27918 15269
rect 27610 15258 27616 15260
rect 27672 15258 27696 15260
rect 27752 15258 27776 15260
rect 27832 15258 27856 15260
rect 27912 15258 27918 15260
rect 27672 15206 27674 15258
rect 27854 15206 27856 15258
rect 27610 15204 27616 15206
rect 27672 15204 27696 15206
rect 27752 15204 27776 15206
rect 27832 15204 27856 15206
rect 27912 15204 27918 15206
rect 27610 15195 27918 15204
rect 27610 14172 27918 14181
rect 27610 14170 27616 14172
rect 27672 14170 27696 14172
rect 27752 14170 27776 14172
rect 27832 14170 27856 14172
rect 27912 14170 27918 14172
rect 27672 14118 27674 14170
rect 27854 14118 27856 14170
rect 27610 14116 27616 14118
rect 27672 14116 27696 14118
rect 27752 14116 27776 14118
rect 27832 14116 27856 14118
rect 27912 14116 27918 14118
rect 27610 14107 27918 14116
rect 27528 13524 27580 13530
rect 27528 13466 27580 13472
rect 27610 13084 27918 13093
rect 27610 13082 27616 13084
rect 27672 13082 27696 13084
rect 27752 13082 27776 13084
rect 27832 13082 27856 13084
rect 27912 13082 27918 13084
rect 27672 13030 27674 13082
rect 27854 13030 27856 13082
rect 27610 13028 27616 13030
rect 27672 13028 27696 13030
rect 27752 13028 27776 13030
rect 27832 13028 27856 13030
rect 27912 13028 27918 13030
rect 27610 13019 27918 13028
rect 26950 12540 27258 12549
rect 26950 12538 26956 12540
rect 27012 12538 27036 12540
rect 27092 12538 27116 12540
rect 27172 12538 27196 12540
rect 27252 12538 27258 12540
rect 27012 12486 27014 12538
rect 27194 12486 27196 12538
rect 26950 12484 26956 12486
rect 27012 12484 27036 12486
rect 27092 12484 27116 12486
rect 27172 12484 27196 12486
rect 27252 12484 27258 12486
rect 26950 12475 27258 12484
rect 27610 11996 27918 12005
rect 27610 11994 27616 11996
rect 27672 11994 27696 11996
rect 27752 11994 27776 11996
rect 27832 11994 27856 11996
rect 27912 11994 27918 11996
rect 27672 11942 27674 11994
rect 27854 11942 27856 11994
rect 27610 11940 27616 11942
rect 27672 11940 27696 11942
rect 27752 11940 27776 11942
rect 27832 11940 27856 11942
rect 27912 11940 27918 11942
rect 27610 11931 27918 11940
rect 26950 11452 27258 11461
rect 26950 11450 26956 11452
rect 27012 11450 27036 11452
rect 27092 11450 27116 11452
rect 27172 11450 27196 11452
rect 27252 11450 27258 11452
rect 27012 11398 27014 11450
rect 27194 11398 27196 11450
rect 26950 11396 26956 11398
rect 27012 11396 27036 11398
rect 27092 11396 27116 11398
rect 27172 11396 27196 11398
rect 27252 11396 27258 11398
rect 26950 11387 27258 11396
rect 27610 10908 27918 10917
rect 27610 10906 27616 10908
rect 27672 10906 27696 10908
rect 27752 10906 27776 10908
rect 27832 10906 27856 10908
rect 27912 10906 27918 10908
rect 27672 10854 27674 10906
rect 27854 10854 27856 10906
rect 27610 10852 27616 10854
rect 27672 10852 27696 10854
rect 27752 10852 27776 10854
rect 27832 10852 27856 10854
rect 27912 10852 27918 10854
rect 27610 10843 27918 10852
rect 26950 10364 27258 10373
rect 26950 10362 26956 10364
rect 27012 10362 27036 10364
rect 27092 10362 27116 10364
rect 27172 10362 27196 10364
rect 27252 10362 27258 10364
rect 27012 10310 27014 10362
rect 27194 10310 27196 10362
rect 26950 10308 26956 10310
rect 27012 10308 27036 10310
rect 27092 10308 27116 10310
rect 27172 10308 27196 10310
rect 27252 10308 27258 10310
rect 26950 10299 27258 10308
rect 27610 9820 27918 9829
rect 27610 9818 27616 9820
rect 27672 9818 27696 9820
rect 27752 9818 27776 9820
rect 27832 9818 27856 9820
rect 27912 9818 27918 9820
rect 27672 9766 27674 9818
rect 27854 9766 27856 9818
rect 27610 9764 27616 9766
rect 27672 9764 27696 9766
rect 27752 9764 27776 9766
rect 27832 9764 27856 9766
rect 27912 9764 27918 9766
rect 27610 9755 27918 9764
rect 26950 9276 27258 9285
rect 26950 9274 26956 9276
rect 27012 9274 27036 9276
rect 27092 9274 27116 9276
rect 27172 9274 27196 9276
rect 27252 9274 27258 9276
rect 27012 9222 27014 9274
rect 27194 9222 27196 9274
rect 26950 9220 26956 9222
rect 27012 9220 27036 9222
rect 27092 9220 27116 9222
rect 27172 9220 27196 9222
rect 27252 9220 27258 9222
rect 26950 9211 27258 9220
rect 27610 8732 27918 8741
rect 27610 8730 27616 8732
rect 27672 8730 27696 8732
rect 27752 8730 27776 8732
rect 27832 8730 27856 8732
rect 27912 8730 27918 8732
rect 27672 8678 27674 8730
rect 27854 8678 27856 8730
rect 27610 8676 27616 8678
rect 27672 8676 27696 8678
rect 27752 8676 27776 8678
rect 27832 8676 27856 8678
rect 27912 8676 27918 8678
rect 27610 8667 27918 8676
rect 26950 8188 27258 8197
rect 26950 8186 26956 8188
rect 27012 8186 27036 8188
rect 27092 8186 27116 8188
rect 27172 8186 27196 8188
rect 27252 8186 27258 8188
rect 27012 8134 27014 8186
rect 27194 8134 27196 8186
rect 26950 8132 26956 8134
rect 27012 8132 27036 8134
rect 27092 8132 27116 8134
rect 27172 8132 27196 8134
rect 27252 8132 27258 8134
rect 26950 8123 27258 8132
rect 27610 7644 27918 7653
rect 27610 7642 27616 7644
rect 27672 7642 27696 7644
rect 27752 7642 27776 7644
rect 27832 7642 27856 7644
rect 27912 7642 27918 7644
rect 27672 7590 27674 7642
rect 27854 7590 27856 7642
rect 27610 7588 27616 7590
rect 27672 7588 27696 7590
rect 27752 7588 27776 7590
rect 27832 7588 27856 7590
rect 27912 7588 27918 7590
rect 27610 7579 27918 7588
rect 26950 7100 27258 7109
rect 26950 7098 26956 7100
rect 27012 7098 27036 7100
rect 27092 7098 27116 7100
rect 27172 7098 27196 7100
rect 27252 7098 27258 7100
rect 27012 7046 27014 7098
rect 27194 7046 27196 7098
rect 26950 7044 26956 7046
rect 27012 7044 27036 7046
rect 27092 7044 27116 7046
rect 27172 7044 27196 7046
rect 27252 7044 27258 7046
rect 26950 7035 27258 7044
rect 27610 6556 27918 6565
rect 27610 6554 27616 6556
rect 27672 6554 27696 6556
rect 27752 6554 27776 6556
rect 27832 6554 27856 6556
rect 27912 6554 27918 6556
rect 27672 6502 27674 6554
rect 27854 6502 27856 6554
rect 27610 6500 27616 6502
rect 27672 6500 27696 6502
rect 27752 6500 27776 6502
rect 27832 6500 27856 6502
rect 27912 6500 27918 6502
rect 27610 6491 27918 6500
rect 26950 6012 27258 6021
rect 26950 6010 26956 6012
rect 27012 6010 27036 6012
rect 27092 6010 27116 6012
rect 27172 6010 27196 6012
rect 27252 6010 27258 6012
rect 27012 5958 27014 6010
rect 27194 5958 27196 6010
rect 26950 5956 26956 5958
rect 27012 5956 27036 5958
rect 27092 5956 27116 5958
rect 27172 5956 27196 5958
rect 27252 5956 27258 5958
rect 26950 5947 27258 5956
rect 27610 5468 27918 5477
rect 27610 5466 27616 5468
rect 27672 5466 27696 5468
rect 27752 5466 27776 5468
rect 27832 5466 27856 5468
rect 27912 5466 27918 5468
rect 27672 5414 27674 5466
rect 27854 5414 27856 5466
rect 27610 5412 27616 5414
rect 27672 5412 27696 5414
rect 27752 5412 27776 5414
rect 27832 5412 27856 5414
rect 27912 5412 27918 5414
rect 27610 5403 27918 5412
rect 26950 4924 27258 4933
rect 26950 4922 26956 4924
rect 27012 4922 27036 4924
rect 27092 4922 27116 4924
rect 27172 4922 27196 4924
rect 27252 4922 27258 4924
rect 27012 4870 27014 4922
rect 27194 4870 27196 4922
rect 26950 4868 26956 4870
rect 27012 4868 27036 4870
rect 27092 4868 27116 4870
rect 27172 4868 27196 4870
rect 27252 4868 27258 4870
rect 26950 4859 27258 4868
rect 26056 4820 26108 4826
rect 26056 4762 26108 4768
rect 28920 4758 28948 17206
rect 29104 17202 29132 25162
rect 29092 17196 29144 17202
rect 29092 17138 29144 17144
rect 28908 4752 28960 4758
rect 28908 4694 28960 4700
rect 25780 4616 25832 4622
rect 25780 4558 25832 4564
rect 23756 4548 23808 4554
rect 23756 4490 23808 4496
rect 22610 4380 22918 4389
rect 22610 4378 22616 4380
rect 22672 4378 22696 4380
rect 22752 4378 22776 4380
rect 22832 4378 22856 4380
rect 22912 4378 22918 4380
rect 22672 4326 22674 4378
rect 22854 4326 22856 4378
rect 22610 4324 22616 4326
rect 22672 4324 22696 4326
rect 22752 4324 22776 4326
rect 22832 4324 22856 4326
rect 22912 4324 22918 4326
rect 22610 4315 22918 4324
rect 27610 4380 27918 4389
rect 27610 4378 27616 4380
rect 27672 4378 27696 4380
rect 27752 4378 27776 4380
rect 27832 4378 27856 4380
rect 27912 4378 27918 4380
rect 27672 4326 27674 4378
rect 27854 4326 27856 4378
rect 27610 4324 27616 4326
rect 27672 4324 27696 4326
rect 27752 4324 27776 4326
rect 27832 4324 27856 4326
rect 27912 4324 27918 4326
rect 27610 4315 27918 4324
rect 21950 3836 22258 3845
rect 21950 3834 21956 3836
rect 22012 3834 22036 3836
rect 22092 3834 22116 3836
rect 22172 3834 22196 3836
rect 22252 3834 22258 3836
rect 22012 3782 22014 3834
rect 22194 3782 22196 3834
rect 21950 3780 21956 3782
rect 22012 3780 22036 3782
rect 22092 3780 22116 3782
rect 22172 3780 22196 3782
rect 22252 3780 22258 3782
rect 21950 3771 22258 3780
rect 26950 3836 27258 3845
rect 26950 3834 26956 3836
rect 27012 3834 27036 3836
rect 27092 3834 27116 3836
rect 27172 3834 27196 3836
rect 27252 3834 27258 3836
rect 27012 3782 27014 3834
rect 27194 3782 27196 3834
rect 26950 3780 26956 3782
rect 27012 3780 27036 3782
rect 27092 3780 27116 3782
rect 27172 3780 27196 3782
rect 27252 3780 27258 3782
rect 26950 3771 27258 3780
rect 22610 3292 22918 3301
rect 22610 3290 22616 3292
rect 22672 3290 22696 3292
rect 22752 3290 22776 3292
rect 22832 3290 22856 3292
rect 22912 3290 22918 3292
rect 22672 3238 22674 3290
rect 22854 3238 22856 3290
rect 22610 3236 22616 3238
rect 22672 3236 22696 3238
rect 22752 3236 22776 3238
rect 22832 3236 22856 3238
rect 22912 3236 22918 3238
rect 22610 3227 22918 3236
rect 27610 3292 27918 3301
rect 27610 3290 27616 3292
rect 27672 3290 27696 3292
rect 27752 3290 27776 3292
rect 27832 3290 27856 3292
rect 27912 3290 27918 3292
rect 27672 3238 27674 3290
rect 27854 3238 27856 3290
rect 27610 3236 27616 3238
rect 27672 3236 27696 3238
rect 27752 3236 27776 3238
rect 27832 3236 27856 3238
rect 27912 3236 27918 3238
rect 27610 3227 27918 3236
rect 29196 3058 29224 56102
rect 29644 55616 29696 55622
rect 29644 55558 29696 55564
rect 29552 50516 29604 50522
rect 29552 50458 29604 50464
rect 29368 49972 29420 49978
rect 29368 49914 29420 49920
rect 29276 43716 29328 43722
rect 29276 43658 29328 43664
rect 29288 30054 29316 43658
rect 29276 30048 29328 30054
rect 29276 29990 29328 29996
rect 29276 28144 29328 28150
rect 29276 28086 29328 28092
rect 29288 25158 29316 28086
rect 29380 25294 29408 49914
rect 29460 31748 29512 31754
rect 29460 31690 29512 31696
rect 29472 31142 29500 31690
rect 29460 31136 29512 31142
rect 29460 31078 29512 31084
rect 29460 28620 29512 28626
rect 29460 28562 29512 28568
rect 29368 25288 29420 25294
rect 29368 25230 29420 25236
rect 29276 25152 29328 25158
rect 29276 25094 29328 25100
rect 29472 3738 29500 28562
rect 29564 28218 29592 50458
rect 29552 28212 29604 28218
rect 29552 28154 29604 28160
rect 29656 11286 29684 55558
rect 29840 51074 29868 56714
rect 29932 55350 29960 67662
rect 31668 57520 31720 57526
rect 31668 57462 31720 57468
rect 30564 56704 30616 56710
rect 30564 56646 30616 56652
rect 29920 55344 29972 55350
rect 29920 55286 29972 55292
rect 30576 55282 30604 56646
rect 30564 55276 30616 55282
rect 30564 55218 30616 55224
rect 29748 51046 29868 51074
rect 29748 48074 29776 51046
rect 30380 48136 30432 48142
rect 30380 48078 30432 48084
rect 29736 48068 29788 48074
rect 29736 48010 29788 48016
rect 29748 45966 29776 48010
rect 30392 47666 30420 48078
rect 30380 47660 30432 47666
rect 30380 47602 30432 47608
rect 30392 47054 30420 47602
rect 30380 47048 30432 47054
rect 30380 46990 30432 46996
rect 30472 47048 30524 47054
rect 30472 46990 30524 46996
rect 29736 45960 29788 45966
rect 29736 45902 29788 45908
rect 29748 39438 29776 45902
rect 30484 41682 30512 46990
rect 30576 44878 30604 55218
rect 31576 53508 31628 53514
rect 31576 53450 31628 53456
rect 31588 53242 31616 53450
rect 31576 53236 31628 53242
rect 31576 53178 31628 53184
rect 31300 51808 31352 51814
rect 31300 51750 31352 51756
rect 30564 44872 30616 44878
rect 30564 44814 30616 44820
rect 30472 41676 30524 41682
rect 30472 41618 30524 41624
rect 30576 41414 30604 44814
rect 30748 41744 30800 41750
rect 30748 41686 30800 41692
rect 30760 41478 30788 41686
rect 30748 41472 30800 41478
rect 30748 41414 30800 41420
rect 30576 41386 30696 41414
rect 29736 39432 29788 39438
rect 29736 39374 29788 39380
rect 29748 13938 29776 39374
rect 30668 36310 30696 41386
rect 31312 40662 31340 51750
rect 31300 40656 31352 40662
rect 31300 40598 31352 40604
rect 30840 39296 30892 39302
rect 30840 39238 30892 39244
rect 30656 36304 30708 36310
rect 30656 36246 30708 36252
rect 29828 35216 29880 35222
rect 29828 35158 29880 35164
rect 29840 31822 29868 35158
rect 29828 31816 29880 31822
rect 29828 31758 29880 31764
rect 30562 28792 30618 28801
rect 30562 28727 30618 28736
rect 30576 28694 30604 28727
rect 30564 28688 30616 28694
rect 30564 28630 30616 28636
rect 30852 19446 30880 39238
rect 31576 37936 31628 37942
rect 31576 37878 31628 37884
rect 31484 36712 31536 36718
rect 31484 36654 31536 36660
rect 31496 36530 31524 36654
rect 31588 36650 31616 37878
rect 31576 36644 31628 36650
rect 31576 36586 31628 36592
rect 31496 36502 31616 36530
rect 31484 32768 31536 32774
rect 31484 32710 31536 32716
rect 31496 32434 31524 32710
rect 31484 32428 31536 32434
rect 31484 32370 31536 32376
rect 31588 31482 31616 36502
rect 31680 33266 31708 57462
rect 31760 49088 31812 49094
rect 31760 49030 31812 49036
rect 31772 33522 31800 49030
rect 31864 37942 31892 68206
rect 31950 68028 32258 68037
rect 31950 68026 31956 68028
rect 32012 68026 32036 68028
rect 32092 68026 32116 68028
rect 32172 68026 32196 68028
rect 32252 68026 32258 68028
rect 32012 67974 32014 68026
rect 32194 67974 32196 68026
rect 31950 67972 31956 67974
rect 32012 67972 32036 67974
rect 32092 67972 32116 67974
rect 32172 67972 32196 67974
rect 32252 67972 32258 67974
rect 31950 67963 32258 67972
rect 32416 67697 32444 68274
rect 32402 67688 32458 67697
rect 32402 67623 32458 67632
rect 32610 67484 32918 67493
rect 32610 67482 32616 67484
rect 32672 67482 32696 67484
rect 32752 67482 32776 67484
rect 32832 67482 32856 67484
rect 32912 67482 32918 67484
rect 32672 67430 32674 67482
rect 32854 67430 32856 67482
rect 32610 67428 32616 67430
rect 32672 67428 32696 67430
rect 32752 67428 32776 67430
rect 32832 67428 32856 67430
rect 32912 67428 32918 67430
rect 32610 67419 32918 67428
rect 31950 66940 32258 66949
rect 31950 66938 31956 66940
rect 32012 66938 32036 66940
rect 32092 66938 32116 66940
rect 32172 66938 32196 66940
rect 32252 66938 32258 66940
rect 32012 66886 32014 66938
rect 32194 66886 32196 66938
rect 31950 66884 31956 66886
rect 32012 66884 32036 66886
rect 32092 66884 32116 66886
rect 32172 66884 32196 66886
rect 32252 66884 32258 66886
rect 31950 66875 32258 66884
rect 32610 66396 32918 66405
rect 32610 66394 32616 66396
rect 32672 66394 32696 66396
rect 32752 66394 32776 66396
rect 32832 66394 32856 66396
rect 32912 66394 32918 66396
rect 32672 66342 32674 66394
rect 32854 66342 32856 66394
rect 32610 66340 32616 66342
rect 32672 66340 32696 66342
rect 32752 66340 32776 66342
rect 32832 66340 32856 66342
rect 32912 66340 32918 66342
rect 32610 66331 32918 66340
rect 31950 65852 32258 65861
rect 31950 65850 31956 65852
rect 32012 65850 32036 65852
rect 32092 65850 32116 65852
rect 32172 65850 32196 65852
rect 32252 65850 32258 65852
rect 32012 65798 32014 65850
rect 32194 65798 32196 65850
rect 31950 65796 31956 65798
rect 32012 65796 32036 65798
rect 32092 65796 32116 65798
rect 32172 65796 32196 65798
rect 32252 65796 32258 65798
rect 31950 65787 32258 65796
rect 32610 65308 32918 65317
rect 32610 65306 32616 65308
rect 32672 65306 32696 65308
rect 32752 65306 32776 65308
rect 32832 65306 32856 65308
rect 32912 65306 32918 65308
rect 32672 65254 32674 65306
rect 32854 65254 32856 65306
rect 32610 65252 32616 65254
rect 32672 65252 32696 65254
rect 32752 65252 32776 65254
rect 32832 65252 32856 65254
rect 32912 65252 32918 65254
rect 32610 65243 32918 65252
rect 31950 64764 32258 64773
rect 31950 64762 31956 64764
rect 32012 64762 32036 64764
rect 32092 64762 32116 64764
rect 32172 64762 32196 64764
rect 32252 64762 32258 64764
rect 32012 64710 32014 64762
rect 32194 64710 32196 64762
rect 31950 64708 31956 64710
rect 32012 64708 32036 64710
rect 32092 64708 32116 64710
rect 32172 64708 32196 64710
rect 32252 64708 32258 64710
rect 31950 64699 32258 64708
rect 32610 64220 32918 64229
rect 32610 64218 32616 64220
rect 32672 64218 32696 64220
rect 32752 64218 32776 64220
rect 32832 64218 32856 64220
rect 32912 64218 32918 64220
rect 32672 64166 32674 64218
rect 32854 64166 32856 64218
rect 32610 64164 32616 64166
rect 32672 64164 32696 64166
rect 32752 64164 32776 64166
rect 32832 64164 32856 64166
rect 32912 64164 32918 64166
rect 32610 64155 32918 64164
rect 32496 63776 32548 63782
rect 32496 63718 32548 63724
rect 31950 63676 32258 63685
rect 31950 63674 31956 63676
rect 32012 63674 32036 63676
rect 32092 63674 32116 63676
rect 32172 63674 32196 63676
rect 32252 63674 32258 63676
rect 32012 63622 32014 63674
rect 32194 63622 32196 63674
rect 31950 63620 31956 63622
rect 32012 63620 32036 63622
rect 32092 63620 32116 63622
rect 32172 63620 32196 63622
rect 32252 63620 32258 63622
rect 31950 63611 32258 63620
rect 31950 62588 32258 62597
rect 31950 62586 31956 62588
rect 32012 62586 32036 62588
rect 32092 62586 32116 62588
rect 32172 62586 32196 62588
rect 32252 62586 32258 62588
rect 32012 62534 32014 62586
rect 32194 62534 32196 62586
rect 31950 62532 31956 62534
rect 32012 62532 32036 62534
rect 32092 62532 32116 62534
rect 32172 62532 32196 62534
rect 32252 62532 32258 62534
rect 31950 62523 32258 62532
rect 31950 61500 32258 61509
rect 31950 61498 31956 61500
rect 32012 61498 32036 61500
rect 32092 61498 32116 61500
rect 32172 61498 32196 61500
rect 32252 61498 32258 61500
rect 32012 61446 32014 61498
rect 32194 61446 32196 61498
rect 31950 61444 31956 61446
rect 32012 61444 32036 61446
rect 32092 61444 32116 61446
rect 32172 61444 32196 61446
rect 32252 61444 32258 61446
rect 31950 61435 32258 61444
rect 31950 60412 32258 60421
rect 31950 60410 31956 60412
rect 32012 60410 32036 60412
rect 32092 60410 32116 60412
rect 32172 60410 32196 60412
rect 32252 60410 32258 60412
rect 32012 60358 32014 60410
rect 32194 60358 32196 60410
rect 31950 60356 31956 60358
rect 32012 60356 32036 60358
rect 32092 60356 32116 60358
rect 32172 60356 32196 60358
rect 32252 60356 32258 60358
rect 31950 60347 32258 60356
rect 31950 59324 32258 59333
rect 31950 59322 31956 59324
rect 32012 59322 32036 59324
rect 32092 59322 32116 59324
rect 32172 59322 32196 59324
rect 32252 59322 32258 59324
rect 32012 59270 32014 59322
rect 32194 59270 32196 59322
rect 31950 59268 31956 59270
rect 32012 59268 32036 59270
rect 32092 59268 32116 59270
rect 32172 59268 32196 59270
rect 32252 59268 32258 59270
rect 31950 59259 32258 59268
rect 31950 58236 32258 58245
rect 31950 58234 31956 58236
rect 32012 58234 32036 58236
rect 32092 58234 32116 58236
rect 32172 58234 32196 58236
rect 32252 58234 32258 58236
rect 32012 58182 32014 58234
rect 32194 58182 32196 58234
rect 31950 58180 31956 58182
rect 32012 58180 32036 58182
rect 32092 58180 32116 58182
rect 32172 58180 32196 58182
rect 32252 58180 32258 58182
rect 31950 58171 32258 58180
rect 31950 57148 32258 57157
rect 31950 57146 31956 57148
rect 32012 57146 32036 57148
rect 32092 57146 32116 57148
rect 32172 57146 32196 57148
rect 32252 57146 32258 57148
rect 32012 57094 32014 57146
rect 32194 57094 32196 57146
rect 31950 57092 31956 57094
rect 32012 57092 32036 57094
rect 32092 57092 32116 57094
rect 32172 57092 32196 57094
rect 32252 57092 32258 57094
rect 31950 57083 32258 57092
rect 31950 56060 32258 56069
rect 31950 56058 31956 56060
rect 32012 56058 32036 56060
rect 32092 56058 32116 56060
rect 32172 56058 32196 56060
rect 32252 56058 32258 56060
rect 32012 56006 32014 56058
rect 32194 56006 32196 56058
rect 31950 56004 31956 56006
rect 32012 56004 32036 56006
rect 32092 56004 32116 56006
rect 32172 56004 32196 56006
rect 32252 56004 32258 56006
rect 31950 55995 32258 56004
rect 31950 54972 32258 54981
rect 31950 54970 31956 54972
rect 32012 54970 32036 54972
rect 32092 54970 32116 54972
rect 32172 54970 32196 54972
rect 32252 54970 32258 54972
rect 32012 54918 32014 54970
rect 32194 54918 32196 54970
rect 31950 54916 31956 54918
rect 32012 54916 32036 54918
rect 32092 54916 32116 54918
rect 32172 54916 32196 54918
rect 32252 54916 32258 54918
rect 31950 54907 32258 54916
rect 31950 53884 32258 53893
rect 31950 53882 31956 53884
rect 32012 53882 32036 53884
rect 32092 53882 32116 53884
rect 32172 53882 32196 53884
rect 32252 53882 32258 53884
rect 32012 53830 32014 53882
rect 32194 53830 32196 53882
rect 31950 53828 31956 53830
rect 32012 53828 32036 53830
rect 32092 53828 32116 53830
rect 32172 53828 32196 53830
rect 32252 53828 32258 53830
rect 31950 53819 32258 53828
rect 31950 52796 32258 52805
rect 31950 52794 31956 52796
rect 32012 52794 32036 52796
rect 32092 52794 32116 52796
rect 32172 52794 32196 52796
rect 32252 52794 32258 52796
rect 32012 52742 32014 52794
rect 32194 52742 32196 52794
rect 31950 52740 31956 52742
rect 32012 52740 32036 52742
rect 32092 52740 32116 52742
rect 32172 52740 32196 52742
rect 32252 52740 32258 52742
rect 31950 52731 32258 52740
rect 32312 52012 32364 52018
rect 32312 51954 32364 51960
rect 31950 51708 32258 51717
rect 31950 51706 31956 51708
rect 32012 51706 32036 51708
rect 32092 51706 32116 51708
rect 32172 51706 32196 51708
rect 32252 51706 32258 51708
rect 32012 51654 32014 51706
rect 32194 51654 32196 51706
rect 31950 51652 31956 51654
rect 32012 51652 32036 51654
rect 32092 51652 32116 51654
rect 32172 51652 32196 51654
rect 32252 51652 32258 51654
rect 31950 51643 32258 51652
rect 31950 50620 32258 50629
rect 31950 50618 31956 50620
rect 32012 50618 32036 50620
rect 32092 50618 32116 50620
rect 32172 50618 32196 50620
rect 32252 50618 32258 50620
rect 32012 50566 32014 50618
rect 32194 50566 32196 50618
rect 31950 50564 31956 50566
rect 32012 50564 32036 50566
rect 32092 50564 32116 50566
rect 32172 50564 32196 50566
rect 32252 50564 32258 50566
rect 31950 50555 32258 50564
rect 31950 49532 32258 49541
rect 31950 49530 31956 49532
rect 32012 49530 32036 49532
rect 32092 49530 32116 49532
rect 32172 49530 32196 49532
rect 32252 49530 32258 49532
rect 32012 49478 32014 49530
rect 32194 49478 32196 49530
rect 31950 49476 31956 49478
rect 32012 49476 32036 49478
rect 32092 49476 32116 49478
rect 32172 49476 32196 49478
rect 32252 49476 32258 49478
rect 31950 49467 32258 49476
rect 31950 48444 32258 48453
rect 31950 48442 31956 48444
rect 32012 48442 32036 48444
rect 32092 48442 32116 48444
rect 32172 48442 32196 48444
rect 32252 48442 32258 48444
rect 32012 48390 32014 48442
rect 32194 48390 32196 48442
rect 31950 48388 31956 48390
rect 32012 48388 32036 48390
rect 32092 48388 32116 48390
rect 32172 48388 32196 48390
rect 32252 48388 32258 48390
rect 31950 48379 32258 48388
rect 31950 47356 32258 47365
rect 31950 47354 31956 47356
rect 32012 47354 32036 47356
rect 32092 47354 32116 47356
rect 32172 47354 32196 47356
rect 32252 47354 32258 47356
rect 32012 47302 32014 47354
rect 32194 47302 32196 47354
rect 31950 47300 31956 47302
rect 32012 47300 32036 47302
rect 32092 47300 32116 47302
rect 32172 47300 32196 47302
rect 32252 47300 32258 47302
rect 31950 47291 32258 47300
rect 31950 46268 32258 46277
rect 31950 46266 31956 46268
rect 32012 46266 32036 46268
rect 32092 46266 32116 46268
rect 32172 46266 32196 46268
rect 32252 46266 32258 46268
rect 32012 46214 32014 46266
rect 32194 46214 32196 46266
rect 31950 46212 31956 46214
rect 32012 46212 32036 46214
rect 32092 46212 32116 46214
rect 32172 46212 32196 46214
rect 32252 46212 32258 46214
rect 31950 46203 32258 46212
rect 31950 45180 32258 45189
rect 31950 45178 31956 45180
rect 32012 45178 32036 45180
rect 32092 45178 32116 45180
rect 32172 45178 32196 45180
rect 32252 45178 32258 45180
rect 32012 45126 32014 45178
rect 32194 45126 32196 45178
rect 31950 45124 31956 45126
rect 32012 45124 32036 45126
rect 32092 45124 32116 45126
rect 32172 45124 32196 45126
rect 32252 45124 32258 45126
rect 31950 45115 32258 45124
rect 31950 44092 32258 44101
rect 31950 44090 31956 44092
rect 32012 44090 32036 44092
rect 32092 44090 32116 44092
rect 32172 44090 32196 44092
rect 32252 44090 32258 44092
rect 32012 44038 32014 44090
rect 32194 44038 32196 44090
rect 31950 44036 31956 44038
rect 32012 44036 32036 44038
rect 32092 44036 32116 44038
rect 32172 44036 32196 44038
rect 32252 44036 32258 44038
rect 31950 44027 32258 44036
rect 31950 43004 32258 43013
rect 31950 43002 31956 43004
rect 32012 43002 32036 43004
rect 32092 43002 32116 43004
rect 32172 43002 32196 43004
rect 32252 43002 32258 43004
rect 32012 42950 32014 43002
rect 32194 42950 32196 43002
rect 31950 42948 31956 42950
rect 32012 42948 32036 42950
rect 32092 42948 32116 42950
rect 32172 42948 32196 42950
rect 32252 42948 32258 42950
rect 31950 42939 32258 42948
rect 31950 41916 32258 41925
rect 31950 41914 31956 41916
rect 32012 41914 32036 41916
rect 32092 41914 32116 41916
rect 32172 41914 32196 41916
rect 32252 41914 32258 41916
rect 32012 41862 32014 41914
rect 32194 41862 32196 41914
rect 31950 41860 31956 41862
rect 32012 41860 32036 41862
rect 32092 41860 32116 41862
rect 32172 41860 32196 41862
rect 32252 41860 32258 41862
rect 31950 41851 32258 41860
rect 31950 40828 32258 40837
rect 31950 40826 31956 40828
rect 32012 40826 32036 40828
rect 32092 40826 32116 40828
rect 32172 40826 32196 40828
rect 32252 40826 32258 40828
rect 32012 40774 32014 40826
rect 32194 40774 32196 40826
rect 31950 40772 31956 40774
rect 32012 40772 32036 40774
rect 32092 40772 32116 40774
rect 32172 40772 32196 40774
rect 32252 40772 32258 40774
rect 31950 40763 32258 40772
rect 31950 39740 32258 39749
rect 31950 39738 31956 39740
rect 32012 39738 32036 39740
rect 32092 39738 32116 39740
rect 32172 39738 32196 39740
rect 32252 39738 32258 39740
rect 32012 39686 32014 39738
rect 32194 39686 32196 39738
rect 31950 39684 31956 39686
rect 32012 39684 32036 39686
rect 32092 39684 32116 39686
rect 32172 39684 32196 39686
rect 32252 39684 32258 39686
rect 31950 39675 32258 39684
rect 31950 38652 32258 38661
rect 31950 38650 31956 38652
rect 32012 38650 32036 38652
rect 32092 38650 32116 38652
rect 32172 38650 32196 38652
rect 32252 38650 32258 38652
rect 32012 38598 32014 38650
rect 32194 38598 32196 38650
rect 31950 38596 31956 38598
rect 32012 38596 32036 38598
rect 32092 38596 32116 38598
rect 32172 38596 32196 38598
rect 32252 38596 32258 38598
rect 31950 38587 32258 38596
rect 31852 37936 31904 37942
rect 31852 37878 31904 37884
rect 31852 37800 31904 37806
rect 31852 37742 31904 37748
rect 31864 36174 31892 37742
rect 31950 37564 32258 37573
rect 31950 37562 31956 37564
rect 32012 37562 32036 37564
rect 32092 37562 32116 37564
rect 32172 37562 32196 37564
rect 32252 37562 32258 37564
rect 32012 37510 32014 37562
rect 32194 37510 32196 37562
rect 31950 37508 31956 37510
rect 32012 37508 32036 37510
rect 32092 37508 32116 37510
rect 32172 37508 32196 37510
rect 32252 37508 32258 37510
rect 31950 37499 32258 37508
rect 31950 36476 32258 36485
rect 31950 36474 31956 36476
rect 32012 36474 32036 36476
rect 32092 36474 32116 36476
rect 32172 36474 32196 36476
rect 32252 36474 32258 36476
rect 32012 36422 32014 36474
rect 32194 36422 32196 36474
rect 31950 36420 31956 36422
rect 32012 36420 32036 36422
rect 32092 36420 32116 36422
rect 32172 36420 32196 36422
rect 32252 36420 32258 36422
rect 31950 36411 32258 36420
rect 32220 36304 32272 36310
rect 32220 36246 32272 36252
rect 31852 36168 31904 36174
rect 31852 36110 31904 36116
rect 32036 36168 32088 36174
rect 32036 36110 32088 36116
rect 32048 35894 32076 36110
rect 32232 36038 32260 36246
rect 32220 36032 32272 36038
rect 32220 35974 32272 35980
rect 31864 35866 32076 35894
rect 31760 33516 31812 33522
rect 31760 33458 31812 33464
rect 31680 33238 31800 33266
rect 31576 31476 31628 31482
rect 31576 31418 31628 31424
rect 31024 29844 31076 29850
rect 31024 29786 31076 29792
rect 30840 19440 30892 19446
rect 30840 19382 30892 19388
rect 30840 16652 30892 16658
rect 30840 16594 30892 16600
rect 29736 13932 29788 13938
rect 29736 13874 29788 13880
rect 29644 11280 29696 11286
rect 29644 11222 29696 11228
rect 30852 11218 30880 16594
rect 31036 14414 31064 29786
rect 31588 28558 31616 31418
rect 31576 28552 31628 28558
rect 31576 28494 31628 28500
rect 31668 27600 31720 27606
rect 31668 27542 31720 27548
rect 31208 24744 31260 24750
rect 31208 24686 31260 24692
rect 31116 21616 31168 21622
rect 31116 21558 31168 21564
rect 31128 16658 31156 21558
rect 31116 16652 31168 16658
rect 31116 16594 31168 16600
rect 31220 15094 31248 24686
rect 31680 21622 31708 27542
rect 31668 21616 31720 21622
rect 31668 21558 31720 21564
rect 31772 21418 31800 33238
rect 31864 31278 31892 35866
rect 31950 35388 32258 35397
rect 31950 35386 31956 35388
rect 32012 35386 32036 35388
rect 32092 35386 32116 35388
rect 32172 35386 32196 35388
rect 32252 35386 32258 35388
rect 32012 35334 32014 35386
rect 32194 35334 32196 35386
rect 31950 35332 31956 35334
rect 32012 35332 32036 35334
rect 32092 35332 32116 35334
rect 32172 35332 32196 35334
rect 32252 35332 32258 35334
rect 31950 35323 32258 35332
rect 31950 34300 32258 34309
rect 31950 34298 31956 34300
rect 32012 34298 32036 34300
rect 32092 34298 32116 34300
rect 32172 34298 32196 34300
rect 32252 34298 32258 34300
rect 32012 34246 32014 34298
rect 32194 34246 32196 34298
rect 31950 34244 31956 34246
rect 32012 34244 32036 34246
rect 32092 34244 32116 34246
rect 32172 34244 32196 34246
rect 32252 34244 32258 34246
rect 31950 34235 32258 34244
rect 31950 33212 32258 33221
rect 31950 33210 31956 33212
rect 32012 33210 32036 33212
rect 32092 33210 32116 33212
rect 32172 33210 32196 33212
rect 32252 33210 32258 33212
rect 32012 33158 32014 33210
rect 32194 33158 32196 33210
rect 31950 33156 31956 33158
rect 32012 33156 32036 33158
rect 32092 33156 32116 33158
rect 32172 33156 32196 33158
rect 32252 33156 32258 33158
rect 31950 33147 32258 33156
rect 31950 32124 32258 32133
rect 31950 32122 31956 32124
rect 32012 32122 32036 32124
rect 32092 32122 32116 32124
rect 32172 32122 32196 32124
rect 32252 32122 32258 32124
rect 32012 32070 32014 32122
rect 32194 32070 32196 32122
rect 31950 32068 31956 32070
rect 32012 32068 32036 32070
rect 32092 32068 32116 32070
rect 32172 32068 32196 32070
rect 32252 32068 32258 32070
rect 31950 32059 32258 32068
rect 31852 31272 31904 31278
rect 31852 31214 31904 31220
rect 31864 28490 31892 31214
rect 31950 31036 32258 31045
rect 31950 31034 31956 31036
rect 32012 31034 32036 31036
rect 32092 31034 32116 31036
rect 32172 31034 32196 31036
rect 32252 31034 32258 31036
rect 32012 30982 32014 31034
rect 32194 30982 32196 31034
rect 31950 30980 31956 30982
rect 32012 30980 32036 30982
rect 32092 30980 32116 30982
rect 32172 30980 32196 30982
rect 32252 30980 32258 30982
rect 31950 30971 32258 30980
rect 31950 29948 32258 29957
rect 31950 29946 31956 29948
rect 32012 29946 32036 29948
rect 32092 29946 32116 29948
rect 32172 29946 32196 29948
rect 32252 29946 32258 29948
rect 32012 29894 32014 29946
rect 32194 29894 32196 29946
rect 31950 29892 31956 29894
rect 32012 29892 32036 29894
rect 32092 29892 32116 29894
rect 32172 29892 32196 29894
rect 32252 29892 32258 29894
rect 31950 29883 32258 29892
rect 31950 28860 32258 28869
rect 31950 28858 31956 28860
rect 32012 28858 32036 28860
rect 32092 28858 32116 28860
rect 32172 28858 32196 28860
rect 32252 28858 32258 28860
rect 32012 28806 32014 28858
rect 32194 28806 32196 28858
rect 31950 28804 31956 28806
rect 32012 28804 32036 28806
rect 32092 28804 32116 28806
rect 32172 28804 32196 28806
rect 32252 28804 32258 28806
rect 31950 28795 32258 28804
rect 31852 28484 31904 28490
rect 31852 28426 31904 28432
rect 31852 28212 31904 28218
rect 31852 28154 31904 28160
rect 31864 25974 31892 28154
rect 31950 27772 32258 27781
rect 31950 27770 31956 27772
rect 32012 27770 32036 27772
rect 32092 27770 32116 27772
rect 32172 27770 32196 27772
rect 32252 27770 32258 27772
rect 32012 27718 32014 27770
rect 32194 27718 32196 27770
rect 31950 27716 31956 27718
rect 32012 27716 32036 27718
rect 32092 27716 32116 27718
rect 32172 27716 32196 27718
rect 32252 27716 32258 27718
rect 31950 27707 32258 27716
rect 31950 26684 32258 26693
rect 31950 26682 31956 26684
rect 32012 26682 32036 26684
rect 32092 26682 32116 26684
rect 32172 26682 32196 26684
rect 32252 26682 32258 26684
rect 32012 26630 32014 26682
rect 32194 26630 32196 26682
rect 31950 26628 31956 26630
rect 32012 26628 32036 26630
rect 32092 26628 32116 26630
rect 32172 26628 32196 26630
rect 32252 26628 32258 26630
rect 31950 26619 32258 26628
rect 31852 25968 31904 25974
rect 31852 25910 31904 25916
rect 32324 25770 32352 51954
rect 32404 37868 32456 37874
rect 32404 37810 32456 37816
rect 32416 36242 32444 37810
rect 32404 36236 32456 36242
rect 32404 36178 32456 36184
rect 32404 36100 32456 36106
rect 32404 36042 32456 36048
rect 32416 30326 32444 36042
rect 32404 30320 32456 30326
rect 32404 30262 32456 30268
rect 32416 28218 32444 30262
rect 32404 28212 32456 28218
rect 32404 28154 32456 28160
rect 32508 27402 32536 63718
rect 32610 63132 32918 63141
rect 32610 63130 32616 63132
rect 32672 63130 32696 63132
rect 32752 63130 32776 63132
rect 32832 63130 32856 63132
rect 32912 63130 32918 63132
rect 32672 63078 32674 63130
rect 32854 63078 32856 63130
rect 32610 63076 32616 63078
rect 32672 63076 32696 63078
rect 32752 63076 32776 63078
rect 32832 63076 32856 63078
rect 32912 63076 32918 63078
rect 32610 63067 32918 63076
rect 32610 62044 32918 62053
rect 32610 62042 32616 62044
rect 32672 62042 32696 62044
rect 32752 62042 32776 62044
rect 32832 62042 32856 62044
rect 32912 62042 32918 62044
rect 32672 61990 32674 62042
rect 32854 61990 32856 62042
rect 32610 61988 32616 61990
rect 32672 61988 32696 61990
rect 32752 61988 32776 61990
rect 32832 61988 32856 61990
rect 32912 61988 32918 61990
rect 32610 61979 32918 61988
rect 32610 60956 32918 60965
rect 32610 60954 32616 60956
rect 32672 60954 32696 60956
rect 32752 60954 32776 60956
rect 32832 60954 32856 60956
rect 32912 60954 32918 60956
rect 32672 60902 32674 60954
rect 32854 60902 32856 60954
rect 32610 60900 32616 60902
rect 32672 60900 32696 60902
rect 32752 60900 32776 60902
rect 32832 60900 32856 60902
rect 32912 60900 32918 60902
rect 32610 60891 32918 60900
rect 32610 59868 32918 59877
rect 32610 59866 32616 59868
rect 32672 59866 32696 59868
rect 32752 59866 32776 59868
rect 32832 59866 32856 59868
rect 32912 59866 32918 59868
rect 32672 59814 32674 59866
rect 32854 59814 32856 59866
rect 32610 59812 32616 59814
rect 32672 59812 32696 59814
rect 32752 59812 32776 59814
rect 32832 59812 32856 59814
rect 32912 59812 32918 59814
rect 32610 59803 32918 59812
rect 32610 58780 32918 58789
rect 32610 58778 32616 58780
rect 32672 58778 32696 58780
rect 32752 58778 32776 58780
rect 32832 58778 32856 58780
rect 32912 58778 32918 58780
rect 32672 58726 32674 58778
rect 32854 58726 32856 58778
rect 32610 58724 32616 58726
rect 32672 58724 32696 58726
rect 32752 58724 32776 58726
rect 32832 58724 32856 58726
rect 32912 58724 32918 58726
rect 32610 58715 32918 58724
rect 32610 57692 32918 57701
rect 32610 57690 32616 57692
rect 32672 57690 32696 57692
rect 32752 57690 32776 57692
rect 32832 57690 32856 57692
rect 32912 57690 32918 57692
rect 32672 57638 32674 57690
rect 32854 57638 32856 57690
rect 32610 57636 32616 57638
rect 32672 57636 32696 57638
rect 32752 57636 32776 57638
rect 32832 57636 32856 57638
rect 32912 57636 32918 57638
rect 32610 57627 32918 57636
rect 32610 56604 32918 56613
rect 32610 56602 32616 56604
rect 32672 56602 32696 56604
rect 32752 56602 32776 56604
rect 32832 56602 32856 56604
rect 32912 56602 32918 56604
rect 32672 56550 32674 56602
rect 32854 56550 32856 56602
rect 32610 56548 32616 56550
rect 32672 56548 32696 56550
rect 32752 56548 32776 56550
rect 32832 56548 32856 56550
rect 32912 56548 32918 56550
rect 32610 56539 32918 56548
rect 32610 55516 32918 55525
rect 32610 55514 32616 55516
rect 32672 55514 32696 55516
rect 32752 55514 32776 55516
rect 32832 55514 32856 55516
rect 32912 55514 32918 55516
rect 32672 55462 32674 55514
rect 32854 55462 32856 55514
rect 32610 55460 32616 55462
rect 32672 55460 32696 55462
rect 32752 55460 32776 55462
rect 32832 55460 32856 55462
rect 32912 55460 32918 55462
rect 32610 55451 32918 55460
rect 32610 54428 32918 54437
rect 32610 54426 32616 54428
rect 32672 54426 32696 54428
rect 32752 54426 32776 54428
rect 32832 54426 32856 54428
rect 32912 54426 32918 54428
rect 32672 54374 32674 54426
rect 32854 54374 32856 54426
rect 32610 54372 32616 54374
rect 32672 54372 32696 54374
rect 32752 54372 32776 54374
rect 32832 54372 32856 54374
rect 32912 54372 32918 54374
rect 32610 54363 32918 54372
rect 32610 53340 32918 53349
rect 32610 53338 32616 53340
rect 32672 53338 32696 53340
rect 32752 53338 32776 53340
rect 32832 53338 32856 53340
rect 32912 53338 32918 53340
rect 32672 53286 32674 53338
rect 32854 53286 32856 53338
rect 32610 53284 32616 53286
rect 32672 53284 32696 53286
rect 32752 53284 32776 53286
rect 32832 53284 32856 53286
rect 32912 53284 32918 53286
rect 32610 53275 32918 53284
rect 33152 52630 33180 69362
rect 36950 69116 37258 69125
rect 36950 69114 36956 69116
rect 37012 69114 37036 69116
rect 37092 69114 37116 69116
rect 37172 69114 37196 69116
rect 37252 69114 37258 69116
rect 37012 69062 37014 69114
rect 37194 69062 37196 69114
rect 36950 69060 36956 69062
rect 37012 69060 37036 69062
rect 37092 69060 37116 69062
rect 37172 69060 37196 69062
rect 37252 69060 37258 69062
rect 36950 69051 37258 69060
rect 36176 68876 36228 68882
rect 36176 68818 36228 68824
rect 35992 68740 36044 68746
rect 35992 68682 36044 68688
rect 34152 68264 34204 68270
rect 34152 68206 34204 68212
rect 34164 67658 34192 68206
rect 34152 67652 34204 67658
rect 34152 67594 34204 67600
rect 34520 67652 34572 67658
rect 34520 67594 34572 67600
rect 33232 63368 33284 63374
rect 33232 63310 33284 63316
rect 33244 58342 33272 63310
rect 33232 58336 33284 58342
rect 33230 58304 33232 58313
rect 33284 58304 33286 58313
rect 33230 58239 33286 58248
rect 34164 56506 34192 67594
rect 33416 56500 33468 56506
rect 33416 56442 33468 56448
rect 34152 56500 34204 56506
rect 34152 56442 34204 56448
rect 33428 55690 33456 56442
rect 33692 56432 33744 56438
rect 33692 56374 33744 56380
rect 33876 56432 33928 56438
rect 33876 56374 33928 56380
rect 33508 56160 33560 56166
rect 33508 56102 33560 56108
rect 33600 56160 33652 56166
rect 33600 56102 33652 56108
rect 33520 55729 33548 56102
rect 33506 55720 33562 55729
rect 33416 55684 33468 55690
rect 33506 55655 33562 55664
rect 33416 55626 33468 55632
rect 33428 55214 33456 55626
rect 33428 55186 33548 55214
rect 33140 52624 33192 52630
rect 33140 52566 33192 52572
rect 32610 52252 32918 52261
rect 32610 52250 32616 52252
rect 32672 52250 32696 52252
rect 32752 52250 32776 52252
rect 32832 52250 32856 52252
rect 32912 52250 32918 52252
rect 32672 52198 32674 52250
rect 32854 52198 32856 52250
rect 32610 52196 32616 52198
rect 32672 52196 32696 52198
rect 32752 52196 32776 52198
rect 32832 52196 32856 52198
rect 32912 52196 32918 52198
rect 32610 52187 32918 52196
rect 33048 51876 33100 51882
rect 33048 51818 33100 51824
rect 32610 51164 32918 51173
rect 32610 51162 32616 51164
rect 32672 51162 32696 51164
rect 32752 51162 32776 51164
rect 32832 51162 32856 51164
rect 32912 51162 32918 51164
rect 32672 51110 32674 51162
rect 32854 51110 32856 51162
rect 32610 51108 32616 51110
rect 32672 51108 32696 51110
rect 32752 51108 32776 51110
rect 32832 51108 32856 51110
rect 32912 51108 32918 51110
rect 32610 51099 32918 51108
rect 32610 50076 32918 50085
rect 32610 50074 32616 50076
rect 32672 50074 32696 50076
rect 32752 50074 32776 50076
rect 32832 50074 32856 50076
rect 32912 50074 32918 50076
rect 32672 50022 32674 50074
rect 32854 50022 32856 50074
rect 32610 50020 32616 50022
rect 32672 50020 32696 50022
rect 32752 50020 32776 50022
rect 32832 50020 32856 50022
rect 32912 50020 32918 50022
rect 32610 50011 32918 50020
rect 32610 48988 32918 48997
rect 32610 48986 32616 48988
rect 32672 48986 32696 48988
rect 32752 48986 32776 48988
rect 32832 48986 32856 48988
rect 32912 48986 32918 48988
rect 32672 48934 32674 48986
rect 32854 48934 32856 48986
rect 32610 48932 32616 48934
rect 32672 48932 32696 48934
rect 32752 48932 32776 48934
rect 32832 48932 32856 48934
rect 32912 48932 32918 48934
rect 32610 48923 32918 48932
rect 32610 47900 32918 47909
rect 32610 47898 32616 47900
rect 32672 47898 32696 47900
rect 32752 47898 32776 47900
rect 32832 47898 32856 47900
rect 32912 47898 32918 47900
rect 32672 47846 32674 47898
rect 32854 47846 32856 47898
rect 32610 47844 32616 47846
rect 32672 47844 32696 47846
rect 32752 47844 32776 47846
rect 32832 47844 32856 47846
rect 32912 47844 32918 47846
rect 32610 47835 32918 47844
rect 33060 47190 33088 51818
rect 33140 51808 33192 51814
rect 33140 51750 33192 51756
rect 33152 51270 33180 51750
rect 33140 51264 33192 51270
rect 33138 51232 33140 51241
rect 33192 51232 33194 51241
rect 33138 51167 33194 51176
rect 33416 49428 33468 49434
rect 33416 49370 33468 49376
rect 33324 49156 33376 49162
rect 33324 49098 33376 49104
rect 33140 49088 33192 49094
rect 33140 49030 33192 49036
rect 33048 47184 33100 47190
rect 33048 47126 33100 47132
rect 32610 46812 32918 46821
rect 32610 46810 32616 46812
rect 32672 46810 32696 46812
rect 32752 46810 32776 46812
rect 32832 46810 32856 46812
rect 32912 46810 32918 46812
rect 32672 46758 32674 46810
rect 32854 46758 32856 46810
rect 32610 46756 32616 46758
rect 32672 46756 32696 46758
rect 32752 46756 32776 46758
rect 32832 46756 32856 46758
rect 32912 46756 32918 46758
rect 32610 46747 32918 46756
rect 32610 45724 32918 45733
rect 32610 45722 32616 45724
rect 32672 45722 32696 45724
rect 32752 45722 32776 45724
rect 32832 45722 32856 45724
rect 32912 45722 32918 45724
rect 32672 45670 32674 45722
rect 32854 45670 32856 45722
rect 32610 45668 32616 45670
rect 32672 45668 32696 45670
rect 32752 45668 32776 45670
rect 32832 45668 32856 45670
rect 32912 45668 32918 45670
rect 32610 45659 32918 45668
rect 32610 44636 32918 44645
rect 32610 44634 32616 44636
rect 32672 44634 32696 44636
rect 32752 44634 32776 44636
rect 32832 44634 32856 44636
rect 32912 44634 32918 44636
rect 32672 44582 32674 44634
rect 32854 44582 32856 44634
rect 32610 44580 32616 44582
rect 32672 44580 32696 44582
rect 32752 44580 32776 44582
rect 32832 44580 32856 44582
rect 32912 44580 32918 44582
rect 32610 44571 32918 44580
rect 32610 43548 32918 43557
rect 32610 43546 32616 43548
rect 32672 43546 32696 43548
rect 32752 43546 32776 43548
rect 32832 43546 32856 43548
rect 32912 43546 32918 43548
rect 32672 43494 32674 43546
rect 32854 43494 32856 43546
rect 32610 43492 32616 43494
rect 32672 43492 32696 43494
rect 32752 43492 32776 43494
rect 32832 43492 32856 43494
rect 32912 43492 32918 43494
rect 32610 43483 32918 43492
rect 32610 42460 32918 42469
rect 32610 42458 32616 42460
rect 32672 42458 32696 42460
rect 32752 42458 32776 42460
rect 32832 42458 32856 42460
rect 32912 42458 32918 42460
rect 32672 42406 32674 42458
rect 32854 42406 32856 42458
rect 32610 42404 32616 42406
rect 32672 42404 32696 42406
rect 32752 42404 32776 42406
rect 32832 42404 32856 42406
rect 32912 42404 32918 42406
rect 32610 42395 32918 42404
rect 32610 41372 32918 41381
rect 32610 41370 32616 41372
rect 32672 41370 32696 41372
rect 32752 41370 32776 41372
rect 32832 41370 32856 41372
rect 32912 41370 32918 41372
rect 32672 41318 32674 41370
rect 32854 41318 32856 41370
rect 32610 41316 32616 41318
rect 32672 41316 32696 41318
rect 32752 41316 32776 41318
rect 32832 41316 32856 41318
rect 32912 41316 32918 41318
rect 32610 41307 32918 41316
rect 32610 40284 32918 40293
rect 32610 40282 32616 40284
rect 32672 40282 32696 40284
rect 32752 40282 32776 40284
rect 32832 40282 32856 40284
rect 32912 40282 32918 40284
rect 32672 40230 32674 40282
rect 32854 40230 32856 40282
rect 32610 40228 32616 40230
rect 32672 40228 32696 40230
rect 32752 40228 32776 40230
rect 32832 40228 32856 40230
rect 32912 40228 32918 40230
rect 32610 40219 32918 40228
rect 32610 39196 32918 39205
rect 32610 39194 32616 39196
rect 32672 39194 32696 39196
rect 32752 39194 32776 39196
rect 32832 39194 32856 39196
rect 32912 39194 32918 39196
rect 32672 39142 32674 39194
rect 32854 39142 32856 39194
rect 32610 39140 32616 39142
rect 32672 39140 32696 39142
rect 32752 39140 32776 39142
rect 32832 39140 32856 39142
rect 32912 39140 32918 39142
rect 32610 39131 32918 39140
rect 32610 38108 32918 38117
rect 32610 38106 32616 38108
rect 32672 38106 32696 38108
rect 32752 38106 32776 38108
rect 32832 38106 32856 38108
rect 32912 38106 32918 38108
rect 32672 38054 32674 38106
rect 32854 38054 32856 38106
rect 32610 38052 32616 38054
rect 32672 38052 32696 38054
rect 32752 38052 32776 38054
rect 32832 38052 32856 38054
rect 32912 38052 32918 38054
rect 32610 38043 32918 38052
rect 32610 37020 32918 37029
rect 32610 37018 32616 37020
rect 32672 37018 32696 37020
rect 32752 37018 32776 37020
rect 32832 37018 32856 37020
rect 32912 37018 32918 37020
rect 32672 36966 32674 37018
rect 32854 36966 32856 37018
rect 32610 36964 32616 36966
rect 32672 36964 32696 36966
rect 32752 36964 32776 36966
rect 32832 36964 32856 36966
rect 32912 36964 32918 36966
rect 32610 36955 32918 36964
rect 33048 36236 33100 36242
rect 33048 36178 33100 36184
rect 32956 36032 33008 36038
rect 32956 35974 33008 35980
rect 32610 35932 32918 35941
rect 32610 35930 32616 35932
rect 32672 35930 32696 35932
rect 32752 35930 32776 35932
rect 32832 35930 32856 35932
rect 32912 35930 32918 35932
rect 32672 35878 32674 35930
rect 32854 35878 32856 35930
rect 32610 35876 32616 35878
rect 32672 35876 32696 35878
rect 32752 35876 32776 35878
rect 32832 35876 32856 35878
rect 32912 35876 32918 35878
rect 32610 35867 32918 35876
rect 32610 34844 32918 34853
rect 32610 34842 32616 34844
rect 32672 34842 32696 34844
rect 32752 34842 32776 34844
rect 32832 34842 32856 34844
rect 32912 34842 32918 34844
rect 32672 34790 32674 34842
rect 32854 34790 32856 34842
rect 32610 34788 32616 34790
rect 32672 34788 32696 34790
rect 32752 34788 32776 34790
rect 32832 34788 32856 34790
rect 32912 34788 32918 34790
rect 32610 34779 32918 34788
rect 32610 33756 32918 33765
rect 32610 33754 32616 33756
rect 32672 33754 32696 33756
rect 32752 33754 32776 33756
rect 32832 33754 32856 33756
rect 32912 33754 32918 33756
rect 32672 33702 32674 33754
rect 32854 33702 32856 33754
rect 32610 33700 32616 33702
rect 32672 33700 32696 33702
rect 32752 33700 32776 33702
rect 32832 33700 32856 33702
rect 32912 33700 32918 33702
rect 32610 33691 32918 33700
rect 32610 32668 32918 32677
rect 32610 32666 32616 32668
rect 32672 32666 32696 32668
rect 32752 32666 32776 32668
rect 32832 32666 32856 32668
rect 32912 32666 32918 32668
rect 32672 32614 32674 32666
rect 32854 32614 32856 32666
rect 32610 32612 32616 32614
rect 32672 32612 32696 32614
rect 32752 32612 32776 32614
rect 32832 32612 32856 32614
rect 32912 32612 32918 32614
rect 32610 32603 32918 32612
rect 32610 31580 32918 31589
rect 32610 31578 32616 31580
rect 32672 31578 32696 31580
rect 32752 31578 32776 31580
rect 32832 31578 32856 31580
rect 32912 31578 32918 31580
rect 32672 31526 32674 31578
rect 32854 31526 32856 31578
rect 32610 31524 32616 31526
rect 32672 31524 32696 31526
rect 32752 31524 32776 31526
rect 32832 31524 32856 31526
rect 32912 31524 32918 31526
rect 32610 31515 32918 31524
rect 32610 30492 32918 30501
rect 32610 30490 32616 30492
rect 32672 30490 32696 30492
rect 32752 30490 32776 30492
rect 32832 30490 32856 30492
rect 32912 30490 32918 30492
rect 32672 30438 32674 30490
rect 32854 30438 32856 30490
rect 32610 30436 32616 30438
rect 32672 30436 32696 30438
rect 32752 30436 32776 30438
rect 32832 30436 32856 30438
rect 32912 30436 32918 30438
rect 32610 30427 32918 30436
rect 32610 29404 32918 29413
rect 32610 29402 32616 29404
rect 32672 29402 32696 29404
rect 32752 29402 32776 29404
rect 32832 29402 32856 29404
rect 32912 29402 32918 29404
rect 32672 29350 32674 29402
rect 32854 29350 32856 29402
rect 32610 29348 32616 29350
rect 32672 29348 32696 29350
rect 32752 29348 32776 29350
rect 32832 29348 32856 29350
rect 32912 29348 32918 29350
rect 32610 29339 32918 29348
rect 32610 28316 32918 28325
rect 32610 28314 32616 28316
rect 32672 28314 32696 28316
rect 32752 28314 32776 28316
rect 32832 28314 32856 28316
rect 32912 28314 32918 28316
rect 32672 28262 32674 28314
rect 32854 28262 32856 28314
rect 32610 28260 32616 28262
rect 32672 28260 32696 28262
rect 32752 28260 32776 28262
rect 32832 28260 32856 28262
rect 32912 28260 32918 28262
rect 32610 28251 32918 28260
rect 32496 27396 32548 27402
rect 32496 27338 32548 27344
rect 32610 27228 32918 27237
rect 32610 27226 32616 27228
rect 32672 27226 32696 27228
rect 32752 27226 32776 27228
rect 32832 27226 32856 27228
rect 32912 27226 32918 27228
rect 32672 27174 32674 27226
rect 32854 27174 32856 27226
rect 32610 27172 32616 27174
rect 32672 27172 32696 27174
rect 32752 27172 32776 27174
rect 32832 27172 32856 27174
rect 32912 27172 32918 27174
rect 32610 27163 32918 27172
rect 32610 26140 32918 26149
rect 32610 26138 32616 26140
rect 32672 26138 32696 26140
rect 32752 26138 32776 26140
rect 32832 26138 32856 26140
rect 32912 26138 32918 26140
rect 32672 26086 32674 26138
rect 32854 26086 32856 26138
rect 32610 26084 32616 26086
rect 32672 26084 32696 26086
rect 32752 26084 32776 26086
rect 32832 26084 32856 26086
rect 32912 26084 32918 26086
rect 32610 26075 32918 26084
rect 32968 25906 32996 35974
rect 32956 25900 33008 25906
rect 32956 25842 33008 25848
rect 33060 25838 33088 36178
rect 33048 25832 33100 25838
rect 33048 25774 33100 25780
rect 32312 25764 32364 25770
rect 32312 25706 32364 25712
rect 31950 25596 32258 25605
rect 31950 25594 31956 25596
rect 32012 25594 32036 25596
rect 32092 25594 32116 25596
rect 32172 25594 32196 25596
rect 32252 25594 32258 25596
rect 32012 25542 32014 25594
rect 32194 25542 32196 25594
rect 31950 25540 31956 25542
rect 32012 25540 32036 25542
rect 32092 25540 32116 25542
rect 32172 25540 32196 25542
rect 32252 25540 32258 25542
rect 31950 25531 32258 25540
rect 32610 25052 32918 25061
rect 32610 25050 32616 25052
rect 32672 25050 32696 25052
rect 32752 25050 32776 25052
rect 32832 25050 32856 25052
rect 32912 25050 32918 25052
rect 32672 24998 32674 25050
rect 32854 24998 32856 25050
rect 32610 24996 32616 24998
rect 32672 24996 32696 24998
rect 32752 24996 32776 24998
rect 32832 24996 32856 24998
rect 32912 24996 32918 24998
rect 32610 24987 32918 24996
rect 31950 24508 32258 24517
rect 31950 24506 31956 24508
rect 32012 24506 32036 24508
rect 32092 24506 32116 24508
rect 32172 24506 32196 24508
rect 32252 24506 32258 24508
rect 32012 24454 32014 24506
rect 32194 24454 32196 24506
rect 31950 24452 31956 24454
rect 32012 24452 32036 24454
rect 32092 24452 32116 24454
rect 32172 24452 32196 24454
rect 32252 24452 32258 24454
rect 31950 24443 32258 24452
rect 32610 23964 32918 23973
rect 32610 23962 32616 23964
rect 32672 23962 32696 23964
rect 32752 23962 32776 23964
rect 32832 23962 32856 23964
rect 32912 23962 32918 23964
rect 32672 23910 32674 23962
rect 32854 23910 32856 23962
rect 32610 23908 32616 23910
rect 32672 23908 32696 23910
rect 32752 23908 32776 23910
rect 32832 23908 32856 23910
rect 32912 23908 32918 23910
rect 32610 23899 32918 23908
rect 31950 23420 32258 23429
rect 31950 23418 31956 23420
rect 32012 23418 32036 23420
rect 32092 23418 32116 23420
rect 32172 23418 32196 23420
rect 32252 23418 32258 23420
rect 32012 23366 32014 23418
rect 32194 23366 32196 23418
rect 31950 23364 31956 23366
rect 32012 23364 32036 23366
rect 32092 23364 32116 23366
rect 32172 23364 32196 23366
rect 32252 23364 32258 23366
rect 31950 23355 32258 23364
rect 32610 22876 32918 22885
rect 32610 22874 32616 22876
rect 32672 22874 32696 22876
rect 32752 22874 32776 22876
rect 32832 22874 32856 22876
rect 32912 22874 32918 22876
rect 32672 22822 32674 22874
rect 32854 22822 32856 22874
rect 32610 22820 32616 22822
rect 32672 22820 32696 22822
rect 32752 22820 32776 22822
rect 32832 22820 32856 22822
rect 32912 22820 32918 22822
rect 32610 22811 32918 22820
rect 31950 22332 32258 22341
rect 31950 22330 31956 22332
rect 32012 22330 32036 22332
rect 32092 22330 32116 22332
rect 32172 22330 32196 22332
rect 32252 22330 32258 22332
rect 32012 22278 32014 22330
rect 32194 22278 32196 22330
rect 31950 22276 31956 22278
rect 32012 22276 32036 22278
rect 32092 22276 32116 22278
rect 32172 22276 32196 22278
rect 32252 22276 32258 22278
rect 31950 22267 32258 22276
rect 32610 21788 32918 21797
rect 32610 21786 32616 21788
rect 32672 21786 32696 21788
rect 32752 21786 32776 21788
rect 32832 21786 32856 21788
rect 32912 21786 32918 21788
rect 32672 21734 32674 21786
rect 32854 21734 32856 21786
rect 32610 21732 32616 21734
rect 32672 21732 32696 21734
rect 32752 21732 32776 21734
rect 32832 21732 32856 21734
rect 32912 21732 32918 21734
rect 32610 21723 32918 21732
rect 31760 21412 31812 21418
rect 31760 21354 31812 21360
rect 32404 21344 32456 21350
rect 32404 21286 32456 21292
rect 31950 21244 32258 21253
rect 31950 21242 31956 21244
rect 32012 21242 32036 21244
rect 32092 21242 32116 21244
rect 32172 21242 32196 21244
rect 32252 21242 32258 21244
rect 32012 21190 32014 21242
rect 32194 21190 32196 21242
rect 31950 21188 31956 21190
rect 32012 21188 32036 21190
rect 32092 21188 32116 21190
rect 32172 21188 32196 21190
rect 32252 21188 32258 21190
rect 31950 21179 32258 21188
rect 31950 20156 32258 20165
rect 31950 20154 31956 20156
rect 32012 20154 32036 20156
rect 32092 20154 32116 20156
rect 32172 20154 32196 20156
rect 32252 20154 32258 20156
rect 32012 20102 32014 20154
rect 32194 20102 32196 20154
rect 31950 20100 31956 20102
rect 32012 20100 32036 20102
rect 32092 20100 32116 20102
rect 32172 20100 32196 20102
rect 32252 20100 32258 20102
rect 31950 20091 32258 20100
rect 31950 19068 32258 19077
rect 31950 19066 31956 19068
rect 32012 19066 32036 19068
rect 32092 19066 32116 19068
rect 32172 19066 32196 19068
rect 32252 19066 32258 19068
rect 32012 19014 32014 19066
rect 32194 19014 32196 19066
rect 31950 19012 31956 19014
rect 32012 19012 32036 19014
rect 32092 19012 32116 19014
rect 32172 19012 32196 19014
rect 32252 19012 32258 19014
rect 31950 19003 32258 19012
rect 31950 17980 32258 17989
rect 31950 17978 31956 17980
rect 32012 17978 32036 17980
rect 32092 17978 32116 17980
rect 32172 17978 32196 17980
rect 32252 17978 32258 17980
rect 32012 17926 32014 17978
rect 32194 17926 32196 17978
rect 31950 17924 31956 17926
rect 32012 17924 32036 17926
rect 32092 17924 32116 17926
rect 32172 17924 32196 17926
rect 32252 17924 32258 17926
rect 31950 17915 32258 17924
rect 31950 16892 32258 16901
rect 31950 16890 31956 16892
rect 32012 16890 32036 16892
rect 32092 16890 32116 16892
rect 32172 16890 32196 16892
rect 32252 16890 32258 16892
rect 32012 16838 32014 16890
rect 32194 16838 32196 16890
rect 31950 16836 31956 16838
rect 32012 16836 32036 16838
rect 32092 16836 32116 16838
rect 32172 16836 32196 16838
rect 32252 16836 32258 16838
rect 31950 16827 32258 16836
rect 31950 15804 32258 15813
rect 31950 15802 31956 15804
rect 32012 15802 32036 15804
rect 32092 15802 32116 15804
rect 32172 15802 32196 15804
rect 32252 15802 32258 15804
rect 32012 15750 32014 15802
rect 32194 15750 32196 15802
rect 31950 15748 31956 15750
rect 32012 15748 32036 15750
rect 32092 15748 32116 15750
rect 32172 15748 32196 15750
rect 32252 15748 32258 15750
rect 31950 15739 32258 15748
rect 32416 15094 32444 21286
rect 32610 20700 32918 20709
rect 32610 20698 32616 20700
rect 32672 20698 32696 20700
rect 32752 20698 32776 20700
rect 32832 20698 32856 20700
rect 32912 20698 32918 20700
rect 32672 20646 32674 20698
rect 32854 20646 32856 20698
rect 32610 20644 32616 20646
rect 32672 20644 32696 20646
rect 32752 20644 32776 20646
rect 32832 20644 32856 20646
rect 32912 20644 32918 20646
rect 32610 20635 32918 20644
rect 32610 19612 32918 19621
rect 32610 19610 32616 19612
rect 32672 19610 32696 19612
rect 32752 19610 32776 19612
rect 32832 19610 32856 19612
rect 32912 19610 32918 19612
rect 32672 19558 32674 19610
rect 32854 19558 32856 19610
rect 32610 19556 32616 19558
rect 32672 19556 32696 19558
rect 32752 19556 32776 19558
rect 32832 19556 32856 19558
rect 32912 19556 32918 19558
rect 32610 19547 32918 19556
rect 32610 18524 32918 18533
rect 32610 18522 32616 18524
rect 32672 18522 32696 18524
rect 32752 18522 32776 18524
rect 32832 18522 32856 18524
rect 32912 18522 32918 18524
rect 32672 18470 32674 18522
rect 32854 18470 32856 18522
rect 32610 18468 32616 18470
rect 32672 18468 32696 18470
rect 32752 18468 32776 18470
rect 32832 18468 32856 18470
rect 32912 18468 32918 18470
rect 32610 18459 32918 18468
rect 32610 17436 32918 17445
rect 32610 17434 32616 17436
rect 32672 17434 32696 17436
rect 32752 17434 32776 17436
rect 32832 17434 32856 17436
rect 32912 17434 32918 17436
rect 32672 17382 32674 17434
rect 32854 17382 32856 17434
rect 32610 17380 32616 17382
rect 32672 17380 32696 17382
rect 32752 17380 32776 17382
rect 32832 17380 32856 17382
rect 32912 17380 32918 17382
rect 32610 17371 32918 17380
rect 32610 16348 32918 16357
rect 32610 16346 32616 16348
rect 32672 16346 32696 16348
rect 32752 16346 32776 16348
rect 32832 16346 32856 16348
rect 32912 16346 32918 16348
rect 32672 16294 32674 16346
rect 32854 16294 32856 16346
rect 32610 16292 32616 16294
rect 32672 16292 32696 16294
rect 32752 16292 32776 16294
rect 32832 16292 32856 16294
rect 32912 16292 32918 16294
rect 32610 16283 32918 16292
rect 32610 15260 32918 15269
rect 32610 15258 32616 15260
rect 32672 15258 32696 15260
rect 32752 15258 32776 15260
rect 32832 15258 32856 15260
rect 32912 15258 32918 15260
rect 32672 15206 32674 15258
rect 32854 15206 32856 15258
rect 32610 15204 32616 15206
rect 32672 15204 32696 15206
rect 32752 15204 32776 15206
rect 32832 15204 32856 15206
rect 32912 15204 32918 15206
rect 32610 15195 32918 15204
rect 31208 15088 31260 15094
rect 31208 15030 31260 15036
rect 32404 15088 32456 15094
rect 32404 15030 32456 15036
rect 31950 14716 32258 14725
rect 31950 14714 31956 14716
rect 32012 14714 32036 14716
rect 32092 14714 32116 14716
rect 32172 14714 32196 14716
rect 32252 14714 32258 14716
rect 32012 14662 32014 14714
rect 32194 14662 32196 14714
rect 31950 14660 31956 14662
rect 32012 14660 32036 14662
rect 32092 14660 32116 14662
rect 32172 14660 32196 14662
rect 32252 14660 32258 14662
rect 31950 14651 32258 14660
rect 31024 14408 31076 14414
rect 31024 14350 31076 14356
rect 32610 14172 32918 14181
rect 32610 14170 32616 14172
rect 32672 14170 32696 14172
rect 32752 14170 32776 14172
rect 32832 14170 32856 14172
rect 32912 14170 32918 14172
rect 32672 14118 32674 14170
rect 32854 14118 32856 14170
rect 32610 14116 32616 14118
rect 32672 14116 32696 14118
rect 32752 14116 32776 14118
rect 32832 14116 32856 14118
rect 32912 14116 32918 14118
rect 32610 14107 32918 14116
rect 31950 13628 32258 13637
rect 31950 13626 31956 13628
rect 32012 13626 32036 13628
rect 32092 13626 32116 13628
rect 32172 13626 32196 13628
rect 32252 13626 32258 13628
rect 32012 13574 32014 13626
rect 32194 13574 32196 13626
rect 31950 13572 31956 13574
rect 32012 13572 32036 13574
rect 32092 13572 32116 13574
rect 32172 13572 32196 13574
rect 32252 13572 32258 13574
rect 31950 13563 32258 13572
rect 32610 13084 32918 13093
rect 32610 13082 32616 13084
rect 32672 13082 32696 13084
rect 32752 13082 32776 13084
rect 32832 13082 32856 13084
rect 32912 13082 32918 13084
rect 32672 13030 32674 13082
rect 32854 13030 32856 13082
rect 32610 13028 32616 13030
rect 32672 13028 32696 13030
rect 32752 13028 32776 13030
rect 32832 13028 32856 13030
rect 32912 13028 32918 13030
rect 32610 13019 32918 13028
rect 31950 12540 32258 12549
rect 31950 12538 31956 12540
rect 32012 12538 32036 12540
rect 32092 12538 32116 12540
rect 32172 12538 32196 12540
rect 32252 12538 32258 12540
rect 32012 12486 32014 12538
rect 32194 12486 32196 12538
rect 31950 12484 31956 12486
rect 32012 12484 32036 12486
rect 32092 12484 32116 12486
rect 32172 12484 32196 12486
rect 32252 12484 32258 12486
rect 31950 12475 32258 12484
rect 32610 11996 32918 12005
rect 32610 11994 32616 11996
rect 32672 11994 32696 11996
rect 32752 11994 32776 11996
rect 32832 11994 32856 11996
rect 32912 11994 32918 11996
rect 32672 11942 32674 11994
rect 32854 11942 32856 11994
rect 32610 11940 32616 11942
rect 32672 11940 32696 11942
rect 32752 11940 32776 11942
rect 32832 11940 32856 11942
rect 32912 11940 32918 11942
rect 32610 11931 32918 11940
rect 31950 11452 32258 11461
rect 31950 11450 31956 11452
rect 32012 11450 32036 11452
rect 32092 11450 32116 11452
rect 32172 11450 32196 11452
rect 32252 11450 32258 11452
rect 32012 11398 32014 11450
rect 32194 11398 32196 11450
rect 31950 11396 31956 11398
rect 32012 11396 32036 11398
rect 32092 11396 32116 11398
rect 32172 11396 32196 11398
rect 32252 11396 32258 11398
rect 31950 11387 32258 11396
rect 33060 11218 33088 25774
rect 33152 12866 33180 49030
rect 33232 31204 33284 31210
rect 33232 31146 33284 31152
rect 33244 30734 33272 31146
rect 33232 30728 33284 30734
rect 33232 30670 33284 30676
rect 33232 23792 33284 23798
rect 33232 23734 33284 23740
rect 33244 15366 33272 23734
rect 33232 15360 33284 15366
rect 33232 15302 33284 15308
rect 33336 14890 33364 49098
rect 33428 48346 33456 49370
rect 33416 48340 33468 48346
rect 33416 48282 33468 48288
rect 33428 23526 33456 48282
rect 33520 31142 33548 55186
rect 33612 49434 33640 56102
rect 33600 49428 33652 49434
rect 33600 49370 33652 49376
rect 33600 48204 33652 48210
rect 33600 48146 33652 48152
rect 33612 31414 33640 48146
rect 33600 31408 33652 31414
rect 33600 31350 33652 31356
rect 33508 31136 33560 31142
rect 33508 31078 33560 31084
rect 33612 28626 33640 31350
rect 33704 29306 33732 56374
rect 33888 55865 33916 56374
rect 33874 55856 33930 55865
rect 33874 55791 33930 55800
rect 34532 55214 34560 67594
rect 35440 65000 35492 65006
rect 35440 64942 35492 64948
rect 35452 58478 35480 64942
rect 35440 58472 35492 58478
rect 35440 58414 35492 58420
rect 34532 55186 34652 55214
rect 34520 53508 34572 53514
rect 34520 53450 34572 53456
rect 34152 52352 34204 52358
rect 34152 52294 34204 52300
rect 34164 51610 34192 52294
rect 34152 51604 34204 51610
rect 34152 51546 34204 51552
rect 34164 50250 34192 51546
rect 34532 51338 34560 53450
rect 34520 51332 34572 51338
rect 34520 51274 34572 51280
rect 34152 50244 34204 50250
rect 34152 50186 34204 50192
rect 33784 50176 33836 50182
rect 33784 50118 33836 50124
rect 33968 50176 34020 50182
rect 33968 50118 34020 50124
rect 33692 29300 33744 29306
rect 33692 29242 33744 29248
rect 33600 28620 33652 28626
rect 33600 28562 33652 28568
rect 33416 23520 33468 23526
rect 33416 23462 33468 23468
rect 33428 18358 33456 23462
rect 33416 18352 33468 18358
rect 33416 18294 33468 18300
rect 33324 14884 33376 14890
rect 33324 14826 33376 14832
rect 33152 12838 33272 12866
rect 30840 11212 30892 11218
rect 30840 11154 30892 11160
rect 33048 11212 33100 11218
rect 33048 11154 33100 11160
rect 33138 10976 33194 10985
rect 32610 10908 32918 10917
rect 33138 10911 33194 10920
rect 32610 10906 32616 10908
rect 32672 10906 32696 10908
rect 32752 10906 32776 10908
rect 32832 10906 32856 10908
rect 32912 10906 32918 10908
rect 32672 10854 32674 10906
rect 32854 10854 32856 10906
rect 32610 10852 32616 10854
rect 32672 10852 32696 10854
rect 32752 10852 32776 10854
rect 32832 10852 32856 10854
rect 32912 10852 32918 10854
rect 32610 10843 32918 10852
rect 33152 10674 33180 10911
rect 33140 10668 33192 10674
rect 33140 10610 33192 10616
rect 31950 10364 32258 10373
rect 31950 10362 31956 10364
rect 32012 10362 32036 10364
rect 32092 10362 32116 10364
rect 32172 10362 32196 10364
rect 32252 10362 32258 10364
rect 32012 10310 32014 10362
rect 32194 10310 32196 10362
rect 31950 10308 31956 10310
rect 32012 10308 32036 10310
rect 32092 10308 32116 10310
rect 32172 10308 32196 10310
rect 32252 10308 32258 10310
rect 31950 10299 32258 10308
rect 32610 9820 32918 9829
rect 32610 9818 32616 9820
rect 32672 9818 32696 9820
rect 32752 9818 32776 9820
rect 32832 9818 32856 9820
rect 32912 9818 32918 9820
rect 32672 9766 32674 9818
rect 32854 9766 32856 9818
rect 32610 9764 32616 9766
rect 32672 9764 32696 9766
rect 32752 9764 32776 9766
rect 32832 9764 32856 9766
rect 32912 9764 32918 9766
rect 32610 9755 32918 9764
rect 31950 9276 32258 9285
rect 31950 9274 31956 9276
rect 32012 9274 32036 9276
rect 32092 9274 32116 9276
rect 32172 9274 32196 9276
rect 32252 9274 32258 9276
rect 32012 9222 32014 9274
rect 32194 9222 32196 9274
rect 31950 9220 31956 9222
rect 32012 9220 32036 9222
rect 32092 9220 32116 9222
rect 32172 9220 32196 9222
rect 32252 9220 32258 9222
rect 31950 9211 32258 9220
rect 33244 9178 33272 12838
rect 33796 10810 33824 50118
rect 33876 48136 33928 48142
rect 33876 48078 33928 48084
rect 33888 41070 33916 48078
rect 33876 41064 33928 41070
rect 33876 41006 33928 41012
rect 33980 17338 34008 50118
rect 34164 30734 34192 50186
rect 34624 46170 34652 55186
rect 34980 54528 35032 54534
rect 34980 54470 35032 54476
rect 34612 46164 34664 46170
rect 34612 46106 34664 46112
rect 34992 35698 35020 54470
rect 35164 47456 35216 47462
rect 35164 47398 35216 47404
rect 35176 45354 35204 47398
rect 35164 45348 35216 45354
rect 35164 45290 35216 45296
rect 34980 35692 35032 35698
rect 34980 35634 35032 35640
rect 34888 31816 34940 31822
rect 34888 31758 34940 31764
rect 34152 30728 34204 30734
rect 34152 30670 34204 30676
rect 34900 24206 34928 31758
rect 34888 24200 34940 24206
rect 34888 24142 34940 24148
rect 33968 17332 34020 17338
rect 33968 17274 34020 17280
rect 34900 13394 34928 24142
rect 34992 16590 35020 35634
rect 35452 35630 35480 58414
rect 36004 44946 36032 68682
rect 36084 62688 36136 62694
rect 36084 62630 36136 62636
rect 36096 53582 36124 62630
rect 36188 57526 36216 68818
rect 36544 68672 36596 68678
rect 36544 68614 36596 68620
rect 36636 68672 36688 68678
rect 36636 68614 36688 68620
rect 37372 68672 37424 68678
rect 37372 68614 37424 68620
rect 36556 64122 36584 68614
rect 36544 64116 36596 64122
rect 36544 64058 36596 64064
rect 36176 57520 36228 57526
rect 36176 57462 36228 57468
rect 36084 53576 36136 53582
rect 36084 53518 36136 53524
rect 35992 44940 36044 44946
rect 35992 44882 36044 44888
rect 35440 35624 35492 35630
rect 35440 35566 35492 35572
rect 35348 35488 35400 35494
rect 35348 35430 35400 35436
rect 35360 32230 35388 35430
rect 35452 34610 35480 35566
rect 35440 34604 35492 34610
rect 35440 34546 35492 34552
rect 35440 32360 35492 32366
rect 35440 32302 35492 32308
rect 35348 32224 35400 32230
rect 35348 32166 35400 32172
rect 35452 31890 35480 32302
rect 35440 31884 35492 31890
rect 35440 31826 35492 31832
rect 36188 22506 36216 57462
rect 36452 57452 36504 57458
rect 36452 57394 36504 57400
rect 36464 56778 36492 57394
rect 36452 56772 36504 56778
rect 36452 56714 36504 56720
rect 36360 52488 36412 52494
rect 36360 52430 36412 52436
rect 36176 22500 36228 22506
rect 36176 22442 36228 22448
rect 34980 16584 35032 16590
rect 34980 16526 35032 16532
rect 34888 13388 34940 13394
rect 34888 13330 34940 13336
rect 33784 10804 33836 10810
rect 33784 10746 33836 10752
rect 36372 10742 36400 52430
rect 36556 50182 36584 64058
rect 36544 50176 36596 50182
rect 36544 50118 36596 50124
rect 36556 49774 36584 50118
rect 36544 49768 36596 49774
rect 36544 49710 36596 49716
rect 36452 31884 36504 31890
rect 36452 31826 36504 31832
rect 36464 17882 36492 31826
rect 36544 31816 36596 31822
rect 36544 31758 36596 31764
rect 36452 17876 36504 17882
rect 36452 17818 36504 17824
rect 36464 13258 36492 17818
rect 36556 17542 36584 31758
rect 36648 26042 36676 68614
rect 36950 68028 37258 68037
rect 36950 68026 36956 68028
rect 37012 68026 37036 68028
rect 37092 68026 37116 68028
rect 37172 68026 37196 68028
rect 37252 68026 37258 68028
rect 37012 67974 37014 68026
rect 37194 67974 37196 68026
rect 36950 67972 36956 67974
rect 37012 67972 37036 67974
rect 37092 67972 37116 67974
rect 37172 67972 37196 67974
rect 37252 67972 37258 67974
rect 36950 67963 37258 67972
rect 36950 66940 37258 66949
rect 36950 66938 36956 66940
rect 37012 66938 37036 66940
rect 37092 66938 37116 66940
rect 37172 66938 37196 66940
rect 37252 66938 37258 66940
rect 37012 66886 37014 66938
rect 37194 66886 37196 66938
rect 36950 66884 36956 66886
rect 37012 66884 37036 66886
rect 37092 66884 37116 66886
rect 37172 66884 37196 66886
rect 37252 66884 37258 66886
rect 36950 66875 37258 66884
rect 36950 65852 37258 65861
rect 36950 65850 36956 65852
rect 37012 65850 37036 65852
rect 37092 65850 37116 65852
rect 37172 65850 37196 65852
rect 37252 65850 37258 65852
rect 37012 65798 37014 65850
rect 37194 65798 37196 65850
rect 36950 65796 36956 65798
rect 37012 65796 37036 65798
rect 37092 65796 37116 65798
rect 37172 65796 37196 65798
rect 37252 65796 37258 65798
rect 36950 65787 37258 65796
rect 36950 64764 37258 64773
rect 36950 64762 36956 64764
rect 37012 64762 37036 64764
rect 37092 64762 37116 64764
rect 37172 64762 37196 64764
rect 37252 64762 37258 64764
rect 37012 64710 37014 64762
rect 37194 64710 37196 64762
rect 36950 64708 36956 64710
rect 37012 64708 37036 64710
rect 37092 64708 37116 64710
rect 37172 64708 37196 64710
rect 37252 64708 37258 64710
rect 36950 64699 37258 64708
rect 36950 63676 37258 63685
rect 36950 63674 36956 63676
rect 37012 63674 37036 63676
rect 37092 63674 37116 63676
rect 37172 63674 37196 63676
rect 37252 63674 37258 63676
rect 37012 63622 37014 63674
rect 37194 63622 37196 63674
rect 36950 63620 36956 63622
rect 37012 63620 37036 63622
rect 37092 63620 37116 63622
rect 37172 63620 37196 63622
rect 37252 63620 37258 63622
rect 36950 63611 37258 63620
rect 36950 62588 37258 62597
rect 36950 62586 36956 62588
rect 37012 62586 37036 62588
rect 37092 62586 37116 62588
rect 37172 62586 37196 62588
rect 37252 62586 37258 62588
rect 37012 62534 37014 62586
rect 37194 62534 37196 62586
rect 36950 62532 36956 62534
rect 37012 62532 37036 62534
rect 37092 62532 37116 62534
rect 37172 62532 37196 62534
rect 37252 62532 37258 62534
rect 36950 62523 37258 62532
rect 36820 62280 36872 62286
rect 36820 62222 36872 62228
rect 36832 57798 36860 62222
rect 36950 61500 37258 61509
rect 36950 61498 36956 61500
rect 37012 61498 37036 61500
rect 37092 61498 37116 61500
rect 37172 61498 37196 61500
rect 37252 61498 37258 61500
rect 37012 61446 37014 61498
rect 37194 61446 37196 61498
rect 36950 61444 36956 61446
rect 37012 61444 37036 61446
rect 37092 61444 37116 61446
rect 37172 61444 37196 61446
rect 37252 61444 37258 61446
rect 36950 61435 37258 61444
rect 36950 60412 37258 60421
rect 36950 60410 36956 60412
rect 37012 60410 37036 60412
rect 37092 60410 37116 60412
rect 37172 60410 37196 60412
rect 37252 60410 37258 60412
rect 37012 60358 37014 60410
rect 37194 60358 37196 60410
rect 36950 60356 36956 60358
rect 37012 60356 37036 60358
rect 37092 60356 37116 60358
rect 37172 60356 37196 60358
rect 37252 60356 37258 60358
rect 36950 60347 37258 60356
rect 36950 59324 37258 59333
rect 36950 59322 36956 59324
rect 37012 59322 37036 59324
rect 37092 59322 37116 59324
rect 37172 59322 37196 59324
rect 37252 59322 37258 59324
rect 37012 59270 37014 59322
rect 37194 59270 37196 59322
rect 36950 59268 36956 59270
rect 37012 59268 37036 59270
rect 37092 59268 37116 59270
rect 37172 59268 37196 59270
rect 37252 59268 37258 59270
rect 36950 59259 37258 59268
rect 36950 58236 37258 58245
rect 36950 58234 36956 58236
rect 37012 58234 37036 58236
rect 37092 58234 37116 58236
rect 37172 58234 37196 58236
rect 37252 58234 37258 58236
rect 37012 58182 37014 58234
rect 37194 58182 37196 58234
rect 36950 58180 36956 58182
rect 37012 58180 37036 58182
rect 37092 58180 37116 58182
rect 37172 58180 37196 58182
rect 37252 58180 37258 58182
rect 36950 58171 37258 58180
rect 36820 57792 36872 57798
rect 36820 57734 36872 57740
rect 37280 57316 37332 57322
rect 37280 57258 37332 57264
rect 36950 57148 37258 57157
rect 36950 57146 36956 57148
rect 37012 57146 37036 57148
rect 37092 57146 37116 57148
rect 37172 57146 37196 57148
rect 37252 57146 37258 57148
rect 37012 57094 37014 57146
rect 37194 57094 37196 57146
rect 36950 57092 36956 57094
rect 37012 57092 37036 57094
rect 37092 57092 37116 57094
rect 37172 57092 37196 57094
rect 37252 57092 37258 57094
rect 36950 57083 37258 57092
rect 37292 56370 37320 57258
rect 37280 56364 37332 56370
rect 37280 56306 37332 56312
rect 36950 56060 37258 56069
rect 36950 56058 36956 56060
rect 37012 56058 37036 56060
rect 37092 56058 37116 56060
rect 37172 56058 37196 56060
rect 37252 56058 37258 56060
rect 37012 56006 37014 56058
rect 37194 56006 37196 56058
rect 36950 56004 36956 56006
rect 37012 56004 37036 56006
rect 37092 56004 37116 56006
rect 37172 56004 37196 56006
rect 37252 56004 37258 56006
rect 36950 55995 37258 56004
rect 36950 54972 37258 54981
rect 36950 54970 36956 54972
rect 37012 54970 37036 54972
rect 37092 54970 37116 54972
rect 37172 54970 37196 54972
rect 37252 54970 37258 54972
rect 37012 54918 37014 54970
rect 37194 54918 37196 54970
rect 36950 54916 36956 54918
rect 37012 54916 37036 54918
rect 37092 54916 37116 54918
rect 37172 54916 37196 54918
rect 37252 54916 37258 54918
rect 36950 54907 37258 54916
rect 36950 53884 37258 53893
rect 36950 53882 36956 53884
rect 37012 53882 37036 53884
rect 37092 53882 37116 53884
rect 37172 53882 37196 53884
rect 37252 53882 37258 53884
rect 37012 53830 37014 53882
rect 37194 53830 37196 53882
rect 36950 53828 36956 53830
rect 37012 53828 37036 53830
rect 37092 53828 37116 53830
rect 37172 53828 37196 53830
rect 37252 53828 37258 53830
rect 36950 53819 37258 53828
rect 36950 52796 37258 52805
rect 36950 52794 36956 52796
rect 37012 52794 37036 52796
rect 37092 52794 37116 52796
rect 37172 52794 37196 52796
rect 37252 52794 37258 52796
rect 37012 52742 37014 52794
rect 37194 52742 37196 52794
rect 36950 52740 36956 52742
rect 37012 52740 37036 52742
rect 37092 52740 37116 52742
rect 37172 52740 37196 52742
rect 37252 52740 37258 52742
rect 36950 52731 37258 52740
rect 36950 51708 37258 51717
rect 36950 51706 36956 51708
rect 37012 51706 37036 51708
rect 37092 51706 37116 51708
rect 37172 51706 37196 51708
rect 37252 51706 37258 51708
rect 37012 51654 37014 51706
rect 37194 51654 37196 51706
rect 36950 51652 36956 51654
rect 37012 51652 37036 51654
rect 37092 51652 37116 51654
rect 37172 51652 37196 51654
rect 37252 51652 37258 51654
rect 36950 51643 37258 51652
rect 36950 50620 37258 50629
rect 36950 50618 36956 50620
rect 37012 50618 37036 50620
rect 37092 50618 37116 50620
rect 37172 50618 37196 50620
rect 37252 50618 37258 50620
rect 37012 50566 37014 50618
rect 37194 50566 37196 50618
rect 36950 50564 36956 50566
rect 37012 50564 37036 50566
rect 37092 50564 37116 50566
rect 37172 50564 37196 50566
rect 37252 50564 37258 50566
rect 36950 50555 37258 50564
rect 36728 49768 36780 49774
rect 36728 49710 36780 49716
rect 36740 35222 36768 49710
rect 36950 49532 37258 49541
rect 36950 49530 36956 49532
rect 37012 49530 37036 49532
rect 37092 49530 37116 49532
rect 37172 49530 37196 49532
rect 37252 49530 37258 49532
rect 37012 49478 37014 49530
rect 37194 49478 37196 49530
rect 36950 49476 36956 49478
rect 37012 49476 37036 49478
rect 37092 49476 37116 49478
rect 37172 49476 37196 49478
rect 37252 49476 37258 49478
rect 36950 49467 37258 49476
rect 36950 48444 37258 48453
rect 36950 48442 36956 48444
rect 37012 48442 37036 48444
rect 37092 48442 37116 48444
rect 37172 48442 37196 48444
rect 37252 48442 37258 48444
rect 37012 48390 37014 48442
rect 37194 48390 37196 48442
rect 36950 48388 36956 48390
rect 37012 48388 37036 48390
rect 37092 48388 37116 48390
rect 37172 48388 37196 48390
rect 37252 48388 37258 48390
rect 36950 48379 37258 48388
rect 36950 47356 37258 47365
rect 36950 47354 36956 47356
rect 37012 47354 37036 47356
rect 37092 47354 37116 47356
rect 37172 47354 37196 47356
rect 37252 47354 37258 47356
rect 37012 47302 37014 47354
rect 37194 47302 37196 47354
rect 36950 47300 36956 47302
rect 37012 47300 37036 47302
rect 37092 47300 37116 47302
rect 37172 47300 37196 47302
rect 37252 47300 37258 47302
rect 36950 47291 37258 47300
rect 36950 46268 37258 46277
rect 36950 46266 36956 46268
rect 37012 46266 37036 46268
rect 37092 46266 37116 46268
rect 37172 46266 37196 46268
rect 37252 46266 37258 46268
rect 37012 46214 37014 46266
rect 37194 46214 37196 46266
rect 36950 46212 36956 46214
rect 37012 46212 37036 46214
rect 37092 46212 37116 46214
rect 37172 46212 37196 46214
rect 37252 46212 37258 46214
rect 36950 46203 37258 46212
rect 36950 45180 37258 45189
rect 36950 45178 36956 45180
rect 37012 45178 37036 45180
rect 37092 45178 37116 45180
rect 37172 45178 37196 45180
rect 37252 45178 37258 45180
rect 37012 45126 37014 45178
rect 37194 45126 37196 45178
rect 36950 45124 36956 45126
rect 37012 45124 37036 45126
rect 37092 45124 37116 45126
rect 37172 45124 37196 45126
rect 37252 45124 37258 45126
rect 36950 45115 37258 45124
rect 36950 44092 37258 44101
rect 36950 44090 36956 44092
rect 37012 44090 37036 44092
rect 37092 44090 37116 44092
rect 37172 44090 37196 44092
rect 37252 44090 37258 44092
rect 37012 44038 37014 44090
rect 37194 44038 37196 44090
rect 36950 44036 36956 44038
rect 37012 44036 37036 44038
rect 37092 44036 37116 44038
rect 37172 44036 37196 44038
rect 37252 44036 37258 44038
rect 36950 44027 37258 44036
rect 36950 43004 37258 43013
rect 36950 43002 36956 43004
rect 37012 43002 37036 43004
rect 37092 43002 37116 43004
rect 37172 43002 37196 43004
rect 37252 43002 37258 43004
rect 37012 42950 37014 43002
rect 37194 42950 37196 43002
rect 36950 42948 36956 42950
rect 37012 42948 37036 42950
rect 37092 42948 37116 42950
rect 37172 42948 37196 42950
rect 37252 42948 37258 42950
rect 36950 42939 37258 42948
rect 36950 41916 37258 41925
rect 36950 41914 36956 41916
rect 37012 41914 37036 41916
rect 37092 41914 37116 41916
rect 37172 41914 37196 41916
rect 37252 41914 37258 41916
rect 37012 41862 37014 41914
rect 37194 41862 37196 41914
rect 36950 41860 36956 41862
rect 37012 41860 37036 41862
rect 37092 41860 37116 41862
rect 37172 41860 37196 41862
rect 37252 41860 37258 41862
rect 36950 41851 37258 41860
rect 36820 41608 36872 41614
rect 36820 41550 36872 41556
rect 36728 35216 36780 35222
rect 36728 35158 36780 35164
rect 36832 32434 36860 41550
rect 37280 41540 37332 41546
rect 37280 41482 37332 41488
rect 36950 40828 37258 40837
rect 36950 40826 36956 40828
rect 37012 40826 37036 40828
rect 37092 40826 37116 40828
rect 37172 40826 37196 40828
rect 37252 40826 37258 40828
rect 37012 40774 37014 40826
rect 37194 40774 37196 40826
rect 36950 40772 36956 40774
rect 37012 40772 37036 40774
rect 37092 40772 37116 40774
rect 37172 40772 37196 40774
rect 37252 40772 37258 40774
rect 36950 40763 37258 40772
rect 36950 39740 37258 39749
rect 36950 39738 36956 39740
rect 37012 39738 37036 39740
rect 37092 39738 37116 39740
rect 37172 39738 37196 39740
rect 37252 39738 37258 39740
rect 37012 39686 37014 39738
rect 37194 39686 37196 39738
rect 36950 39684 36956 39686
rect 37012 39684 37036 39686
rect 37092 39684 37116 39686
rect 37172 39684 37196 39686
rect 37252 39684 37258 39686
rect 36950 39675 37258 39684
rect 36950 38652 37258 38661
rect 36950 38650 36956 38652
rect 37012 38650 37036 38652
rect 37092 38650 37116 38652
rect 37172 38650 37196 38652
rect 37252 38650 37258 38652
rect 37012 38598 37014 38650
rect 37194 38598 37196 38650
rect 36950 38596 36956 38598
rect 37012 38596 37036 38598
rect 37092 38596 37116 38598
rect 37172 38596 37196 38598
rect 37252 38596 37258 38598
rect 36950 38587 37258 38596
rect 37292 37670 37320 41482
rect 37280 37664 37332 37670
rect 37280 37606 37332 37612
rect 36950 37564 37258 37573
rect 36950 37562 36956 37564
rect 37012 37562 37036 37564
rect 37092 37562 37116 37564
rect 37172 37562 37196 37564
rect 37252 37562 37258 37564
rect 37012 37510 37014 37562
rect 37194 37510 37196 37562
rect 36950 37508 36956 37510
rect 37012 37508 37036 37510
rect 37092 37508 37116 37510
rect 37172 37508 37196 37510
rect 37252 37508 37258 37510
rect 36950 37499 37258 37508
rect 36950 36476 37258 36485
rect 36950 36474 36956 36476
rect 37012 36474 37036 36476
rect 37092 36474 37116 36476
rect 37172 36474 37196 36476
rect 37252 36474 37258 36476
rect 37012 36422 37014 36474
rect 37194 36422 37196 36474
rect 36950 36420 36956 36422
rect 37012 36420 37036 36422
rect 37092 36420 37116 36422
rect 37172 36420 37196 36422
rect 37252 36420 37258 36422
rect 36950 36411 37258 36420
rect 36950 35388 37258 35397
rect 36950 35386 36956 35388
rect 37012 35386 37036 35388
rect 37092 35386 37116 35388
rect 37172 35386 37196 35388
rect 37252 35386 37258 35388
rect 37012 35334 37014 35386
rect 37194 35334 37196 35386
rect 36950 35332 36956 35334
rect 37012 35332 37036 35334
rect 37092 35332 37116 35334
rect 37172 35332 37196 35334
rect 37252 35332 37258 35334
rect 36950 35323 37258 35332
rect 36950 34300 37258 34309
rect 36950 34298 36956 34300
rect 37012 34298 37036 34300
rect 37092 34298 37116 34300
rect 37172 34298 37196 34300
rect 37252 34298 37258 34300
rect 37012 34246 37014 34298
rect 37194 34246 37196 34298
rect 36950 34244 36956 34246
rect 37012 34244 37036 34246
rect 37092 34244 37116 34246
rect 37172 34244 37196 34246
rect 37252 34244 37258 34246
rect 36950 34235 37258 34244
rect 36950 33212 37258 33221
rect 36950 33210 36956 33212
rect 37012 33210 37036 33212
rect 37092 33210 37116 33212
rect 37172 33210 37196 33212
rect 37252 33210 37258 33212
rect 37012 33158 37014 33210
rect 37194 33158 37196 33210
rect 36950 33156 36956 33158
rect 37012 33156 37036 33158
rect 37092 33156 37116 33158
rect 37172 33156 37196 33158
rect 37252 33156 37258 33158
rect 36950 33147 37258 33156
rect 36820 32428 36872 32434
rect 36820 32370 36872 32376
rect 36950 32124 37258 32133
rect 36950 32122 36956 32124
rect 37012 32122 37036 32124
rect 37092 32122 37116 32124
rect 37172 32122 37196 32124
rect 37252 32122 37258 32124
rect 37012 32070 37014 32122
rect 37194 32070 37196 32122
rect 36950 32068 36956 32070
rect 37012 32068 37036 32070
rect 37092 32068 37116 32070
rect 37172 32068 37196 32070
rect 37252 32068 37258 32070
rect 36950 32059 37258 32068
rect 36950 31036 37258 31045
rect 36950 31034 36956 31036
rect 37012 31034 37036 31036
rect 37092 31034 37116 31036
rect 37172 31034 37196 31036
rect 37252 31034 37258 31036
rect 37012 30982 37014 31034
rect 37194 30982 37196 31034
rect 36950 30980 36956 30982
rect 37012 30980 37036 30982
rect 37092 30980 37116 30982
rect 37172 30980 37196 30982
rect 37252 30980 37258 30982
rect 36950 30971 37258 30980
rect 36950 29948 37258 29957
rect 36950 29946 36956 29948
rect 37012 29946 37036 29948
rect 37092 29946 37116 29948
rect 37172 29946 37196 29948
rect 37252 29946 37258 29948
rect 37012 29894 37014 29946
rect 37194 29894 37196 29946
rect 36950 29892 36956 29894
rect 37012 29892 37036 29894
rect 37092 29892 37116 29894
rect 37172 29892 37196 29894
rect 37252 29892 37258 29894
rect 36950 29883 37258 29892
rect 36950 28860 37258 28869
rect 36950 28858 36956 28860
rect 37012 28858 37036 28860
rect 37092 28858 37116 28860
rect 37172 28858 37196 28860
rect 37252 28858 37258 28860
rect 37012 28806 37014 28858
rect 37194 28806 37196 28858
rect 36950 28804 36956 28806
rect 37012 28804 37036 28806
rect 37092 28804 37116 28806
rect 37172 28804 37196 28806
rect 37252 28804 37258 28806
rect 36950 28795 37258 28804
rect 36950 27772 37258 27781
rect 36950 27770 36956 27772
rect 37012 27770 37036 27772
rect 37092 27770 37116 27772
rect 37172 27770 37196 27772
rect 37252 27770 37258 27772
rect 37012 27718 37014 27770
rect 37194 27718 37196 27770
rect 36950 27716 36956 27718
rect 37012 27716 37036 27718
rect 37092 27716 37116 27718
rect 37172 27716 37196 27718
rect 37252 27716 37258 27718
rect 36950 27707 37258 27716
rect 36950 26684 37258 26693
rect 36950 26682 36956 26684
rect 37012 26682 37036 26684
rect 37092 26682 37116 26684
rect 37172 26682 37196 26684
rect 37252 26682 37258 26684
rect 37012 26630 37014 26682
rect 37194 26630 37196 26682
rect 36950 26628 36956 26630
rect 37012 26628 37036 26630
rect 37092 26628 37116 26630
rect 37172 26628 37196 26630
rect 37252 26628 37258 26630
rect 36950 26619 37258 26628
rect 36636 26036 36688 26042
rect 36636 25978 36688 25984
rect 36950 25596 37258 25605
rect 36950 25594 36956 25596
rect 37012 25594 37036 25596
rect 37092 25594 37116 25596
rect 37172 25594 37196 25596
rect 37252 25594 37258 25596
rect 37012 25542 37014 25594
rect 37194 25542 37196 25594
rect 36950 25540 36956 25542
rect 37012 25540 37036 25542
rect 37092 25540 37116 25542
rect 37172 25540 37196 25542
rect 37252 25540 37258 25542
rect 36950 25531 37258 25540
rect 36950 24508 37258 24517
rect 36950 24506 36956 24508
rect 37012 24506 37036 24508
rect 37092 24506 37116 24508
rect 37172 24506 37196 24508
rect 37252 24506 37258 24508
rect 37012 24454 37014 24506
rect 37194 24454 37196 24506
rect 36950 24452 36956 24454
rect 37012 24452 37036 24454
rect 37092 24452 37116 24454
rect 37172 24452 37196 24454
rect 37252 24452 37258 24454
rect 36950 24443 37258 24452
rect 36950 23420 37258 23429
rect 36950 23418 36956 23420
rect 37012 23418 37036 23420
rect 37092 23418 37116 23420
rect 37172 23418 37196 23420
rect 37252 23418 37258 23420
rect 37012 23366 37014 23418
rect 37194 23366 37196 23418
rect 36950 23364 36956 23366
rect 37012 23364 37036 23366
rect 37092 23364 37116 23366
rect 37172 23364 37196 23366
rect 37252 23364 37258 23366
rect 36950 23355 37258 23364
rect 36950 22332 37258 22341
rect 36950 22330 36956 22332
rect 37012 22330 37036 22332
rect 37092 22330 37116 22332
rect 37172 22330 37196 22332
rect 37252 22330 37258 22332
rect 37012 22278 37014 22330
rect 37194 22278 37196 22330
rect 36950 22276 36956 22278
rect 37012 22276 37036 22278
rect 37092 22276 37116 22278
rect 37172 22276 37196 22278
rect 37252 22276 37258 22278
rect 36950 22267 37258 22276
rect 37384 21554 37412 68614
rect 37610 68572 37918 68581
rect 37610 68570 37616 68572
rect 37672 68570 37696 68572
rect 37752 68570 37776 68572
rect 37832 68570 37856 68572
rect 37912 68570 37918 68572
rect 37672 68518 37674 68570
rect 37854 68518 37856 68570
rect 37610 68516 37616 68518
rect 37672 68516 37696 68518
rect 37752 68516 37776 68518
rect 37832 68516 37856 68518
rect 37912 68516 37918 68518
rect 37610 68507 37918 68516
rect 37464 67788 37516 67794
rect 37464 67730 37516 67736
rect 37476 60042 37504 67730
rect 37610 67484 37918 67493
rect 37610 67482 37616 67484
rect 37672 67482 37696 67484
rect 37752 67482 37776 67484
rect 37832 67482 37856 67484
rect 37912 67482 37918 67484
rect 37672 67430 37674 67482
rect 37854 67430 37856 67482
rect 37610 67428 37616 67430
rect 37672 67428 37696 67430
rect 37752 67428 37776 67430
rect 37832 67428 37856 67430
rect 37912 67428 37918 67430
rect 37610 67419 37918 67428
rect 37610 66396 37918 66405
rect 37610 66394 37616 66396
rect 37672 66394 37696 66396
rect 37752 66394 37776 66396
rect 37832 66394 37856 66396
rect 37912 66394 37918 66396
rect 37672 66342 37674 66394
rect 37854 66342 37856 66394
rect 37610 66340 37616 66342
rect 37672 66340 37696 66342
rect 37752 66340 37776 66342
rect 37832 66340 37856 66342
rect 37912 66340 37918 66342
rect 37610 66331 37918 66340
rect 37610 65308 37918 65317
rect 37610 65306 37616 65308
rect 37672 65306 37696 65308
rect 37752 65306 37776 65308
rect 37832 65306 37856 65308
rect 37912 65306 37918 65308
rect 37672 65254 37674 65306
rect 37854 65254 37856 65306
rect 37610 65252 37616 65254
rect 37672 65252 37696 65254
rect 37752 65252 37776 65254
rect 37832 65252 37856 65254
rect 37912 65252 37918 65254
rect 37610 65243 37918 65252
rect 37610 64220 37918 64229
rect 37610 64218 37616 64220
rect 37672 64218 37696 64220
rect 37752 64218 37776 64220
rect 37832 64218 37856 64220
rect 37912 64218 37918 64220
rect 37672 64166 37674 64218
rect 37854 64166 37856 64218
rect 37610 64164 37616 64166
rect 37672 64164 37696 64166
rect 37752 64164 37776 64166
rect 37832 64164 37856 64166
rect 37912 64164 37918 64166
rect 37610 64155 37918 64164
rect 37610 63132 37918 63141
rect 37610 63130 37616 63132
rect 37672 63130 37696 63132
rect 37752 63130 37776 63132
rect 37832 63130 37856 63132
rect 37912 63130 37918 63132
rect 37672 63078 37674 63130
rect 37854 63078 37856 63130
rect 37610 63076 37616 63078
rect 37672 63076 37696 63078
rect 37752 63076 37776 63078
rect 37832 63076 37856 63078
rect 37912 63076 37918 63078
rect 37610 63067 37918 63076
rect 37610 62044 37918 62053
rect 37610 62042 37616 62044
rect 37672 62042 37696 62044
rect 37752 62042 37776 62044
rect 37832 62042 37856 62044
rect 37912 62042 37918 62044
rect 37672 61990 37674 62042
rect 37854 61990 37856 62042
rect 37610 61988 37616 61990
rect 37672 61988 37696 61990
rect 37752 61988 37776 61990
rect 37832 61988 37856 61990
rect 37912 61988 37918 61990
rect 37610 61979 37918 61988
rect 37610 60956 37918 60965
rect 37610 60954 37616 60956
rect 37672 60954 37696 60956
rect 37752 60954 37776 60956
rect 37832 60954 37856 60956
rect 37912 60954 37918 60956
rect 37672 60902 37674 60954
rect 37854 60902 37856 60954
rect 37610 60900 37616 60902
rect 37672 60900 37696 60902
rect 37752 60900 37776 60902
rect 37832 60900 37856 60902
rect 37912 60900 37918 60902
rect 37610 60891 37918 60900
rect 38476 60308 38528 60314
rect 38476 60250 38528 60256
rect 37464 60036 37516 60042
rect 37464 59978 37516 59984
rect 38200 60036 38252 60042
rect 38200 59978 38252 59984
rect 37610 59868 37918 59877
rect 37610 59866 37616 59868
rect 37672 59866 37696 59868
rect 37752 59866 37776 59868
rect 37832 59866 37856 59868
rect 37912 59866 37918 59868
rect 37672 59814 37674 59866
rect 37854 59814 37856 59866
rect 37610 59812 37616 59814
rect 37672 59812 37696 59814
rect 37752 59812 37776 59814
rect 37832 59812 37856 59814
rect 37912 59812 37918 59814
rect 37610 59803 37918 59812
rect 37610 58780 37918 58789
rect 37610 58778 37616 58780
rect 37672 58778 37696 58780
rect 37752 58778 37776 58780
rect 37832 58778 37856 58780
rect 37912 58778 37918 58780
rect 37672 58726 37674 58778
rect 37854 58726 37856 58778
rect 37610 58724 37616 58726
rect 37672 58724 37696 58726
rect 37752 58724 37776 58726
rect 37832 58724 37856 58726
rect 37912 58724 37918 58726
rect 37610 58715 37918 58724
rect 37610 57692 37918 57701
rect 37610 57690 37616 57692
rect 37672 57690 37696 57692
rect 37752 57690 37776 57692
rect 37832 57690 37856 57692
rect 37912 57690 37918 57692
rect 37672 57638 37674 57690
rect 37854 57638 37856 57690
rect 37610 57636 37616 57638
rect 37672 57636 37696 57638
rect 37752 57636 37776 57638
rect 37832 57636 37856 57638
rect 37912 57636 37918 57638
rect 37610 57627 37918 57636
rect 37610 56604 37918 56613
rect 37610 56602 37616 56604
rect 37672 56602 37696 56604
rect 37752 56602 37776 56604
rect 37832 56602 37856 56604
rect 37912 56602 37918 56604
rect 37672 56550 37674 56602
rect 37854 56550 37856 56602
rect 37610 56548 37616 56550
rect 37672 56548 37696 56550
rect 37752 56548 37776 56550
rect 37832 56548 37856 56550
rect 37912 56548 37918 56550
rect 37610 56539 37918 56548
rect 37464 56432 37516 56438
rect 37464 56374 37516 56380
rect 37476 53514 37504 56374
rect 38016 56296 38068 56302
rect 38016 56238 38068 56244
rect 38108 56296 38160 56302
rect 38108 56238 38160 56244
rect 37610 55516 37918 55525
rect 37610 55514 37616 55516
rect 37672 55514 37696 55516
rect 37752 55514 37776 55516
rect 37832 55514 37856 55516
rect 37912 55514 37918 55516
rect 37672 55462 37674 55514
rect 37854 55462 37856 55514
rect 37610 55460 37616 55462
rect 37672 55460 37696 55462
rect 37752 55460 37776 55462
rect 37832 55460 37856 55462
rect 37912 55460 37918 55462
rect 37610 55451 37918 55460
rect 37610 54428 37918 54437
rect 37610 54426 37616 54428
rect 37672 54426 37696 54428
rect 37752 54426 37776 54428
rect 37832 54426 37856 54428
rect 37912 54426 37918 54428
rect 37672 54374 37674 54426
rect 37854 54374 37856 54426
rect 37610 54372 37616 54374
rect 37672 54372 37696 54374
rect 37752 54372 37776 54374
rect 37832 54372 37856 54374
rect 37912 54372 37918 54374
rect 37610 54363 37918 54372
rect 37464 53508 37516 53514
rect 37464 53450 37516 53456
rect 37476 50386 37504 53450
rect 37610 53340 37918 53349
rect 37610 53338 37616 53340
rect 37672 53338 37696 53340
rect 37752 53338 37776 53340
rect 37832 53338 37856 53340
rect 37912 53338 37918 53340
rect 37672 53286 37674 53338
rect 37854 53286 37856 53338
rect 37610 53284 37616 53286
rect 37672 53284 37696 53286
rect 37752 53284 37776 53286
rect 37832 53284 37856 53286
rect 37912 53284 37918 53286
rect 37610 53275 37918 53284
rect 37610 52252 37918 52261
rect 37610 52250 37616 52252
rect 37672 52250 37696 52252
rect 37752 52250 37776 52252
rect 37832 52250 37856 52252
rect 37912 52250 37918 52252
rect 37672 52198 37674 52250
rect 37854 52198 37856 52250
rect 37610 52196 37616 52198
rect 37672 52196 37696 52198
rect 37752 52196 37776 52198
rect 37832 52196 37856 52198
rect 37912 52196 37918 52198
rect 37610 52187 37918 52196
rect 37610 51164 37918 51173
rect 37610 51162 37616 51164
rect 37672 51162 37696 51164
rect 37752 51162 37776 51164
rect 37832 51162 37856 51164
rect 37912 51162 37918 51164
rect 37672 51110 37674 51162
rect 37854 51110 37856 51162
rect 37610 51108 37616 51110
rect 37672 51108 37696 51110
rect 37752 51108 37776 51110
rect 37832 51108 37856 51110
rect 37912 51108 37918 51110
rect 37610 51099 37918 51108
rect 37464 50380 37516 50386
rect 37464 50322 37516 50328
rect 37610 50076 37918 50085
rect 37610 50074 37616 50076
rect 37672 50074 37696 50076
rect 37752 50074 37776 50076
rect 37832 50074 37856 50076
rect 37912 50074 37918 50076
rect 37672 50022 37674 50074
rect 37854 50022 37856 50074
rect 37610 50020 37616 50022
rect 37672 50020 37696 50022
rect 37752 50020 37776 50022
rect 37832 50020 37856 50022
rect 37912 50020 37918 50022
rect 37610 50011 37918 50020
rect 37610 48988 37918 48997
rect 37610 48986 37616 48988
rect 37672 48986 37696 48988
rect 37752 48986 37776 48988
rect 37832 48986 37856 48988
rect 37912 48986 37918 48988
rect 37672 48934 37674 48986
rect 37854 48934 37856 48986
rect 37610 48932 37616 48934
rect 37672 48932 37696 48934
rect 37752 48932 37776 48934
rect 37832 48932 37856 48934
rect 37912 48932 37918 48934
rect 37610 48923 37918 48932
rect 37610 47900 37918 47909
rect 37610 47898 37616 47900
rect 37672 47898 37696 47900
rect 37752 47898 37776 47900
rect 37832 47898 37856 47900
rect 37912 47898 37918 47900
rect 37672 47846 37674 47898
rect 37854 47846 37856 47898
rect 37610 47844 37616 47846
rect 37672 47844 37696 47846
rect 37752 47844 37776 47846
rect 37832 47844 37856 47846
rect 37912 47844 37918 47846
rect 37610 47835 37918 47844
rect 37610 46812 37918 46821
rect 37610 46810 37616 46812
rect 37672 46810 37696 46812
rect 37752 46810 37776 46812
rect 37832 46810 37856 46812
rect 37912 46810 37918 46812
rect 37672 46758 37674 46810
rect 37854 46758 37856 46810
rect 37610 46756 37616 46758
rect 37672 46756 37696 46758
rect 37752 46756 37776 46758
rect 37832 46756 37856 46758
rect 37912 46756 37918 46758
rect 37610 46747 37918 46756
rect 37610 45724 37918 45733
rect 37610 45722 37616 45724
rect 37672 45722 37696 45724
rect 37752 45722 37776 45724
rect 37832 45722 37856 45724
rect 37912 45722 37918 45724
rect 37672 45670 37674 45722
rect 37854 45670 37856 45722
rect 37610 45668 37616 45670
rect 37672 45668 37696 45670
rect 37752 45668 37776 45670
rect 37832 45668 37856 45670
rect 37912 45668 37918 45670
rect 37610 45659 37918 45668
rect 37610 44636 37918 44645
rect 37610 44634 37616 44636
rect 37672 44634 37696 44636
rect 37752 44634 37776 44636
rect 37832 44634 37856 44636
rect 37912 44634 37918 44636
rect 37672 44582 37674 44634
rect 37854 44582 37856 44634
rect 37610 44580 37616 44582
rect 37672 44580 37696 44582
rect 37752 44580 37776 44582
rect 37832 44580 37856 44582
rect 37912 44580 37918 44582
rect 37610 44571 37918 44580
rect 37610 43548 37918 43557
rect 37610 43546 37616 43548
rect 37672 43546 37696 43548
rect 37752 43546 37776 43548
rect 37832 43546 37856 43548
rect 37912 43546 37918 43548
rect 37672 43494 37674 43546
rect 37854 43494 37856 43546
rect 37610 43492 37616 43494
rect 37672 43492 37696 43494
rect 37752 43492 37776 43494
rect 37832 43492 37856 43494
rect 37912 43492 37918 43494
rect 37610 43483 37918 43492
rect 37610 42460 37918 42469
rect 37610 42458 37616 42460
rect 37672 42458 37696 42460
rect 37752 42458 37776 42460
rect 37832 42458 37856 42460
rect 37912 42458 37918 42460
rect 37672 42406 37674 42458
rect 37854 42406 37856 42458
rect 37610 42404 37616 42406
rect 37672 42404 37696 42406
rect 37752 42404 37776 42406
rect 37832 42404 37856 42406
rect 37912 42404 37918 42406
rect 37610 42395 37918 42404
rect 37610 41372 37918 41381
rect 37610 41370 37616 41372
rect 37672 41370 37696 41372
rect 37752 41370 37776 41372
rect 37832 41370 37856 41372
rect 37912 41370 37918 41372
rect 37672 41318 37674 41370
rect 37854 41318 37856 41370
rect 37610 41316 37616 41318
rect 37672 41316 37696 41318
rect 37752 41316 37776 41318
rect 37832 41316 37856 41318
rect 37912 41316 37918 41318
rect 37610 41307 37918 41316
rect 37610 40284 37918 40293
rect 37610 40282 37616 40284
rect 37672 40282 37696 40284
rect 37752 40282 37776 40284
rect 37832 40282 37856 40284
rect 37912 40282 37918 40284
rect 37672 40230 37674 40282
rect 37854 40230 37856 40282
rect 37610 40228 37616 40230
rect 37672 40228 37696 40230
rect 37752 40228 37776 40230
rect 37832 40228 37856 40230
rect 37912 40228 37918 40230
rect 37610 40219 37918 40228
rect 37610 39196 37918 39205
rect 37610 39194 37616 39196
rect 37672 39194 37696 39196
rect 37752 39194 37776 39196
rect 37832 39194 37856 39196
rect 37912 39194 37918 39196
rect 37672 39142 37674 39194
rect 37854 39142 37856 39194
rect 37610 39140 37616 39142
rect 37672 39140 37696 39142
rect 37752 39140 37776 39142
rect 37832 39140 37856 39142
rect 37912 39140 37918 39142
rect 37610 39131 37918 39140
rect 37610 38108 37918 38117
rect 37610 38106 37616 38108
rect 37672 38106 37696 38108
rect 37752 38106 37776 38108
rect 37832 38106 37856 38108
rect 37912 38106 37918 38108
rect 37672 38054 37674 38106
rect 37854 38054 37856 38106
rect 37610 38052 37616 38054
rect 37672 38052 37696 38054
rect 37752 38052 37776 38054
rect 37832 38052 37856 38054
rect 37912 38052 37918 38054
rect 37610 38043 37918 38052
rect 37610 37020 37918 37029
rect 37610 37018 37616 37020
rect 37672 37018 37696 37020
rect 37752 37018 37776 37020
rect 37832 37018 37856 37020
rect 37912 37018 37918 37020
rect 37672 36966 37674 37018
rect 37854 36966 37856 37018
rect 37610 36964 37616 36966
rect 37672 36964 37696 36966
rect 37752 36964 37776 36966
rect 37832 36964 37856 36966
rect 37912 36964 37918 36966
rect 37610 36955 37918 36964
rect 37610 35932 37918 35941
rect 37610 35930 37616 35932
rect 37672 35930 37696 35932
rect 37752 35930 37776 35932
rect 37832 35930 37856 35932
rect 37912 35930 37918 35932
rect 37672 35878 37674 35930
rect 37854 35878 37856 35930
rect 37610 35876 37616 35878
rect 37672 35876 37696 35878
rect 37752 35876 37776 35878
rect 37832 35876 37856 35878
rect 37912 35876 37918 35878
rect 37610 35867 37918 35876
rect 37610 34844 37918 34853
rect 37610 34842 37616 34844
rect 37672 34842 37696 34844
rect 37752 34842 37776 34844
rect 37832 34842 37856 34844
rect 37912 34842 37918 34844
rect 37672 34790 37674 34842
rect 37854 34790 37856 34842
rect 37610 34788 37616 34790
rect 37672 34788 37696 34790
rect 37752 34788 37776 34790
rect 37832 34788 37856 34790
rect 37912 34788 37918 34790
rect 37610 34779 37918 34788
rect 37610 33756 37918 33765
rect 37610 33754 37616 33756
rect 37672 33754 37696 33756
rect 37752 33754 37776 33756
rect 37832 33754 37856 33756
rect 37912 33754 37918 33756
rect 37672 33702 37674 33754
rect 37854 33702 37856 33754
rect 37610 33700 37616 33702
rect 37672 33700 37696 33702
rect 37752 33700 37776 33702
rect 37832 33700 37856 33702
rect 37912 33700 37918 33702
rect 37610 33691 37918 33700
rect 37610 32668 37918 32677
rect 37610 32666 37616 32668
rect 37672 32666 37696 32668
rect 37752 32666 37776 32668
rect 37832 32666 37856 32668
rect 37912 32666 37918 32668
rect 37672 32614 37674 32666
rect 37854 32614 37856 32666
rect 37610 32612 37616 32614
rect 37672 32612 37696 32614
rect 37752 32612 37776 32614
rect 37832 32612 37856 32614
rect 37912 32612 37918 32614
rect 37610 32603 37918 32612
rect 37610 31580 37918 31589
rect 37610 31578 37616 31580
rect 37672 31578 37696 31580
rect 37752 31578 37776 31580
rect 37832 31578 37856 31580
rect 37912 31578 37918 31580
rect 37672 31526 37674 31578
rect 37854 31526 37856 31578
rect 37610 31524 37616 31526
rect 37672 31524 37696 31526
rect 37752 31524 37776 31526
rect 37832 31524 37856 31526
rect 37912 31524 37918 31526
rect 37610 31515 37918 31524
rect 37610 30492 37918 30501
rect 37610 30490 37616 30492
rect 37672 30490 37696 30492
rect 37752 30490 37776 30492
rect 37832 30490 37856 30492
rect 37912 30490 37918 30492
rect 37672 30438 37674 30490
rect 37854 30438 37856 30490
rect 37610 30436 37616 30438
rect 37672 30436 37696 30438
rect 37752 30436 37776 30438
rect 37832 30436 37856 30438
rect 37912 30436 37918 30438
rect 37610 30427 37918 30436
rect 37610 29404 37918 29413
rect 37610 29402 37616 29404
rect 37672 29402 37696 29404
rect 37752 29402 37776 29404
rect 37832 29402 37856 29404
rect 37912 29402 37918 29404
rect 37672 29350 37674 29402
rect 37854 29350 37856 29402
rect 37610 29348 37616 29350
rect 37672 29348 37696 29350
rect 37752 29348 37776 29350
rect 37832 29348 37856 29350
rect 37912 29348 37918 29350
rect 37610 29339 37918 29348
rect 37610 28316 37918 28325
rect 37610 28314 37616 28316
rect 37672 28314 37696 28316
rect 37752 28314 37776 28316
rect 37832 28314 37856 28316
rect 37912 28314 37918 28316
rect 37672 28262 37674 28314
rect 37854 28262 37856 28314
rect 37610 28260 37616 28262
rect 37672 28260 37696 28262
rect 37752 28260 37776 28262
rect 37832 28260 37856 28262
rect 37912 28260 37918 28262
rect 37610 28251 37918 28260
rect 38028 27334 38056 56238
rect 38120 55894 38148 56238
rect 38108 55888 38160 55894
rect 38108 55830 38160 55836
rect 38120 51074 38148 55830
rect 38212 52426 38240 59978
rect 38292 59968 38344 59974
rect 38292 59910 38344 59916
rect 38304 53786 38332 59910
rect 38292 53780 38344 53786
rect 38292 53722 38344 53728
rect 38200 52420 38252 52426
rect 38200 52362 38252 52368
rect 38120 51046 38240 51074
rect 38108 47252 38160 47258
rect 38108 47194 38160 47200
rect 38120 32774 38148 47194
rect 38212 47054 38240 51046
rect 38384 50380 38436 50386
rect 38384 50322 38436 50328
rect 38200 47048 38252 47054
rect 38200 46990 38252 46996
rect 38108 32768 38160 32774
rect 38108 32710 38160 32716
rect 38016 27328 38068 27334
rect 38016 27270 38068 27276
rect 37610 27228 37918 27237
rect 37610 27226 37616 27228
rect 37672 27226 37696 27228
rect 37752 27226 37776 27228
rect 37832 27226 37856 27228
rect 37912 27226 37918 27228
rect 37672 27174 37674 27226
rect 37854 27174 37856 27226
rect 37610 27172 37616 27174
rect 37672 27172 37696 27174
rect 37752 27172 37776 27174
rect 37832 27172 37856 27174
rect 37912 27172 37918 27174
rect 37610 27163 37918 27172
rect 37610 26140 37918 26149
rect 37610 26138 37616 26140
rect 37672 26138 37696 26140
rect 37752 26138 37776 26140
rect 37832 26138 37856 26140
rect 37912 26138 37918 26140
rect 37672 26086 37674 26138
rect 37854 26086 37856 26138
rect 37610 26084 37616 26086
rect 37672 26084 37696 26086
rect 37752 26084 37776 26086
rect 37832 26084 37856 26086
rect 37912 26084 37918 26086
rect 37610 26075 37918 26084
rect 37610 25052 37918 25061
rect 37610 25050 37616 25052
rect 37672 25050 37696 25052
rect 37752 25050 37776 25052
rect 37832 25050 37856 25052
rect 37912 25050 37918 25052
rect 37672 24998 37674 25050
rect 37854 24998 37856 25050
rect 37610 24996 37616 24998
rect 37672 24996 37696 24998
rect 37752 24996 37776 24998
rect 37832 24996 37856 24998
rect 37912 24996 37918 24998
rect 37610 24987 37918 24996
rect 37610 23964 37918 23973
rect 37610 23962 37616 23964
rect 37672 23962 37696 23964
rect 37752 23962 37776 23964
rect 37832 23962 37856 23964
rect 37912 23962 37918 23964
rect 37672 23910 37674 23962
rect 37854 23910 37856 23962
rect 37610 23908 37616 23910
rect 37672 23908 37696 23910
rect 37752 23908 37776 23910
rect 37832 23908 37856 23910
rect 37912 23908 37918 23910
rect 37610 23899 37918 23908
rect 37610 22876 37918 22885
rect 37610 22874 37616 22876
rect 37672 22874 37696 22876
rect 37752 22874 37776 22876
rect 37832 22874 37856 22876
rect 37912 22874 37918 22876
rect 37672 22822 37674 22874
rect 37854 22822 37856 22874
rect 37610 22820 37616 22822
rect 37672 22820 37696 22822
rect 37752 22820 37776 22822
rect 37832 22820 37856 22822
rect 37912 22820 37918 22822
rect 37610 22811 37918 22820
rect 37610 21788 37918 21797
rect 37610 21786 37616 21788
rect 37672 21786 37696 21788
rect 37752 21786 37776 21788
rect 37832 21786 37856 21788
rect 37912 21786 37918 21788
rect 37672 21734 37674 21786
rect 37854 21734 37856 21786
rect 37610 21732 37616 21734
rect 37672 21732 37696 21734
rect 37752 21732 37776 21734
rect 37832 21732 37856 21734
rect 37912 21732 37918 21734
rect 37610 21723 37918 21732
rect 37372 21548 37424 21554
rect 37372 21490 37424 21496
rect 36636 21480 36688 21486
rect 36636 21422 36688 21428
rect 36648 18426 36676 21422
rect 36950 21244 37258 21253
rect 36950 21242 36956 21244
rect 37012 21242 37036 21244
rect 37092 21242 37116 21244
rect 37172 21242 37196 21244
rect 37252 21242 37258 21244
rect 37012 21190 37014 21242
rect 37194 21190 37196 21242
rect 36950 21188 36956 21190
rect 37012 21188 37036 21190
rect 37092 21188 37116 21190
rect 37172 21188 37196 21190
rect 37252 21188 37258 21190
rect 36950 21179 37258 21188
rect 37610 20700 37918 20709
rect 37610 20698 37616 20700
rect 37672 20698 37696 20700
rect 37752 20698 37776 20700
rect 37832 20698 37856 20700
rect 37912 20698 37918 20700
rect 37672 20646 37674 20698
rect 37854 20646 37856 20698
rect 37610 20644 37616 20646
rect 37672 20644 37696 20646
rect 37752 20644 37776 20646
rect 37832 20644 37856 20646
rect 37912 20644 37918 20646
rect 37610 20635 37918 20644
rect 36950 20156 37258 20165
rect 36950 20154 36956 20156
rect 37012 20154 37036 20156
rect 37092 20154 37116 20156
rect 37172 20154 37196 20156
rect 37252 20154 37258 20156
rect 37012 20102 37014 20154
rect 37194 20102 37196 20154
rect 36950 20100 36956 20102
rect 37012 20100 37036 20102
rect 37092 20100 37116 20102
rect 37172 20100 37196 20102
rect 37252 20100 37258 20102
rect 36950 20091 37258 20100
rect 37610 19612 37918 19621
rect 37610 19610 37616 19612
rect 37672 19610 37696 19612
rect 37752 19610 37776 19612
rect 37832 19610 37856 19612
rect 37912 19610 37918 19612
rect 37672 19558 37674 19610
rect 37854 19558 37856 19610
rect 37610 19556 37616 19558
rect 37672 19556 37696 19558
rect 37752 19556 37776 19558
rect 37832 19556 37856 19558
rect 37912 19556 37918 19558
rect 37610 19547 37918 19556
rect 36950 19068 37258 19077
rect 36950 19066 36956 19068
rect 37012 19066 37036 19068
rect 37092 19066 37116 19068
rect 37172 19066 37196 19068
rect 37252 19066 37258 19068
rect 37012 19014 37014 19066
rect 37194 19014 37196 19066
rect 36950 19012 36956 19014
rect 37012 19012 37036 19014
rect 37092 19012 37116 19014
rect 37172 19012 37196 19014
rect 37252 19012 37258 19014
rect 36950 19003 37258 19012
rect 37610 18524 37918 18533
rect 37610 18522 37616 18524
rect 37672 18522 37696 18524
rect 37752 18522 37776 18524
rect 37832 18522 37856 18524
rect 37912 18522 37918 18524
rect 37672 18470 37674 18522
rect 37854 18470 37856 18522
rect 37610 18468 37616 18470
rect 37672 18468 37696 18470
rect 37752 18468 37776 18470
rect 37832 18468 37856 18470
rect 37912 18468 37918 18470
rect 37610 18459 37918 18468
rect 36636 18420 36688 18426
rect 36636 18362 36688 18368
rect 36544 17536 36596 17542
rect 36544 17478 36596 17484
rect 36452 13252 36504 13258
rect 36452 13194 36504 13200
rect 36360 10736 36412 10742
rect 36360 10678 36412 10684
rect 36464 10674 36492 13194
rect 36452 10668 36504 10674
rect 36452 10610 36504 10616
rect 33232 9172 33284 9178
rect 33232 9114 33284 9120
rect 32610 8732 32918 8741
rect 32610 8730 32616 8732
rect 32672 8730 32696 8732
rect 32752 8730 32776 8732
rect 32832 8730 32856 8732
rect 32912 8730 32918 8732
rect 32672 8678 32674 8730
rect 32854 8678 32856 8730
rect 32610 8676 32616 8678
rect 32672 8676 32696 8678
rect 32752 8676 32776 8678
rect 32832 8676 32856 8678
rect 32912 8676 32918 8678
rect 32610 8667 32918 8676
rect 31950 8188 32258 8197
rect 31950 8186 31956 8188
rect 32012 8186 32036 8188
rect 32092 8186 32116 8188
rect 32172 8186 32196 8188
rect 32252 8186 32258 8188
rect 32012 8134 32014 8186
rect 32194 8134 32196 8186
rect 31950 8132 31956 8134
rect 32012 8132 32036 8134
rect 32092 8132 32116 8134
rect 32172 8132 32196 8134
rect 32252 8132 32258 8134
rect 31950 8123 32258 8132
rect 32610 7644 32918 7653
rect 32610 7642 32616 7644
rect 32672 7642 32696 7644
rect 32752 7642 32776 7644
rect 32832 7642 32856 7644
rect 32912 7642 32918 7644
rect 32672 7590 32674 7642
rect 32854 7590 32856 7642
rect 32610 7588 32616 7590
rect 32672 7588 32696 7590
rect 32752 7588 32776 7590
rect 32832 7588 32856 7590
rect 32912 7588 32918 7590
rect 32610 7579 32918 7588
rect 31950 7100 32258 7109
rect 31950 7098 31956 7100
rect 32012 7098 32036 7100
rect 32092 7098 32116 7100
rect 32172 7098 32196 7100
rect 32252 7098 32258 7100
rect 32012 7046 32014 7098
rect 32194 7046 32196 7098
rect 31950 7044 31956 7046
rect 32012 7044 32036 7046
rect 32092 7044 32116 7046
rect 32172 7044 32196 7046
rect 32252 7044 32258 7046
rect 31950 7035 32258 7044
rect 32610 6556 32918 6565
rect 32610 6554 32616 6556
rect 32672 6554 32696 6556
rect 32752 6554 32776 6556
rect 32832 6554 32856 6556
rect 32912 6554 32918 6556
rect 32672 6502 32674 6554
rect 32854 6502 32856 6554
rect 32610 6500 32616 6502
rect 32672 6500 32696 6502
rect 32752 6500 32776 6502
rect 32832 6500 32856 6502
rect 32912 6500 32918 6502
rect 32610 6491 32918 6500
rect 31950 6012 32258 6021
rect 31950 6010 31956 6012
rect 32012 6010 32036 6012
rect 32092 6010 32116 6012
rect 32172 6010 32196 6012
rect 32252 6010 32258 6012
rect 32012 5958 32014 6010
rect 32194 5958 32196 6010
rect 31950 5956 31956 5958
rect 32012 5956 32036 5958
rect 32092 5956 32116 5958
rect 32172 5956 32196 5958
rect 32252 5956 32258 5958
rect 31950 5947 32258 5956
rect 32610 5468 32918 5477
rect 32610 5466 32616 5468
rect 32672 5466 32696 5468
rect 32752 5466 32776 5468
rect 32832 5466 32856 5468
rect 32912 5466 32918 5468
rect 32672 5414 32674 5466
rect 32854 5414 32856 5466
rect 32610 5412 32616 5414
rect 32672 5412 32696 5414
rect 32752 5412 32776 5414
rect 32832 5412 32856 5414
rect 32912 5412 32918 5414
rect 32610 5403 32918 5412
rect 31950 4924 32258 4933
rect 31950 4922 31956 4924
rect 32012 4922 32036 4924
rect 32092 4922 32116 4924
rect 32172 4922 32196 4924
rect 32252 4922 32258 4924
rect 32012 4870 32014 4922
rect 32194 4870 32196 4922
rect 31950 4868 31956 4870
rect 32012 4868 32036 4870
rect 32092 4868 32116 4870
rect 32172 4868 32196 4870
rect 32252 4868 32258 4870
rect 31950 4859 32258 4868
rect 32610 4380 32918 4389
rect 32610 4378 32616 4380
rect 32672 4378 32696 4380
rect 32752 4378 32776 4380
rect 32832 4378 32856 4380
rect 32912 4378 32918 4380
rect 32672 4326 32674 4378
rect 32854 4326 32856 4378
rect 32610 4324 32616 4326
rect 32672 4324 32696 4326
rect 32752 4324 32776 4326
rect 32832 4324 32856 4326
rect 32912 4324 32918 4326
rect 32610 4315 32918 4324
rect 31950 3836 32258 3845
rect 31950 3834 31956 3836
rect 32012 3834 32036 3836
rect 32092 3834 32116 3836
rect 32172 3834 32196 3836
rect 32252 3834 32258 3836
rect 32012 3782 32014 3834
rect 32194 3782 32196 3834
rect 31950 3780 31956 3782
rect 32012 3780 32036 3782
rect 32092 3780 32116 3782
rect 32172 3780 32196 3782
rect 32252 3780 32258 3782
rect 31950 3771 32258 3780
rect 29460 3732 29512 3738
rect 29460 3674 29512 3680
rect 32610 3292 32918 3301
rect 32610 3290 32616 3292
rect 32672 3290 32696 3292
rect 32752 3290 32776 3292
rect 32832 3290 32856 3292
rect 32912 3290 32918 3292
rect 32672 3238 32674 3290
rect 32854 3238 32856 3290
rect 32610 3236 32616 3238
rect 32672 3236 32696 3238
rect 32752 3236 32776 3238
rect 32832 3236 32856 3238
rect 32912 3236 32918 3238
rect 32610 3227 32918 3236
rect 21824 3052 21876 3058
rect 21824 2994 21876 3000
rect 29184 3052 29236 3058
rect 29184 2994 29236 3000
rect 21640 2848 21692 2854
rect 21640 2790 21692 2796
rect 21950 2748 22258 2757
rect 21950 2746 21956 2748
rect 22012 2746 22036 2748
rect 22092 2746 22116 2748
rect 22172 2746 22196 2748
rect 22252 2746 22258 2748
rect 22012 2694 22014 2746
rect 22194 2694 22196 2746
rect 21950 2692 21956 2694
rect 22012 2692 22036 2694
rect 22092 2692 22116 2694
rect 22172 2692 22196 2694
rect 22252 2692 22258 2694
rect 21950 2683 22258 2692
rect 26950 2748 27258 2757
rect 26950 2746 26956 2748
rect 27012 2746 27036 2748
rect 27092 2746 27116 2748
rect 27172 2746 27196 2748
rect 27252 2746 27258 2748
rect 27012 2694 27014 2746
rect 27194 2694 27196 2746
rect 26950 2692 26956 2694
rect 27012 2692 27036 2694
rect 27092 2692 27116 2694
rect 27172 2692 27196 2694
rect 27252 2692 27258 2694
rect 26950 2683 27258 2692
rect 31950 2748 32258 2757
rect 31950 2746 31956 2748
rect 32012 2746 32036 2748
rect 32092 2746 32116 2748
rect 32172 2746 32196 2748
rect 32252 2746 32258 2748
rect 32012 2694 32014 2746
rect 32194 2694 32196 2746
rect 31950 2692 31956 2694
rect 32012 2692 32036 2694
rect 32092 2692 32116 2694
rect 32172 2692 32196 2694
rect 32252 2692 32258 2694
rect 31950 2683 32258 2692
rect 36648 2650 36676 18362
rect 36950 17980 37258 17989
rect 36950 17978 36956 17980
rect 37012 17978 37036 17980
rect 37092 17978 37116 17980
rect 37172 17978 37196 17980
rect 37252 17978 37258 17980
rect 37012 17926 37014 17978
rect 37194 17926 37196 17978
rect 36950 17924 36956 17926
rect 37012 17924 37036 17926
rect 37092 17924 37116 17926
rect 37172 17924 37196 17926
rect 37252 17924 37258 17926
rect 36950 17915 37258 17924
rect 38212 17610 38240 46990
rect 38292 32360 38344 32366
rect 38292 32302 38344 32308
rect 38200 17604 38252 17610
rect 38200 17546 38252 17552
rect 37610 17436 37918 17445
rect 37610 17434 37616 17436
rect 37672 17434 37696 17436
rect 37752 17434 37776 17436
rect 37832 17434 37856 17436
rect 37912 17434 37918 17436
rect 37672 17382 37674 17434
rect 37854 17382 37856 17434
rect 37610 17380 37616 17382
rect 37672 17380 37696 17382
rect 37752 17380 37776 17382
rect 37832 17380 37856 17382
rect 37912 17380 37918 17382
rect 37610 17371 37918 17380
rect 36950 16892 37258 16901
rect 36950 16890 36956 16892
rect 37012 16890 37036 16892
rect 37092 16890 37116 16892
rect 37172 16890 37196 16892
rect 37252 16890 37258 16892
rect 37012 16838 37014 16890
rect 37194 16838 37196 16890
rect 36950 16836 36956 16838
rect 37012 16836 37036 16838
rect 37092 16836 37116 16838
rect 37172 16836 37196 16838
rect 37252 16836 37258 16838
rect 36950 16827 37258 16836
rect 37610 16348 37918 16357
rect 37610 16346 37616 16348
rect 37672 16346 37696 16348
rect 37752 16346 37776 16348
rect 37832 16346 37856 16348
rect 37912 16346 37918 16348
rect 37672 16294 37674 16346
rect 37854 16294 37856 16346
rect 37610 16292 37616 16294
rect 37672 16292 37696 16294
rect 37752 16292 37776 16294
rect 37832 16292 37856 16294
rect 37912 16292 37918 16294
rect 37610 16283 37918 16292
rect 38200 15904 38252 15910
rect 38200 15846 38252 15852
rect 36950 15804 37258 15813
rect 36950 15802 36956 15804
rect 37012 15802 37036 15804
rect 37092 15802 37116 15804
rect 37172 15802 37196 15804
rect 37252 15802 37258 15804
rect 37012 15750 37014 15802
rect 37194 15750 37196 15802
rect 36950 15748 36956 15750
rect 37012 15748 37036 15750
rect 37092 15748 37116 15750
rect 37172 15748 37196 15750
rect 37252 15748 37258 15750
rect 36950 15739 37258 15748
rect 37610 15260 37918 15269
rect 37610 15258 37616 15260
rect 37672 15258 37696 15260
rect 37752 15258 37776 15260
rect 37832 15258 37856 15260
rect 37912 15258 37918 15260
rect 37672 15206 37674 15258
rect 37854 15206 37856 15258
rect 37610 15204 37616 15206
rect 37672 15204 37696 15206
rect 37752 15204 37776 15206
rect 37832 15204 37856 15206
rect 37912 15204 37918 15206
rect 37610 15195 37918 15204
rect 38212 15026 38240 15846
rect 38016 15020 38068 15026
rect 38016 14962 38068 14968
rect 38200 15020 38252 15026
rect 38200 14962 38252 14968
rect 36950 14716 37258 14725
rect 36950 14714 36956 14716
rect 37012 14714 37036 14716
rect 37092 14714 37116 14716
rect 37172 14714 37196 14716
rect 37252 14714 37258 14716
rect 37012 14662 37014 14714
rect 37194 14662 37196 14714
rect 36950 14660 36956 14662
rect 37012 14660 37036 14662
rect 37092 14660 37116 14662
rect 37172 14660 37196 14662
rect 37252 14660 37258 14662
rect 36950 14651 37258 14660
rect 37610 14172 37918 14181
rect 37610 14170 37616 14172
rect 37672 14170 37696 14172
rect 37752 14170 37776 14172
rect 37832 14170 37856 14172
rect 37912 14170 37918 14172
rect 37672 14118 37674 14170
rect 37854 14118 37856 14170
rect 37610 14116 37616 14118
rect 37672 14116 37696 14118
rect 37752 14116 37776 14118
rect 37832 14116 37856 14118
rect 37912 14116 37918 14118
rect 37610 14107 37918 14116
rect 36950 13628 37258 13637
rect 36950 13626 36956 13628
rect 37012 13626 37036 13628
rect 37092 13626 37116 13628
rect 37172 13626 37196 13628
rect 37252 13626 37258 13628
rect 37012 13574 37014 13626
rect 37194 13574 37196 13626
rect 36950 13572 36956 13574
rect 37012 13572 37036 13574
rect 37092 13572 37116 13574
rect 37172 13572 37196 13574
rect 37252 13572 37258 13574
rect 36950 13563 37258 13572
rect 37610 13084 37918 13093
rect 37610 13082 37616 13084
rect 37672 13082 37696 13084
rect 37752 13082 37776 13084
rect 37832 13082 37856 13084
rect 37912 13082 37918 13084
rect 37672 13030 37674 13082
rect 37854 13030 37856 13082
rect 37610 13028 37616 13030
rect 37672 13028 37696 13030
rect 37752 13028 37776 13030
rect 37832 13028 37856 13030
rect 37912 13028 37918 13030
rect 37610 13019 37918 13028
rect 36950 12540 37258 12549
rect 36950 12538 36956 12540
rect 37012 12538 37036 12540
rect 37092 12538 37116 12540
rect 37172 12538 37196 12540
rect 37252 12538 37258 12540
rect 37012 12486 37014 12538
rect 37194 12486 37196 12538
rect 36950 12484 36956 12486
rect 37012 12484 37036 12486
rect 37092 12484 37116 12486
rect 37172 12484 37196 12486
rect 37252 12484 37258 12486
rect 36950 12475 37258 12484
rect 37610 11996 37918 12005
rect 37610 11994 37616 11996
rect 37672 11994 37696 11996
rect 37752 11994 37776 11996
rect 37832 11994 37856 11996
rect 37912 11994 37918 11996
rect 37672 11942 37674 11994
rect 37854 11942 37856 11994
rect 37610 11940 37616 11942
rect 37672 11940 37696 11942
rect 37752 11940 37776 11942
rect 37832 11940 37856 11942
rect 37912 11940 37918 11942
rect 37610 11931 37918 11940
rect 36950 11452 37258 11461
rect 36950 11450 36956 11452
rect 37012 11450 37036 11452
rect 37092 11450 37116 11452
rect 37172 11450 37196 11452
rect 37252 11450 37258 11452
rect 37012 11398 37014 11450
rect 37194 11398 37196 11450
rect 36950 11396 36956 11398
rect 37012 11396 37036 11398
rect 37092 11396 37116 11398
rect 37172 11396 37196 11398
rect 37252 11396 37258 11398
rect 36950 11387 37258 11396
rect 37610 10908 37918 10917
rect 37610 10906 37616 10908
rect 37672 10906 37696 10908
rect 37752 10906 37776 10908
rect 37832 10906 37856 10908
rect 37912 10906 37918 10908
rect 37672 10854 37674 10906
rect 37854 10854 37856 10906
rect 37610 10852 37616 10854
rect 37672 10852 37696 10854
rect 37752 10852 37776 10854
rect 37832 10852 37856 10854
rect 37912 10852 37918 10854
rect 37610 10843 37918 10852
rect 36950 10364 37258 10373
rect 36950 10362 36956 10364
rect 37012 10362 37036 10364
rect 37092 10362 37116 10364
rect 37172 10362 37196 10364
rect 37252 10362 37258 10364
rect 37012 10310 37014 10362
rect 37194 10310 37196 10362
rect 36950 10308 36956 10310
rect 37012 10308 37036 10310
rect 37092 10308 37116 10310
rect 37172 10308 37196 10310
rect 37252 10308 37258 10310
rect 36950 10299 37258 10308
rect 37610 9820 37918 9829
rect 37610 9818 37616 9820
rect 37672 9818 37696 9820
rect 37752 9818 37776 9820
rect 37832 9818 37856 9820
rect 37912 9818 37918 9820
rect 37672 9766 37674 9818
rect 37854 9766 37856 9818
rect 37610 9764 37616 9766
rect 37672 9764 37696 9766
rect 37752 9764 37776 9766
rect 37832 9764 37856 9766
rect 37912 9764 37918 9766
rect 37610 9755 37918 9764
rect 36950 9276 37258 9285
rect 36950 9274 36956 9276
rect 37012 9274 37036 9276
rect 37092 9274 37116 9276
rect 37172 9274 37196 9276
rect 37252 9274 37258 9276
rect 37012 9222 37014 9274
rect 37194 9222 37196 9274
rect 36950 9220 36956 9222
rect 37012 9220 37036 9222
rect 37092 9220 37116 9222
rect 37172 9220 37196 9222
rect 37252 9220 37258 9222
rect 36950 9211 37258 9220
rect 38028 8974 38056 14962
rect 38016 8968 38068 8974
rect 38016 8910 38068 8916
rect 38212 8906 38240 14962
rect 38200 8900 38252 8906
rect 38200 8842 38252 8848
rect 37610 8732 37918 8741
rect 37610 8730 37616 8732
rect 37672 8730 37696 8732
rect 37752 8730 37776 8732
rect 37832 8730 37856 8732
rect 37912 8730 37918 8732
rect 37672 8678 37674 8730
rect 37854 8678 37856 8730
rect 37610 8676 37616 8678
rect 37672 8676 37696 8678
rect 37752 8676 37776 8678
rect 37832 8676 37856 8678
rect 37912 8676 37918 8678
rect 37610 8667 37918 8676
rect 36950 8188 37258 8197
rect 36950 8186 36956 8188
rect 37012 8186 37036 8188
rect 37092 8186 37116 8188
rect 37172 8186 37196 8188
rect 37252 8186 37258 8188
rect 37012 8134 37014 8186
rect 37194 8134 37196 8186
rect 36950 8132 36956 8134
rect 37012 8132 37036 8134
rect 37092 8132 37116 8134
rect 37172 8132 37196 8134
rect 37252 8132 37258 8134
rect 36950 8123 37258 8132
rect 37610 7644 37918 7653
rect 37610 7642 37616 7644
rect 37672 7642 37696 7644
rect 37752 7642 37776 7644
rect 37832 7642 37856 7644
rect 37912 7642 37918 7644
rect 37672 7590 37674 7642
rect 37854 7590 37856 7642
rect 37610 7588 37616 7590
rect 37672 7588 37696 7590
rect 37752 7588 37776 7590
rect 37832 7588 37856 7590
rect 37912 7588 37918 7590
rect 37610 7579 37918 7588
rect 36950 7100 37258 7109
rect 36950 7098 36956 7100
rect 37012 7098 37036 7100
rect 37092 7098 37116 7100
rect 37172 7098 37196 7100
rect 37252 7098 37258 7100
rect 37012 7046 37014 7098
rect 37194 7046 37196 7098
rect 36950 7044 36956 7046
rect 37012 7044 37036 7046
rect 37092 7044 37116 7046
rect 37172 7044 37196 7046
rect 37252 7044 37258 7046
rect 36950 7035 37258 7044
rect 37610 6556 37918 6565
rect 37610 6554 37616 6556
rect 37672 6554 37696 6556
rect 37752 6554 37776 6556
rect 37832 6554 37856 6556
rect 37912 6554 37918 6556
rect 37672 6502 37674 6554
rect 37854 6502 37856 6554
rect 37610 6500 37616 6502
rect 37672 6500 37696 6502
rect 37752 6500 37776 6502
rect 37832 6500 37856 6502
rect 37912 6500 37918 6502
rect 37610 6491 37918 6500
rect 36950 6012 37258 6021
rect 36950 6010 36956 6012
rect 37012 6010 37036 6012
rect 37092 6010 37116 6012
rect 37172 6010 37196 6012
rect 37252 6010 37258 6012
rect 37012 5958 37014 6010
rect 37194 5958 37196 6010
rect 36950 5956 36956 5958
rect 37012 5956 37036 5958
rect 37092 5956 37116 5958
rect 37172 5956 37196 5958
rect 37252 5956 37258 5958
rect 36950 5947 37258 5956
rect 37610 5468 37918 5477
rect 37610 5466 37616 5468
rect 37672 5466 37696 5468
rect 37752 5466 37776 5468
rect 37832 5466 37856 5468
rect 37912 5466 37918 5468
rect 37672 5414 37674 5466
rect 37854 5414 37856 5466
rect 37610 5412 37616 5414
rect 37672 5412 37696 5414
rect 37752 5412 37776 5414
rect 37832 5412 37856 5414
rect 37912 5412 37918 5414
rect 37610 5403 37918 5412
rect 36950 4924 37258 4933
rect 36950 4922 36956 4924
rect 37012 4922 37036 4924
rect 37092 4922 37116 4924
rect 37172 4922 37196 4924
rect 37252 4922 37258 4924
rect 37012 4870 37014 4922
rect 37194 4870 37196 4922
rect 36950 4868 36956 4870
rect 37012 4868 37036 4870
rect 37092 4868 37116 4870
rect 37172 4868 37196 4870
rect 37252 4868 37258 4870
rect 36950 4859 37258 4868
rect 37610 4380 37918 4389
rect 37610 4378 37616 4380
rect 37672 4378 37696 4380
rect 37752 4378 37776 4380
rect 37832 4378 37856 4380
rect 37912 4378 37918 4380
rect 37672 4326 37674 4378
rect 37854 4326 37856 4378
rect 37610 4324 37616 4326
rect 37672 4324 37696 4326
rect 37752 4324 37776 4326
rect 37832 4324 37856 4326
rect 37912 4324 37918 4326
rect 37610 4315 37918 4324
rect 36950 3836 37258 3845
rect 36950 3834 36956 3836
rect 37012 3834 37036 3836
rect 37092 3834 37116 3836
rect 37172 3834 37196 3836
rect 37252 3834 37258 3836
rect 37012 3782 37014 3834
rect 37194 3782 37196 3834
rect 36950 3780 36956 3782
rect 37012 3780 37036 3782
rect 37092 3780 37116 3782
rect 37172 3780 37196 3782
rect 37252 3780 37258 3782
rect 36950 3771 37258 3780
rect 37610 3292 37918 3301
rect 37610 3290 37616 3292
rect 37672 3290 37696 3292
rect 37752 3290 37776 3292
rect 37832 3290 37856 3292
rect 37912 3290 37918 3292
rect 37672 3238 37674 3290
rect 37854 3238 37856 3290
rect 37610 3236 37616 3238
rect 37672 3236 37696 3238
rect 37752 3236 37776 3238
rect 37832 3236 37856 3238
rect 37912 3236 37918 3238
rect 37610 3227 37918 3236
rect 38304 3058 38332 32302
rect 38396 10538 38424 50322
rect 38488 12170 38516 60250
rect 38936 58540 38988 58546
rect 38936 58482 38988 58488
rect 38844 56432 38896 56438
rect 38844 56374 38896 56380
rect 38660 50244 38712 50250
rect 38660 50186 38712 50192
rect 38672 41414 38700 50186
rect 38672 41386 38792 41414
rect 38568 32768 38620 32774
rect 38568 32710 38620 32716
rect 38580 32366 38608 32710
rect 38660 32428 38712 32434
rect 38660 32370 38712 32376
rect 38568 32360 38620 32366
rect 38568 32302 38620 32308
rect 38580 27946 38608 32302
rect 38568 27940 38620 27946
rect 38568 27882 38620 27888
rect 38672 22982 38700 32370
rect 38660 22976 38712 22982
rect 38660 22918 38712 22924
rect 38476 12164 38528 12170
rect 38476 12106 38528 12112
rect 38384 10532 38436 10538
rect 38384 10474 38436 10480
rect 38764 4486 38792 41386
rect 38856 9382 38884 56374
rect 38948 51074 38976 58482
rect 39028 57860 39080 57866
rect 39028 57802 39080 57808
rect 39040 54738 39068 57802
rect 39028 54732 39080 54738
rect 39028 54674 39080 54680
rect 38948 51046 39068 51074
rect 39040 35494 39068 51046
rect 39028 35488 39080 35494
rect 39028 35430 39080 35436
rect 39132 30705 39160 69362
rect 39764 62280 39816 62286
rect 39764 62222 39816 62228
rect 39948 62280 40000 62286
rect 39948 62222 40000 62228
rect 39304 62212 39356 62218
rect 39304 62154 39356 62160
rect 39488 62212 39540 62218
rect 39488 62154 39540 62160
rect 39212 57928 39264 57934
rect 39212 57870 39264 57876
rect 39224 54670 39252 57870
rect 39316 57866 39344 62154
rect 39304 57860 39356 57866
rect 39304 57802 39356 57808
rect 39500 57050 39528 62154
rect 39672 57792 39724 57798
rect 39672 57734 39724 57740
rect 39488 57044 39540 57050
rect 39488 56986 39540 56992
rect 39212 54664 39264 54670
rect 39212 54606 39264 54612
rect 39500 32026 39528 56986
rect 39684 54670 39712 57734
rect 39672 54664 39724 54670
rect 39672 54606 39724 54612
rect 39580 54528 39632 54534
rect 39580 54470 39632 54476
rect 39488 32020 39540 32026
rect 39488 31962 39540 31968
rect 39118 30696 39174 30705
rect 39118 30631 39174 30640
rect 39592 20262 39620 54470
rect 39672 32020 39724 32026
rect 39672 31962 39724 31968
rect 39580 20256 39632 20262
rect 39580 20198 39632 20204
rect 38936 14408 38988 14414
rect 38934 14376 38936 14385
rect 38988 14376 38990 14385
rect 38934 14311 38990 14320
rect 39684 13394 39712 31962
rect 39776 31822 39804 62222
rect 39960 57458 39988 62222
rect 40408 62144 40460 62150
rect 40408 62086 40460 62092
rect 40132 57928 40184 57934
rect 40132 57870 40184 57876
rect 40144 57594 40172 57870
rect 40132 57588 40184 57594
rect 40132 57530 40184 57536
rect 39948 57452 40000 57458
rect 39948 57394 40000 57400
rect 39960 55282 39988 57394
rect 39856 55276 39908 55282
rect 39856 55218 39908 55224
rect 39948 55276 40000 55282
rect 39948 55218 40000 55224
rect 39764 31816 39816 31822
rect 39764 31758 39816 31764
rect 39776 16454 39804 31758
rect 39868 18698 39896 55218
rect 40224 47660 40276 47666
rect 40224 47602 40276 47608
rect 40040 37460 40092 37466
rect 40040 37402 40092 37408
rect 40052 30666 40080 37402
rect 40236 36242 40264 47602
rect 40224 36236 40276 36242
rect 40224 36178 40276 36184
rect 40132 32564 40184 32570
rect 40132 32506 40184 32512
rect 40144 32026 40172 32506
rect 40132 32020 40184 32026
rect 40132 31962 40184 31968
rect 40040 30660 40092 30666
rect 40040 30602 40092 30608
rect 40236 29170 40264 36178
rect 40224 29164 40276 29170
rect 40224 29106 40276 29112
rect 40420 20534 40448 62086
rect 40500 36168 40552 36174
rect 40500 36110 40552 36116
rect 40512 36009 40540 36110
rect 40498 36000 40554 36009
rect 40498 35935 40554 35944
rect 40408 20528 40460 20534
rect 40408 20470 40460 20476
rect 39856 18692 39908 18698
rect 39856 18634 39908 18640
rect 39764 16448 39816 16454
rect 39764 16390 39816 16396
rect 39672 13388 39724 13394
rect 39672 13330 39724 13336
rect 38844 9376 38896 9382
rect 38844 9318 38896 9324
rect 38752 4480 38804 4486
rect 38752 4422 38804 4428
rect 38292 3052 38344 3058
rect 38292 2994 38344 3000
rect 36950 2748 37258 2757
rect 36950 2746 36956 2748
rect 37012 2746 37036 2748
rect 37092 2746 37116 2748
rect 37172 2746 37196 2748
rect 37252 2746 37258 2748
rect 37012 2694 37014 2746
rect 37194 2694 37196 2746
rect 36950 2692 36956 2694
rect 37012 2692 37036 2694
rect 37092 2692 37116 2694
rect 37172 2692 37196 2694
rect 37252 2692 37258 2694
rect 36950 2683 37258 2692
rect 36636 2644 36688 2650
rect 36636 2586 36688 2592
rect 30852 2514 31156 2530
rect 18604 2508 18656 2514
rect 18604 2450 18656 2456
rect 30840 2508 31156 2514
rect 30892 2502 31156 2508
rect 30840 2450 30892 2456
rect 31128 2446 31156 2502
rect 31116 2440 31168 2446
rect 31116 2382 31168 2388
rect 39304 2440 39356 2446
rect 39304 2382 39356 2388
rect 10232 2372 10284 2378
rect 10232 2314 10284 2320
rect 8024 2304 8076 2310
rect 8024 2246 8076 2252
rect 13084 2304 13136 2310
rect 13084 2246 13136 2252
rect 18328 2304 18380 2310
rect 18328 2246 18380 2252
rect 23572 2304 23624 2310
rect 23572 2246 23624 2252
rect 28816 2304 28868 2310
rect 28816 2246 28868 2252
rect 34060 2304 34112 2310
rect 34060 2246 34112 2252
rect 2610 2204 2918 2213
rect 2610 2202 2616 2204
rect 2672 2202 2696 2204
rect 2752 2202 2776 2204
rect 2832 2202 2856 2204
rect 2912 2202 2918 2204
rect 2672 2150 2674 2202
rect 2854 2150 2856 2202
rect 2610 2148 2616 2150
rect 2672 2148 2696 2150
rect 2752 2148 2776 2150
rect 2832 2148 2856 2150
rect 2912 2148 2918 2150
rect 2610 2139 2918 2148
rect 7610 2204 7918 2213
rect 7610 2202 7616 2204
rect 7672 2202 7696 2204
rect 7752 2202 7776 2204
rect 7832 2202 7856 2204
rect 7912 2202 7918 2204
rect 7672 2150 7674 2202
rect 7854 2150 7856 2202
rect 7610 2148 7616 2150
rect 7672 2148 7696 2150
rect 7752 2148 7776 2150
rect 7832 2148 7856 2150
rect 7912 2148 7918 2150
rect 7610 2139 7918 2148
rect 2516 1278 2636 1306
rect 2608 800 2636 1278
rect 8036 1170 8064 2246
rect 12610 2204 12918 2213
rect 12610 2202 12616 2204
rect 12672 2202 12696 2204
rect 12752 2202 12776 2204
rect 12832 2202 12856 2204
rect 12912 2202 12918 2204
rect 12672 2150 12674 2202
rect 12854 2150 12856 2202
rect 12610 2148 12616 2150
rect 12672 2148 12696 2150
rect 12752 2148 12776 2150
rect 12832 2148 12856 2150
rect 12912 2148 12918 2150
rect 12610 2139 12918 2148
rect 7852 1142 8064 1170
rect 7852 800 7880 1142
rect 13096 800 13124 2246
rect 17610 2204 17918 2213
rect 17610 2202 17616 2204
rect 17672 2202 17696 2204
rect 17752 2202 17776 2204
rect 17832 2202 17856 2204
rect 17912 2202 17918 2204
rect 17672 2150 17674 2202
rect 17854 2150 17856 2202
rect 17610 2148 17616 2150
rect 17672 2148 17696 2150
rect 17752 2148 17776 2150
rect 17832 2148 17856 2150
rect 17912 2148 17918 2150
rect 17610 2139 17918 2148
rect 18340 800 18368 2246
rect 22610 2204 22918 2213
rect 22610 2202 22616 2204
rect 22672 2202 22696 2204
rect 22752 2202 22776 2204
rect 22832 2202 22856 2204
rect 22912 2202 22918 2204
rect 22672 2150 22674 2202
rect 22854 2150 22856 2202
rect 22610 2148 22616 2150
rect 22672 2148 22696 2150
rect 22752 2148 22776 2150
rect 22832 2148 22856 2150
rect 22912 2148 22918 2150
rect 22610 2139 22918 2148
rect 23584 800 23612 2246
rect 27610 2204 27918 2213
rect 27610 2202 27616 2204
rect 27672 2202 27696 2204
rect 27752 2202 27776 2204
rect 27832 2202 27856 2204
rect 27912 2202 27918 2204
rect 27672 2150 27674 2202
rect 27854 2150 27856 2202
rect 27610 2148 27616 2150
rect 27672 2148 27696 2150
rect 27752 2148 27776 2150
rect 27832 2148 27856 2150
rect 27912 2148 27918 2150
rect 27610 2139 27918 2148
rect 28828 800 28856 2246
rect 32610 2204 32918 2213
rect 32610 2202 32616 2204
rect 32672 2202 32696 2204
rect 32752 2202 32776 2204
rect 32832 2202 32856 2204
rect 32912 2202 32918 2204
rect 32672 2150 32674 2202
rect 32854 2150 32856 2202
rect 32610 2148 32616 2150
rect 32672 2148 32696 2150
rect 32752 2148 32776 2150
rect 32832 2148 32856 2150
rect 32912 2148 32918 2150
rect 32610 2139 32918 2148
rect 34072 800 34100 2246
rect 37610 2204 37918 2213
rect 37610 2202 37616 2204
rect 37672 2202 37696 2204
rect 37752 2202 37776 2204
rect 37832 2202 37856 2204
rect 37912 2202 37918 2204
rect 37672 2150 37674 2202
rect 37854 2150 37856 2202
rect 37610 2148 37616 2150
rect 37672 2148 37696 2150
rect 37752 2148 37776 2150
rect 37832 2148 37856 2150
rect 37912 2148 37918 2150
rect 37610 2139 37918 2148
rect 39316 800 39344 2382
rect 2594 0 2650 800
rect 7838 0 7894 800
rect 13082 0 13138 800
rect 18326 0 18382 800
rect 23570 0 23626 800
rect 28814 0 28870 800
rect 34058 0 34114 800
rect 39302 0 39358 800
<< via2 >>
rect 2616 69658 2672 69660
rect 2696 69658 2752 69660
rect 2776 69658 2832 69660
rect 2856 69658 2912 69660
rect 2616 69606 2662 69658
rect 2662 69606 2672 69658
rect 2696 69606 2726 69658
rect 2726 69606 2738 69658
rect 2738 69606 2752 69658
rect 2776 69606 2790 69658
rect 2790 69606 2802 69658
rect 2802 69606 2832 69658
rect 2856 69606 2866 69658
rect 2866 69606 2912 69658
rect 2616 69604 2672 69606
rect 2696 69604 2752 69606
rect 2776 69604 2832 69606
rect 2856 69604 2912 69606
rect 7616 69658 7672 69660
rect 7696 69658 7752 69660
rect 7776 69658 7832 69660
rect 7856 69658 7912 69660
rect 7616 69606 7662 69658
rect 7662 69606 7672 69658
rect 7696 69606 7726 69658
rect 7726 69606 7738 69658
rect 7738 69606 7752 69658
rect 7776 69606 7790 69658
rect 7790 69606 7802 69658
rect 7802 69606 7832 69658
rect 7856 69606 7866 69658
rect 7866 69606 7912 69658
rect 7616 69604 7672 69606
rect 7696 69604 7752 69606
rect 7776 69604 7832 69606
rect 7856 69604 7912 69606
rect 12616 69658 12672 69660
rect 12696 69658 12752 69660
rect 12776 69658 12832 69660
rect 12856 69658 12912 69660
rect 12616 69606 12662 69658
rect 12662 69606 12672 69658
rect 12696 69606 12726 69658
rect 12726 69606 12738 69658
rect 12738 69606 12752 69658
rect 12776 69606 12790 69658
rect 12790 69606 12802 69658
rect 12802 69606 12832 69658
rect 12856 69606 12866 69658
rect 12866 69606 12912 69658
rect 12616 69604 12672 69606
rect 12696 69604 12752 69606
rect 12776 69604 12832 69606
rect 12856 69604 12912 69606
rect 17616 69658 17672 69660
rect 17696 69658 17752 69660
rect 17776 69658 17832 69660
rect 17856 69658 17912 69660
rect 17616 69606 17662 69658
rect 17662 69606 17672 69658
rect 17696 69606 17726 69658
rect 17726 69606 17738 69658
rect 17738 69606 17752 69658
rect 17776 69606 17790 69658
rect 17790 69606 17802 69658
rect 17802 69606 17832 69658
rect 17856 69606 17866 69658
rect 17866 69606 17912 69658
rect 17616 69604 17672 69606
rect 17696 69604 17752 69606
rect 17776 69604 17832 69606
rect 17856 69604 17912 69606
rect 22616 69658 22672 69660
rect 22696 69658 22752 69660
rect 22776 69658 22832 69660
rect 22856 69658 22912 69660
rect 22616 69606 22662 69658
rect 22662 69606 22672 69658
rect 22696 69606 22726 69658
rect 22726 69606 22738 69658
rect 22738 69606 22752 69658
rect 22776 69606 22790 69658
rect 22790 69606 22802 69658
rect 22802 69606 22832 69658
rect 22856 69606 22866 69658
rect 22866 69606 22912 69658
rect 22616 69604 22672 69606
rect 22696 69604 22752 69606
rect 22776 69604 22832 69606
rect 22856 69604 22912 69606
rect 27616 69658 27672 69660
rect 27696 69658 27752 69660
rect 27776 69658 27832 69660
rect 27856 69658 27912 69660
rect 27616 69606 27662 69658
rect 27662 69606 27672 69658
rect 27696 69606 27726 69658
rect 27726 69606 27738 69658
rect 27738 69606 27752 69658
rect 27776 69606 27790 69658
rect 27790 69606 27802 69658
rect 27802 69606 27832 69658
rect 27856 69606 27866 69658
rect 27866 69606 27912 69658
rect 27616 69604 27672 69606
rect 27696 69604 27752 69606
rect 27776 69604 27832 69606
rect 27856 69604 27912 69606
rect 32616 69658 32672 69660
rect 32696 69658 32752 69660
rect 32776 69658 32832 69660
rect 32856 69658 32912 69660
rect 32616 69606 32662 69658
rect 32662 69606 32672 69658
rect 32696 69606 32726 69658
rect 32726 69606 32738 69658
rect 32738 69606 32752 69658
rect 32776 69606 32790 69658
rect 32790 69606 32802 69658
rect 32802 69606 32832 69658
rect 32856 69606 32866 69658
rect 32866 69606 32912 69658
rect 32616 69604 32672 69606
rect 32696 69604 32752 69606
rect 32776 69604 32832 69606
rect 32856 69604 32912 69606
rect 37616 69658 37672 69660
rect 37696 69658 37752 69660
rect 37776 69658 37832 69660
rect 37856 69658 37912 69660
rect 37616 69606 37662 69658
rect 37662 69606 37672 69658
rect 37696 69606 37726 69658
rect 37726 69606 37738 69658
rect 37738 69606 37752 69658
rect 37776 69606 37790 69658
rect 37790 69606 37802 69658
rect 37802 69606 37832 69658
rect 37856 69606 37866 69658
rect 37866 69606 37912 69658
rect 37616 69604 37672 69606
rect 37696 69604 37752 69606
rect 37776 69604 37832 69606
rect 37856 69604 37912 69606
rect 1956 69114 2012 69116
rect 2036 69114 2092 69116
rect 2116 69114 2172 69116
rect 2196 69114 2252 69116
rect 1956 69062 2002 69114
rect 2002 69062 2012 69114
rect 2036 69062 2066 69114
rect 2066 69062 2078 69114
rect 2078 69062 2092 69114
rect 2116 69062 2130 69114
rect 2130 69062 2142 69114
rect 2142 69062 2172 69114
rect 2196 69062 2206 69114
rect 2206 69062 2252 69114
rect 1956 69060 2012 69062
rect 2036 69060 2092 69062
rect 2116 69060 2172 69062
rect 2196 69060 2252 69062
rect 2616 68570 2672 68572
rect 2696 68570 2752 68572
rect 2776 68570 2832 68572
rect 2856 68570 2912 68572
rect 2616 68518 2662 68570
rect 2662 68518 2672 68570
rect 2696 68518 2726 68570
rect 2726 68518 2738 68570
rect 2738 68518 2752 68570
rect 2776 68518 2790 68570
rect 2790 68518 2802 68570
rect 2802 68518 2832 68570
rect 2856 68518 2866 68570
rect 2866 68518 2912 68570
rect 2616 68516 2672 68518
rect 2696 68516 2752 68518
rect 2776 68516 2832 68518
rect 2856 68516 2912 68518
rect 1956 68026 2012 68028
rect 2036 68026 2092 68028
rect 2116 68026 2172 68028
rect 2196 68026 2252 68028
rect 1956 67974 2002 68026
rect 2002 67974 2012 68026
rect 2036 67974 2066 68026
rect 2066 67974 2078 68026
rect 2078 67974 2092 68026
rect 2116 67974 2130 68026
rect 2130 67974 2142 68026
rect 2142 67974 2172 68026
rect 2196 67974 2206 68026
rect 2206 67974 2252 68026
rect 1956 67972 2012 67974
rect 2036 67972 2092 67974
rect 2116 67972 2172 67974
rect 2196 67972 2252 67974
rect 1956 66938 2012 66940
rect 2036 66938 2092 66940
rect 2116 66938 2172 66940
rect 2196 66938 2252 66940
rect 1956 66886 2002 66938
rect 2002 66886 2012 66938
rect 2036 66886 2066 66938
rect 2066 66886 2078 66938
rect 2078 66886 2092 66938
rect 2116 66886 2130 66938
rect 2130 66886 2142 66938
rect 2142 66886 2172 66938
rect 2196 66886 2206 66938
rect 2206 66886 2252 66938
rect 1956 66884 2012 66886
rect 2036 66884 2092 66886
rect 2116 66884 2172 66886
rect 2196 66884 2252 66886
rect 1956 65850 2012 65852
rect 2036 65850 2092 65852
rect 2116 65850 2172 65852
rect 2196 65850 2252 65852
rect 1956 65798 2002 65850
rect 2002 65798 2012 65850
rect 2036 65798 2066 65850
rect 2066 65798 2078 65850
rect 2078 65798 2092 65850
rect 2116 65798 2130 65850
rect 2130 65798 2142 65850
rect 2142 65798 2172 65850
rect 2196 65798 2206 65850
rect 2206 65798 2252 65850
rect 1956 65796 2012 65798
rect 2036 65796 2092 65798
rect 2116 65796 2172 65798
rect 2196 65796 2252 65798
rect 1956 64762 2012 64764
rect 2036 64762 2092 64764
rect 2116 64762 2172 64764
rect 2196 64762 2252 64764
rect 1956 64710 2002 64762
rect 2002 64710 2012 64762
rect 2036 64710 2066 64762
rect 2066 64710 2078 64762
rect 2078 64710 2092 64762
rect 2116 64710 2130 64762
rect 2130 64710 2142 64762
rect 2142 64710 2172 64762
rect 2196 64710 2206 64762
rect 2206 64710 2252 64762
rect 1956 64708 2012 64710
rect 2036 64708 2092 64710
rect 2116 64708 2172 64710
rect 2196 64708 2252 64710
rect 1956 63674 2012 63676
rect 2036 63674 2092 63676
rect 2116 63674 2172 63676
rect 2196 63674 2252 63676
rect 1956 63622 2002 63674
rect 2002 63622 2012 63674
rect 2036 63622 2066 63674
rect 2066 63622 2078 63674
rect 2078 63622 2092 63674
rect 2116 63622 2130 63674
rect 2130 63622 2142 63674
rect 2142 63622 2172 63674
rect 2196 63622 2206 63674
rect 2206 63622 2252 63674
rect 1956 63620 2012 63622
rect 2036 63620 2092 63622
rect 2116 63620 2172 63622
rect 2196 63620 2252 63622
rect 1956 62586 2012 62588
rect 2036 62586 2092 62588
rect 2116 62586 2172 62588
rect 2196 62586 2252 62588
rect 1956 62534 2002 62586
rect 2002 62534 2012 62586
rect 2036 62534 2066 62586
rect 2066 62534 2078 62586
rect 2078 62534 2092 62586
rect 2116 62534 2130 62586
rect 2130 62534 2142 62586
rect 2142 62534 2172 62586
rect 2196 62534 2206 62586
rect 2206 62534 2252 62586
rect 1956 62532 2012 62534
rect 2036 62532 2092 62534
rect 2116 62532 2172 62534
rect 2196 62532 2252 62534
rect 1956 61498 2012 61500
rect 2036 61498 2092 61500
rect 2116 61498 2172 61500
rect 2196 61498 2252 61500
rect 1956 61446 2002 61498
rect 2002 61446 2012 61498
rect 2036 61446 2066 61498
rect 2066 61446 2078 61498
rect 2078 61446 2092 61498
rect 2116 61446 2130 61498
rect 2130 61446 2142 61498
rect 2142 61446 2172 61498
rect 2196 61446 2206 61498
rect 2206 61446 2252 61498
rect 1956 61444 2012 61446
rect 2036 61444 2092 61446
rect 2116 61444 2172 61446
rect 2196 61444 2252 61446
rect 1956 60410 2012 60412
rect 2036 60410 2092 60412
rect 2116 60410 2172 60412
rect 2196 60410 2252 60412
rect 1956 60358 2002 60410
rect 2002 60358 2012 60410
rect 2036 60358 2066 60410
rect 2066 60358 2078 60410
rect 2078 60358 2092 60410
rect 2116 60358 2130 60410
rect 2130 60358 2142 60410
rect 2142 60358 2172 60410
rect 2196 60358 2206 60410
rect 2206 60358 2252 60410
rect 1956 60356 2012 60358
rect 2036 60356 2092 60358
rect 2116 60356 2172 60358
rect 2196 60356 2252 60358
rect 1956 59322 2012 59324
rect 2036 59322 2092 59324
rect 2116 59322 2172 59324
rect 2196 59322 2252 59324
rect 1956 59270 2002 59322
rect 2002 59270 2012 59322
rect 2036 59270 2066 59322
rect 2066 59270 2078 59322
rect 2078 59270 2092 59322
rect 2116 59270 2130 59322
rect 2130 59270 2142 59322
rect 2142 59270 2172 59322
rect 2196 59270 2206 59322
rect 2206 59270 2252 59322
rect 1956 59268 2012 59270
rect 2036 59268 2092 59270
rect 2116 59268 2172 59270
rect 2196 59268 2252 59270
rect 1956 58234 2012 58236
rect 2036 58234 2092 58236
rect 2116 58234 2172 58236
rect 2196 58234 2252 58236
rect 1956 58182 2002 58234
rect 2002 58182 2012 58234
rect 2036 58182 2066 58234
rect 2066 58182 2078 58234
rect 2078 58182 2092 58234
rect 2116 58182 2130 58234
rect 2130 58182 2142 58234
rect 2142 58182 2172 58234
rect 2196 58182 2206 58234
rect 2206 58182 2252 58234
rect 1956 58180 2012 58182
rect 2036 58180 2092 58182
rect 2116 58180 2172 58182
rect 2196 58180 2252 58182
rect 1956 57146 2012 57148
rect 2036 57146 2092 57148
rect 2116 57146 2172 57148
rect 2196 57146 2252 57148
rect 1956 57094 2002 57146
rect 2002 57094 2012 57146
rect 2036 57094 2066 57146
rect 2066 57094 2078 57146
rect 2078 57094 2092 57146
rect 2116 57094 2130 57146
rect 2130 57094 2142 57146
rect 2142 57094 2172 57146
rect 2196 57094 2206 57146
rect 2206 57094 2252 57146
rect 1956 57092 2012 57094
rect 2036 57092 2092 57094
rect 2116 57092 2172 57094
rect 2196 57092 2252 57094
rect 1956 56058 2012 56060
rect 2036 56058 2092 56060
rect 2116 56058 2172 56060
rect 2196 56058 2252 56060
rect 1956 56006 2002 56058
rect 2002 56006 2012 56058
rect 2036 56006 2066 56058
rect 2066 56006 2078 56058
rect 2078 56006 2092 56058
rect 2116 56006 2130 56058
rect 2130 56006 2142 56058
rect 2142 56006 2172 56058
rect 2196 56006 2206 56058
rect 2206 56006 2252 56058
rect 1956 56004 2012 56006
rect 2036 56004 2092 56006
rect 2116 56004 2172 56006
rect 2196 56004 2252 56006
rect 1956 54970 2012 54972
rect 2036 54970 2092 54972
rect 2116 54970 2172 54972
rect 2196 54970 2252 54972
rect 1956 54918 2002 54970
rect 2002 54918 2012 54970
rect 2036 54918 2066 54970
rect 2066 54918 2078 54970
rect 2078 54918 2092 54970
rect 2116 54918 2130 54970
rect 2130 54918 2142 54970
rect 2142 54918 2172 54970
rect 2196 54918 2206 54970
rect 2206 54918 2252 54970
rect 1956 54916 2012 54918
rect 2036 54916 2092 54918
rect 2116 54916 2172 54918
rect 2196 54916 2252 54918
rect 1956 53882 2012 53884
rect 2036 53882 2092 53884
rect 2116 53882 2172 53884
rect 2196 53882 2252 53884
rect 1956 53830 2002 53882
rect 2002 53830 2012 53882
rect 2036 53830 2066 53882
rect 2066 53830 2078 53882
rect 2078 53830 2092 53882
rect 2116 53830 2130 53882
rect 2130 53830 2142 53882
rect 2142 53830 2172 53882
rect 2196 53830 2206 53882
rect 2206 53830 2252 53882
rect 1956 53828 2012 53830
rect 2036 53828 2092 53830
rect 2116 53828 2172 53830
rect 2196 53828 2252 53830
rect 1956 52794 2012 52796
rect 2036 52794 2092 52796
rect 2116 52794 2172 52796
rect 2196 52794 2252 52796
rect 1956 52742 2002 52794
rect 2002 52742 2012 52794
rect 2036 52742 2066 52794
rect 2066 52742 2078 52794
rect 2078 52742 2092 52794
rect 2116 52742 2130 52794
rect 2130 52742 2142 52794
rect 2142 52742 2172 52794
rect 2196 52742 2206 52794
rect 2206 52742 2252 52794
rect 1956 52740 2012 52742
rect 2036 52740 2092 52742
rect 2116 52740 2172 52742
rect 2196 52740 2252 52742
rect 1956 51706 2012 51708
rect 2036 51706 2092 51708
rect 2116 51706 2172 51708
rect 2196 51706 2252 51708
rect 1956 51654 2002 51706
rect 2002 51654 2012 51706
rect 2036 51654 2066 51706
rect 2066 51654 2078 51706
rect 2078 51654 2092 51706
rect 2116 51654 2130 51706
rect 2130 51654 2142 51706
rect 2142 51654 2172 51706
rect 2196 51654 2206 51706
rect 2206 51654 2252 51706
rect 1956 51652 2012 51654
rect 2036 51652 2092 51654
rect 2116 51652 2172 51654
rect 2196 51652 2252 51654
rect 1956 50618 2012 50620
rect 2036 50618 2092 50620
rect 2116 50618 2172 50620
rect 2196 50618 2252 50620
rect 1956 50566 2002 50618
rect 2002 50566 2012 50618
rect 2036 50566 2066 50618
rect 2066 50566 2078 50618
rect 2078 50566 2092 50618
rect 2116 50566 2130 50618
rect 2130 50566 2142 50618
rect 2142 50566 2172 50618
rect 2196 50566 2206 50618
rect 2206 50566 2252 50618
rect 1956 50564 2012 50566
rect 2036 50564 2092 50566
rect 2116 50564 2172 50566
rect 2196 50564 2252 50566
rect 1956 49530 2012 49532
rect 2036 49530 2092 49532
rect 2116 49530 2172 49532
rect 2196 49530 2252 49532
rect 1956 49478 2002 49530
rect 2002 49478 2012 49530
rect 2036 49478 2066 49530
rect 2066 49478 2078 49530
rect 2078 49478 2092 49530
rect 2116 49478 2130 49530
rect 2130 49478 2142 49530
rect 2142 49478 2172 49530
rect 2196 49478 2206 49530
rect 2206 49478 2252 49530
rect 1956 49476 2012 49478
rect 2036 49476 2092 49478
rect 2116 49476 2172 49478
rect 2196 49476 2252 49478
rect 1956 48442 2012 48444
rect 2036 48442 2092 48444
rect 2116 48442 2172 48444
rect 2196 48442 2252 48444
rect 1956 48390 2002 48442
rect 2002 48390 2012 48442
rect 2036 48390 2066 48442
rect 2066 48390 2078 48442
rect 2078 48390 2092 48442
rect 2116 48390 2130 48442
rect 2130 48390 2142 48442
rect 2142 48390 2172 48442
rect 2196 48390 2206 48442
rect 2206 48390 2252 48442
rect 1956 48388 2012 48390
rect 2036 48388 2092 48390
rect 2116 48388 2172 48390
rect 2196 48388 2252 48390
rect 1956 47354 2012 47356
rect 2036 47354 2092 47356
rect 2116 47354 2172 47356
rect 2196 47354 2252 47356
rect 1956 47302 2002 47354
rect 2002 47302 2012 47354
rect 2036 47302 2066 47354
rect 2066 47302 2078 47354
rect 2078 47302 2092 47354
rect 2116 47302 2130 47354
rect 2130 47302 2142 47354
rect 2142 47302 2172 47354
rect 2196 47302 2206 47354
rect 2206 47302 2252 47354
rect 1956 47300 2012 47302
rect 2036 47300 2092 47302
rect 2116 47300 2172 47302
rect 2196 47300 2252 47302
rect 1956 46266 2012 46268
rect 2036 46266 2092 46268
rect 2116 46266 2172 46268
rect 2196 46266 2252 46268
rect 1956 46214 2002 46266
rect 2002 46214 2012 46266
rect 2036 46214 2066 46266
rect 2066 46214 2078 46266
rect 2078 46214 2092 46266
rect 2116 46214 2130 46266
rect 2130 46214 2142 46266
rect 2142 46214 2172 46266
rect 2196 46214 2206 46266
rect 2206 46214 2252 46266
rect 1956 46212 2012 46214
rect 2036 46212 2092 46214
rect 2116 46212 2172 46214
rect 2196 46212 2252 46214
rect 1956 45178 2012 45180
rect 2036 45178 2092 45180
rect 2116 45178 2172 45180
rect 2196 45178 2252 45180
rect 1956 45126 2002 45178
rect 2002 45126 2012 45178
rect 2036 45126 2066 45178
rect 2066 45126 2078 45178
rect 2078 45126 2092 45178
rect 2116 45126 2130 45178
rect 2130 45126 2142 45178
rect 2142 45126 2172 45178
rect 2196 45126 2206 45178
rect 2206 45126 2252 45178
rect 1956 45124 2012 45126
rect 2036 45124 2092 45126
rect 2116 45124 2172 45126
rect 2196 45124 2252 45126
rect 1956 44090 2012 44092
rect 2036 44090 2092 44092
rect 2116 44090 2172 44092
rect 2196 44090 2252 44092
rect 1956 44038 2002 44090
rect 2002 44038 2012 44090
rect 2036 44038 2066 44090
rect 2066 44038 2078 44090
rect 2078 44038 2092 44090
rect 2116 44038 2130 44090
rect 2130 44038 2142 44090
rect 2142 44038 2172 44090
rect 2196 44038 2206 44090
rect 2206 44038 2252 44090
rect 1956 44036 2012 44038
rect 2036 44036 2092 44038
rect 2116 44036 2172 44038
rect 2196 44036 2252 44038
rect 1956 43002 2012 43004
rect 2036 43002 2092 43004
rect 2116 43002 2172 43004
rect 2196 43002 2252 43004
rect 1956 42950 2002 43002
rect 2002 42950 2012 43002
rect 2036 42950 2066 43002
rect 2066 42950 2078 43002
rect 2078 42950 2092 43002
rect 2116 42950 2130 43002
rect 2130 42950 2142 43002
rect 2142 42950 2172 43002
rect 2196 42950 2206 43002
rect 2206 42950 2252 43002
rect 1956 42948 2012 42950
rect 2036 42948 2092 42950
rect 2116 42948 2172 42950
rect 2196 42948 2252 42950
rect 1956 41914 2012 41916
rect 2036 41914 2092 41916
rect 2116 41914 2172 41916
rect 2196 41914 2252 41916
rect 1956 41862 2002 41914
rect 2002 41862 2012 41914
rect 2036 41862 2066 41914
rect 2066 41862 2078 41914
rect 2078 41862 2092 41914
rect 2116 41862 2130 41914
rect 2130 41862 2142 41914
rect 2142 41862 2172 41914
rect 2196 41862 2206 41914
rect 2206 41862 2252 41914
rect 1956 41860 2012 41862
rect 2036 41860 2092 41862
rect 2116 41860 2172 41862
rect 2196 41860 2252 41862
rect 1956 40826 2012 40828
rect 2036 40826 2092 40828
rect 2116 40826 2172 40828
rect 2196 40826 2252 40828
rect 1956 40774 2002 40826
rect 2002 40774 2012 40826
rect 2036 40774 2066 40826
rect 2066 40774 2078 40826
rect 2078 40774 2092 40826
rect 2116 40774 2130 40826
rect 2130 40774 2142 40826
rect 2142 40774 2172 40826
rect 2196 40774 2206 40826
rect 2206 40774 2252 40826
rect 1956 40772 2012 40774
rect 2036 40772 2092 40774
rect 2116 40772 2172 40774
rect 2196 40772 2252 40774
rect 1956 39738 2012 39740
rect 2036 39738 2092 39740
rect 2116 39738 2172 39740
rect 2196 39738 2252 39740
rect 1956 39686 2002 39738
rect 2002 39686 2012 39738
rect 2036 39686 2066 39738
rect 2066 39686 2078 39738
rect 2078 39686 2092 39738
rect 2116 39686 2130 39738
rect 2130 39686 2142 39738
rect 2142 39686 2172 39738
rect 2196 39686 2206 39738
rect 2206 39686 2252 39738
rect 1956 39684 2012 39686
rect 2036 39684 2092 39686
rect 2116 39684 2172 39686
rect 2196 39684 2252 39686
rect 1956 38650 2012 38652
rect 2036 38650 2092 38652
rect 2116 38650 2172 38652
rect 2196 38650 2252 38652
rect 1956 38598 2002 38650
rect 2002 38598 2012 38650
rect 2036 38598 2066 38650
rect 2066 38598 2078 38650
rect 2078 38598 2092 38650
rect 2116 38598 2130 38650
rect 2130 38598 2142 38650
rect 2142 38598 2172 38650
rect 2196 38598 2206 38650
rect 2206 38598 2252 38650
rect 1956 38596 2012 38598
rect 2036 38596 2092 38598
rect 2116 38596 2172 38598
rect 2196 38596 2252 38598
rect 1956 37562 2012 37564
rect 2036 37562 2092 37564
rect 2116 37562 2172 37564
rect 2196 37562 2252 37564
rect 1956 37510 2002 37562
rect 2002 37510 2012 37562
rect 2036 37510 2066 37562
rect 2066 37510 2078 37562
rect 2078 37510 2092 37562
rect 2116 37510 2130 37562
rect 2130 37510 2142 37562
rect 2142 37510 2172 37562
rect 2196 37510 2206 37562
rect 2206 37510 2252 37562
rect 1956 37508 2012 37510
rect 2036 37508 2092 37510
rect 2116 37508 2172 37510
rect 2196 37508 2252 37510
rect 1956 36474 2012 36476
rect 2036 36474 2092 36476
rect 2116 36474 2172 36476
rect 2196 36474 2252 36476
rect 1956 36422 2002 36474
rect 2002 36422 2012 36474
rect 2036 36422 2066 36474
rect 2066 36422 2078 36474
rect 2078 36422 2092 36474
rect 2116 36422 2130 36474
rect 2130 36422 2142 36474
rect 2142 36422 2172 36474
rect 2196 36422 2206 36474
rect 2206 36422 2252 36474
rect 1956 36420 2012 36422
rect 2036 36420 2092 36422
rect 2116 36420 2172 36422
rect 2196 36420 2252 36422
rect 1956 35386 2012 35388
rect 2036 35386 2092 35388
rect 2116 35386 2172 35388
rect 2196 35386 2252 35388
rect 1956 35334 2002 35386
rect 2002 35334 2012 35386
rect 2036 35334 2066 35386
rect 2066 35334 2078 35386
rect 2078 35334 2092 35386
rect 2116 35334 2130 35386
rect 2130 35334 2142 35386
rect 2142 35334 2172 35386
rect 2196 35334 2206 35386
rect 2206 35334 2252 35386
rect 1956 35332 2012 35334
rect 2036 35332 2092 35334
rect 2116 35332 2172 35334
rect 2196 35332 2252 35334
rect 1956 34298 2012 34300
rect 2036 34298 2092 34300
rect 2116 34298 2172 34300
rect 2196 34298 2252 34300
rect 1956 34246 2002 34298
rect 2002 34246 2012 34298
rect 2036 34246 2066 34298
rect 2066 34246 2078 34298
rect 2078 34246 2092 34298
rect 2116 34246 2130 34298
rect 2130 34246 2142 34298
rect 2142 34246 2172 34298
rect 2196 34246 2206 34298
rect 2206 34246 2252 34298
rect 1956 34244 2012 34246
rect 2036 34244 2092 34246
rect 2116 34244 2172 34246
rect 2196 34244 2252 34246
rect 1956 33210 2012 33212
rect 2036 33210 2092 33212
rect 2116 33210 2172 33212
rect 2196 33210 2252 33212
rect 1956 33158 2002 33210
rect 2002 33158 2012 33210
rect 2036 33158 2066 33210
rect 2066 33158 2078 33210
rect 2078 33158 2092 33210
rect 2116 33158 2130 33210
rect 2130 33158 2142 33210
rect 2142 33158 2172 33210
rect 2196 33158 2206 33210
rect 2206 33158 2252 33210
rect 1956 33156 2012 33158
rect 2036 33156 2092 33158
rect 2116 33156 2172 33158
rect 2196 33156 2252 33158
rect 1956 32122 2012 32124
rect 2036 32122 2092 32124
rect 2116 32122 2172 32124
rect 2196 32122 2252 32124
rect 1956 32070 2002 32122
rect 2002 32070 2012 32122
rect 2036 32070 2066 32122
rect 2066 32070 2078 32122
rect 2078 32070 2092 32122
rect 2116 32070 2130 32122
rect 2130 32070 2142 32122
rect 2142 32070 2172 32122
rect 2196 32070 2206 32122
rect 2206 32070 2252 32122
rect 1956 32068 2012 32070
rect 2036 32068 2092 32070
rect 2116 32068 2172 32070
rect 2196 32068 2252 32070
rect 1956 31034 2012 31036
rect 2036 31034 2092 31036
rect 2116 31034 2172 31036
rect 2196 31034 2252 31036
rect 1956 30982 2002 31034
rect 2002 30982 2012 31034
rect 2036 30982 2066 31034
rect 2066 30982 2078 31034
rect 2078 30982 2092 31034
rect 2116 30982 2130 31034
rect 2130 30982 2142 31034
rect 2142 30982 2172 31034
rect 2196 30982 2206 31034
rect 2206 30982 2252 31034
rect 1956 30980 2012 30982
rect 2036 30980 2092 30982
rect 2116 30980 2172 30982
rect 2196 30980 2252 30982
rect 1956 29946 2012 29948
rect 2036 29946 2092 29948
rect 2116 29946 2172 29948
rect 2196 29946 2252 29948
rect 1956 29894 2002 29946
rect 2002 29894 2012 29946
rect 2036 29894 2066 29946
rect 2066 29894 2078 29946
rect 2078 29894 2092 29946
rect 2116 29894 2130 29946
rect 2130 29894 2142 29946
rect 2142 29894 2172 29946
rect 2196 29894 2206 29946
rect 2206 29894 2252 29946
rect 1956 29892 2012 29894
rect 2036 29892 2092 29894
rect 2116 29892 2172 29894
rect 2196 29892 2252 29894
rect 1956 28858 2012 28860
rect 2036 28858 2092 28860
rect 2116 28858 2172 28860
rect 2196 28858 2252 28860
rect 1956 28806 2002 28858
rect 2002 28806 2012 28858
rect 2036 28806 2066 28858
rect 2066 28806 2078 28858
rect 2078 28806 2092 28858
rect 2116 28806 2130 28858
rect 2130 28806 2142 28858
rect 2142 28806 2172 28858
rect 2196 28806 2206 28858
rect 2206 28806 2252 28858
rect 1956 28804 2012 28806
rect 2036 28804 2092 28806
rect 2116 28804 2172 28806
rect 2196 28804 2252 28806
rect 1956 27770 2012 27772
rect 2036 27770 2092 27772
rect 2116 27770 2172 27772
rect 2196 27770 2252 27772
rect 1956 27718 2002 27770
rect 2002 27718 2012 27770
rect 2036 27718 2066 27770
rect 2066 27718 2078 27770
rect 2078 27718 2092 27770
rect 2116 27718 2130 27770
rect 2130 27718 2142 27770
rect 2142 27718 2172 27770
rect 2196 27718 2206 27770
rect 2206 27718 2252 27770
rect 1956 27716 2012 27718
rect 2036 27716 2092 27718
rect 2116 27716 2172 27718
rect 2196 27716 2252 27718
rect 1956 26682 2012 26684
rect 2036 26682 2092 26684
rect 2116 26682 2172 26684
rect 2196 26682 2252 26684
rect 1956 26630 2002 26682
rect 2002 26630 2012 26682
rect 2036 26630 2066 26682
rect 2066 26630 2078 26682
rect 2078 26630 2092 26682
rect 2116 26630 2130 26682
rect 2130 26630 2142 26682
rect 2142 26630 2172 26682
rect 2196 26630 2206 26682
rect 2206 26630 2252 26682
rect 1956 26628 2012 26630
rect 2036 26628 2092 26630
rect 2116 26628 2172 26630
rect 2196 26628 2252 26630
rect 1956 25594 2012 25596
rect 2036 25594 2092 25596
rect 2116 25594 2172 25596
rect 2196 25594 2252 25596
rect 1956 25542 2002 25594
rect 2002 25542 2012 25594
rect 2036 25542 2066 25594
rect 2066 25542 2078 25594
rect 2078 25542 2092 25594
rect 2116 25542 2130 25594
rect 2130 25542 2142 25594
rect 2142 25542 2172 25594
rect 2196 25542 2206 25594
rect 2206 25542 2252 25594
rect 1956 25540 2012 25542
rect 2036 25540 2092 25542
rect 2116 25540 2172 25542
rect 2196 25540 2252 25542
rect 1956 24506 2012 24508
rect 2036 24506 2092 24508
rect 2116 24506 2172 24508
rect 2196 24506 2252 24508
rect 1956 24454 2002 24506
rect 2002 24454 2012 24506
rect 2036 24454 2066 24506
rect 2066 24454 2078 24506
rect 2078 24454 2092 24506
rect 2116 24454 2130 24506
rect 2130 24454 2142 24506
rect 2142 24454 2172 24506
rect 2196 24454 2206 24506
rect 2206 24454 2252 24506
rect 1956 24452 2012 24454
rect 2036 24452 2092 24454
rect 2116 24452 2172 24454
rect 2196 24452 2252 24454
rect 2616 67482 2672 67484
rect 2696 67482 2752 67484
rect 2776 67482 2832 67484
rect 2856 67482 2912 67484
rect 2616 67430 2662 67482
rect 2662 67430 2672 67482
rect 2696 67430 2726 67482
rect 2726 67430 2738 67482
rect 2738 67430 2752 67482
rect 2776 67430 2790 67482
rect 2790 67430 2802 67482
rect 2802 67430 2832 67482
rect 2856 67430 2866 67482
rect 2866 67430 2912 67482
rect 2616 67428 2672 67430
rect 2696 67428 2752 67430
rect 2776 67428 2832 67430
rect 2856 67428 2912 67430
rect 2616 66394 2672 66396
rect 2696 66394 2752 66396
rect 2776 66394 2832 66396
rect 2856 66394 2912 66396
rect 2616 66342 2662 66394
rect 2662 66342 2672 66394
rect 2696 66342 2726 66394
rect 2726 66342 2738 66394
rect 2738 66342 2752 66394
rect 2776 66342 2790 66394
rect 2790 66342 2802 66394
rect 2802 66342 2832 66394
rect 2856 66342 2866 66394
rect 2866 66342 2912 66394
rect 2616 66340 2672 66342
rect 2696 66340 2752 66342
rect 2776 66340 2832 66342
rect 2856 66340 2912 66342
rect 2616 65306 2672 65308
rect 2696 65306 2752 65308
rect 2776 65306 2832 65308
rect 2856 65306 2912 65308
rect 2616 65254 2662 65306
rect 2662 65254 2672 65306
rect 2696 65254 2726 65306
rect 2726 65254 2738 65306
rect 2738 65254 2752 65306
rect 2776 65254 2790 65306
rect 2790 65254 2802 65306
rect 2802 65254 2832 65306
rect 2856 65254 2866 65306
rect 2866 65254 2912 65306
rect 2616 65252 2672 65254
rect 2696 65252 2752 65254
rect 2776 65252 2832 65254
rect 2856 65252 2912 65254
rect 2616 64218 2672 64220
rect 2696 64218 2752 64220
rect 2776 64218 2832 64220
rect 2856 64218 2912 64220
rect 2616 64166 2662 64218
rect 2662 64166 2672 64218
rect 2696 64166 2726 64218
rect 2726 64166 2738 64218
rect 2738 64166 2752 64218
rect 2776 64166 2790 64218
rect 2790 64166 2802 64218
rect 2802 64166 2832 64218
rect 2856 64166 2866 64218
rect 2866 64166 2912 64218
rect 2616 64164 2672 64166
rect 2696 64164 2752 64166
rect 2776 64164 2832 64166
rect 2856 64164 2912 64166
rect 2616 63130 2672 63132
rect 2696 63130 2752 63132
rect 2776 63130 2832 63132
rect 2856 63130 2912 63132
rect 2616 63078 2662 63130
rect 2662 63078 2672 63130
rect 2696 63078 2726 63130
rect 2726 63078 2738 63130
rect 2738 63078 2752 63130
rect 2776 63078 2790 63130
rect 2790 63078 2802 63130
rect 2802 63078 2832 63130
rect 2856 63078 2866 63130
rect 2866 63078 2912 63130
rect 2616 63076 2672 63078
rect 2696 63076 2752 63078
rect 2776 63076 2832 63078
rect 2856 63076 2912 63078
rect 2616 62042 2672 62044
rect 2696 62042 2752 62044
rect 2776 62042 2832 62044
rect 2856 62042 2912 62044
rect 2616 61990 2662 62042
rect 2662 61990 2672 62042
rect 2696 61990 2726 62042
rect 2726 61990 2738 62042
rect 2738 61990 2752 62042
rect 2776 61990 2790 62042
rect 2790 61990 2802 62042
rect 2802 61990 2832 62042
rect 2856 61990 2866 62042
rect 2866 61990 2912 62042
rect 2616 61988 2672 61990
rect 2696 61988 2752 61990
rect 2776 61988 2832 61990
rect 2856 61988 2912 61990
rect 2616 60954 2672 60956
rect 2696 60954 2752 60956
rect 2776 60954 2832 60956
rect 2856 60954 2912 60956
rect 2616 60902 2662 60954
rect 2662 60902 2672 60954
rect 2696 60902 2726 60954
rect 2726 60902 2738 60954
rect 2738 60902 2752 60954
rect 2776 60902 2790 60954
rect 2790 60902 2802 60954
rect 2802 60902 2832 60954
rect 2856 60902 2866 60954
rect 2866 60902 2912 60954
rect 2616 60900 2672 60902
rect 2696 60900 2752 60902
rect 2776 60900 2832 60902
rect 2856 60900 2912 60902
rect 2616 59866 2672 59868
rect 2696 59866 2752 59868
rect 2776 59866 2832 59868
rect 2856 59866 2912 59868
rect 2616 59814 2662 59866
rect 2662 59814 2672 59866
rect 2696 59814 2726 59866
rect 2726 59814 2738 59866
rect 2738 59814 2752 59866
rect 2776 59814 2790 59866
rect 2790 59814 2802 59866
rect 2802 59814 2832 59866
rect 2856 59814 2866 59866
rect 2866 59814 2912 59866
rect 2616 59812 2672 59814
rect 2696 59812 2752 59814
rect 2776 59812 2832 59814
rect 2856 59812 2912 59814
rect 2616 58778 2672 58780
rect 2696 58778 2752 58780
rect 2776 58778 2832 58780
rect 2856 58778 2912 58780
rect 2616 58726 2662 58778
rect 2662 58726 2672 58778
rect 2696 58726 2726 58778
rect 2726 58726 2738 58778
rect 2738 58726 2752 58778
rect 2776 58726 2790 58778
rect 2790 58726 2802 58778
rect 2802 58726 2832 58778
rect 2856 58726 2866 58778
rect 2866 58726 2912 58778
rect 2616 58724 2672 58726
rect 2696 58724 2752 58726
rect 2776 58724 2832 58726
rect 2856 58724 2912 58726
rect 6956 69114 7012 69116
rect 7036 69114 7092 69116
rect 7116 69114 7172 69116
rect 7196 69114 7252 69116
rect 6956 69062 7002 69114
rect 7002 69062 7012 69114
rect 7036 69062 7066 69114
rect 7066 69062 7078 69114
rect 7078 69062 7092 69114
rect 7116 69062 7130 69114
rect 7130 69062 7142 69114
rect 7142 69062 7172 69114
rect 7196 69062 7206 69114
rect 7206 69062 7252 69114
rect 6956 69060 7012 69062
rect 7036 69060 7092 69062
rect 7116 69060 7172 69062
rect 7196 69060 7252 69062
rect 7616 68570 7672 68572
rect 7696 68570 7752 68572
rect 7776 68570 7832 68572
rect 7856 68570 7912 68572
rect 7616 68518 7662 68570
rect 7662 68518 7672 68570
rect 7696 68518 7726 68570
rect 7726 68518 7738 68570
rect 7738 68518 7752 68570
rect 7776 68518 7790 68570
rect 7790 68518 7802 68570
rect 7802 68518 7832 68570
rect 7856 68518 7866 68570
rect 7866 68518 7912 68570
rect 7616 68516 7672 68518
rect 7696 68516 7752 68518
rect 7776 68516 7832 68518
rect 7856 68516 7912 68518
rect 2616 57690 2672 57692
rect 2696 57690 2752 57692
rect 2776 57690 2832 57692
rect 2856 57690 2912 57692
rect 2616 57638 2662 57690
rect 2662 57638 2672 57690
rect 2696 57638 2726 57690
rect 2726 57638 2738 57690
rect 2738 57638 2752 57690
rect 2776 57638 2790 57690
rect 2790 57638 2802 57690
rect 2802 57638 2832 57690
rect 2856 57638 2866 57690
rect 2866 57638 2912 57690
rect 2616 57636 2672 57638
rect 2696 57636 2752 57638
rect 2776 57636 2832 57638
rect 2856 57636 2912 57638
rect 2616 56602 2672 56604
rect 2696 56602 2752 56604
rect 2776 56602 2832 56604
rect 2856 56602 2912 56604
rect 2616 56550 2662 56602
rect 2662 56550 2672 56602
rect 2696 56550 2726 56602
rect 2726 56550 2738 56602
rect 2738 56550 2752 56602
rect 2776 56550 2790 56602
rect 2790 56550 2802 56602
rect 2802 56550 2832 56602
rect 2856 56550 2866 56602
rect 2866 56550 2912 56602
rect 2616 56548 2672 56550
rect 2696 56548 2752 56550
rect 2776 56548 2832 56550
rect 2856 56548 2912 56550
rect 2616 55514 2672 55516
rect 2696 55514 2752 55516
rect 2776 55514 2832 55516
rect 2856 55514 2912 55516
rect 2616 55462 2662 55514
rect 2662 55462 2672 55514
rect 2696 55462 2726 55514
rect 2726 55462 2738 55514
rect 2738 55462 2752 55514
rect 2776 55462 2790 55514
rect 2790 55462 2802 55514
rect 2802 55462 2832 55514
rect 2856 55462 2866 55514
rect 2866 55462 2912 55514
rect 2616 55460 2672 55462
rect 2696 55460 2752 55462
rect 2776 55460 2832 55462
rect 2856 55460 2912 55462
rect 2616 54426 2672 54428
rect 2696 54426 2752 54428
rect 2776 54426 2832 54428
rect 2856 54426 2912 54428
rect 2616 54374 2662 54426
rect 2662 54374 2672 54426
rect 2696 54374 2726 54426
rect 2726 54374 2738 54426
rect 2738 54374 2752 54426
rect 2776 54374 2790 54426
rect 2790 54374 2802 54426
rect 2802 54374 2832 54426
rect 2856 54374 2866 54426
rect 2866 54374 2912 54426
rect 2616 54372 2672 54374
rect 2696 54372 2752 54374
rect 2776 54372 2832 54374
rect 2856 54372 2912 54374
rect 2616 53338 2672 53340
rect 2696 53338 2752 53340
rect 2776 53338 2832 53340
rect 2856 53338 2912 53340
rect 2616 53286 2662 53338
rect 2662 53286 2672 53338
rect 2696 53286 2726 53338
rect 2726 53286 2738 53338
rect 2738 53286 2752 53338
rect 2776 53286 2790 53338
rect 2790 53286 2802 53338
rect 2802 53286 2832 53338
rect 2856 53286 2866 53338
rect 2866 53286 2912 53338
rect 2616 53284 2672 53286
rect 2696 53284 2752 53286
rect 2776 53284 2832 53286
rect 2856 53284 2912 53286
rect 2616 52250 2672 52252
rect 2696 52250 2752 52252
rect 2776 52250 2832 52252
rect 2856 52250 2912 52252
rect 2616 52198 2662 52250
rect 2662 52198 2672 52250
rect 2696 52198 2726 52250
rect 2726 52198 2738 52250
rect 2738 52198 2752 52250
rect 2776 52198 2790 52250
rect 2790 52198 2802 52250
rect 2802 52198 2832 52250
rect 2856 52198 2866 52250
rect 2866 52198 2912 52250
rect 2616 52196 2672 52198
rect 2696 52196 2752 52198
rect 2776 52196 2832 52198
rect 2856 52196 2912 52198
rect 2616 51162 2672 51164
rect 2696 51162 2752 51164
rect 2776 51162 2832 51164
rect 2856 51162 2912 51164
rect 2616 51110 2662 51162
rect 2662 51110 2672 51162
rect 2696 51110 2726 51162
rect 2726 51110 2738 51162
rect 2738 51110 2752 51162
rect 2776 51110 2790 51162
rect 2790 51110 2802 51162
rect 2802 51110 2832 51162
rect 2856 51110 2866 51162
rect 2866 51110 2912 51162
rect 2616 51108 2672 51110
rect 2696 51108 2752 51110
rect 2776 51108 2832 51110
rect 2856 51108 2912 51110
rect 2616 50074 2672 50076
rect 2696 50074 2752 50076
rect 2776 50074 2832 50076
rect 2856 50074 2912 50076
rect 2616 50022 2662 50074
rect 2662 50022 2672 50074
rect 2696 50022 2726 50074
rect 2726 50022 2738 50074
rect 2738 50022 2752 50074
rect 2776 50022 2790 50074
rect 2790 50022 2802 50074
rect 2802 50022 2832 50074
rect 2856 50022 2866 50074
rect 2866 50022 2912 50074
rect 2616 50020 2672 50022
rect 2696 50020 2752 50022
rect 2776 50020 2832 50022
rect 2856 50020 2912 50022
rect 2616 48986 2672 48988
rect 2696 48986 2752 48988
rect 2776 48986 2832 48988
rect 2856 48986 2912 48988
rect 2616 48934 2662 48986
rect 2662 48934 2672 48986
rect 2696 48934 2726 48986
rect 2726 48934 2738 48986
rect 2738 48934 2752 48986
rect 2776 48934 2790 48986
rect 2790 48934 2802 48986
rect 2802 48934 2832 48986
rect 2856 48934 2866 48986
rect 2866 48934 2912 48986
rect 2616 48932 2672 48934
rect 2696 48932 2752 48934
rect 2776 48932 2832 48934
rect 2856 48932 2912 48934
rect 2616 47898 2672 47900
rect 2696 47898 2752 47900
rect 2776 47898 2832 47900
rect 2856 47898 2912 47900
rect 2616 47846 2662 47898
rect 2662 47846 2672 47898
rect 2696 47846 2726 47898
rect 2726 47846 2738 47898
rect 2738 47846 2752 47898
rect 2776 47846 2790 47898
rect 2790 47846 2802 47898
rect 2802 47846 2832 47898
rect 2856 47846 2866 47898
rect 2866 47846 2912 47898
rect 2616 47844 2672 47846
rect 2696 47844 2752 47846
rect 2776 47844 2832 47846
rect 2856 47844 2912 47846
rect 2616 46810 2672 46812
rect 2696 46810 2752 46812
rect 2776 46810 2832 46812
rect 2856 46810 2912 46812
rect 2616 46758 2662 46810
rect 2662 46758 2672 46810
rect 2696 46758 2726 46810
rect 2726 46758 2738 46810
rect 2738 46758 2752 46810
rect 2776 46758 2790 46810
rect 2790 46758 2802 46810
rect 2802 46758 2832 46810
rect 2856 46758 2866 46810
rect 2866 46758 2912 46810
rect 2616 46756 2672 46758
rect 2696 46756 2752 46758
rect 2776 46756 2832 46758
rect 2856 46756 2912 46758
rect 2616 45722 2672 45724
rect 2696 45722 2752 45724
rect 2776 45722 2832 45724
rect 2856 45722 2912 45724
rect 2616 45670 2662 45722
rect 2662 45670 2672 45722
rect 2696 45670 2726 45722
rect 2726 45670 2738 45722
rect 2738 45670 2752 45722
rect 2776 45670 2790 45722
rect 2790 45670 2802 45722
rect 2802 45670 2832 45722
rect 2856 45670 2866 45722
rect 2866 45670 2912 45722
rect 2616 45668 2672 45670
rect 2696 45668 2752 45670
rect 2776 45668 2832 45670
rect 2856 45668 2912 45670
rect 1956 23418 2012 23420
rect 2036 23418 2092 23420
rect 2116 23418 2172 23420
rect 2196 23418 2252 23420
rect 1956 23366 2002 23418
rect 2002 23366 2012 23418
rect 2036 23366 2066 23418
rect 2066 23366 2078 23418
rect 2078 23366 2092 23418
rect 2116 23366 2130 23418
rect 2130 23366 2142 23418
rect 2142 23366 2172 23418
rect 2196 23366 2206 23418
rect 2206 23366 2252 23418
rect 1956 23364 2012 23366
rect 2036 23364 2092 23366
rect 2116 23364 2172 23366
rect 2196 23364 2252 23366
rect 1956 22330 2012 22332
rect 2036 22330 2092 22332
rect 2116 22330 2172 22332
rect 2196 22330 2252 22332
rect 1956 22278 2002 22330
rect 2002 22278 2012 22330
rect 2036 22278 2066 22330
rect 2066 22278 2078 22330
rect 2078 22278 2092 22330
rect 2116 22278 2130 22330
rect 2130 22278 2142 22330
rect 2142 22278 2172 22330
rect 2196 22278 2206 22330
rect 2206 22278 2252 22330
rect 1956 22276 2012 22278
rect 2036 22276 2092 22278
rect 2116 22276 2172 22278
rect 2196 22276 2252 22278
rect 1956 21242 2012 21244
rect 2036 21242 2092 21244
rect 2116 21242 2172 21244
rect 2196 21242 2252 21244
rect 1956 21190 2002 21242
rect 2002 21190 2012 21242
rect 2036 21190 2066 21242
rect 2066 21190 2078 21242
rect 2078 21190 2092 21242
rect 2116 21190 2130 21242
rect 2130 21190 2142 21242
rect 2142 21190 2172 21242
rect 2196 21190 2206 21242
rect 2206 21190 2252 21242
rect 1956 21188 2012 21190
rect 2036 21188 2092 21190
rect 2116 21188 2172 21190
rect 2196 21188 2252 21190
rect 1956 20154 2012 20156
rect 2036 20154 2092 20156
rect 2116 20154 2172 20156
rect 2196 20154 2252 20156
rect 1956 20102 2002 20154
rect 2002 20102 2012 20154
rect 2036 20102 2066 20154
rect 2066 20102 2078 20154
rect 2078 20102 2092 20154
rect 2116 20102 2130 20154
rect 2130 20102 2142 20154
rect 2142 20102 2172 20154
rect 2196 20102 2206 20154
rect 2206 20102 2252 20154
rect 1956 20100 2012 20102
rect 2036 20100 2092 20102
rect 2116 20100 2172 20102
rect 2196 20100 2252 20102
rect 1956 19066 2012 19068
rect 2036 19066 2092 19068
rect 2116 19066 2172 19068
rect 2196 19066 2252 19068
rect 1956 19014 2002 19066
rect 2002 19014 2012 19066
rect 2036 19014 2066 19066
rect 2066 19014 2078 19066
rect 2078 19014 2092 19066
rect 2116 19014 2130 19066
rect 2130 19014 2142 19066
rect 2142 19014 2172 19066
rect 2196 19014 2206 19066
rect 2206 19014 2252 19066
rect 1956 19012 2012 19014
rect 2036 19012 2092 19014
rect 2116 19012 2172 19014
rect 2196 19012 2252 19014
rect 1956 17978 2012 17980
rect 2036 17978 2092 17980
rect 2116 17978 2172 17980
rect 2196 17978 2252 17980
rect 1956 17926 2002 17978
rect 2002 17926 2012 17978
rect 2036 17926 2066 17978
rect 2066 17926 2078 17978
rect 2078 17926 2092 17978
rect 2116 17926 2130 17978
rect 2130 17926 2142 17978
rect 2142 17926 2172 17978
rect 2196 17926 2206 17978
rect 2206 17926 2252 17978
rect 1956 17924 2012 17926
rect 2036 17924 2092 17926
rect 2116 17924 2172 17926
rect 2196 17924 2252 17926
rect 1956 16890 2012 16892
rect 2036 16890 2092 16892
rect 2116 16890 2172 16892
rect 2196 16890 2252 16892
rect 1956 16838 2002 16890
rect 2002 16838 2012 16890
rect 2036 16838 2066 16890
rect 2066 16838 2078 16890
rect 2078 16838 2092 16890
rect 2116 16838 2130 16890
rect 2130 16838 2142 16890
rect 2142 16838 2172 16890
rect 2196 16838 2206 16890
rect 2206 16838 2252 16890
rect 1956 16836 2012 16838
rect 2036 16836 2092 16838
rect 2116 16836 2172 16838
rect 2196 16836 2252 16838
rect 1956 15802 2012 15804
rect 2036 15802 2092 15804
rect 2116 15802 2172 15804
rect 2196 15802 2252 15804
rect 1956 15750 2002 15802
rect 2002 15750 2012 15802
rect 2036 15750 2066 15802
rect 2066 15750 2078 15802
rect 2078 15750 2092 15802
rect 2116 15750 2130 15802
rect 2130 15750 2142 15802
rect 2142 15750 2172 15802
rect 2196 15750 2206 15802
rect 2206 15750 2252 15802
rect 1956 15748 2012 15750
rect 2036 15748 2092 15750
rect 2116 15748 2172 15750
rect 2196 15748 2252 15750
rect 1956 14714 2012 14716
rect 2036 14714 2092 14716
rect 2116 14714 2172 14716
rect 2196 14714 2252 14716
rect 1956 14662 2002 14714
rect 2002 14662 2012 14714
rect 2036 14662 2066 14714
rect 2066 14662 2078 14714
rect 2078 14662 2092 14714
rect 2116 14662 2130 14714
rect 2130 14662 2142 14714
rect 2142 14662 2172 14714
rect 2196 14662 2206 14714
rect 2206 14662 2252 14714
rect 1956 14660 2012 14662
rect 2036 14660 2092 14662
rect 2116 14660 2172 14662
rect 2196 14660 2252 14662
rect 1956 13626 2012 13628
rect 2036 13626 2092 13628
rect 2116 13626 2172 13628
rect 2196 13626 2252 13628
rect 1956 13574 2002 13626
rect 2002 13574 2012 13626
rect 2036 13574 2066 13626
rect 2066 13574 2078 13626
rect 2078 13574 2092 13626
rect 2116 13574 2130 13626
rect 2130 13574 2142 13626
rect 2142 13574 2172 13626
rect 2196 13574 2206 13626
rect 2206 13574 2252 13626
rect 1956 13572 2012 13574
rect 2036 13572 2092 13574
rect 2116 13572 2172 13574
rect 2196 13572 2252 13574
rect 1956 12538 2012 12540
rect 2036 12538 2092 12540
rect 2116 12538 2172 12540
rect 2196 12538 2252 12540
rect 1956 12486 2002 12538
rect 2002 12486 2012 12538
rect 2036 12486 2066 12538
rect 2066 12486 2078 12538
rect 2078 12486 2092 12538
rect 2116 12486 2130 12538
rect 2130 12486 2142 12538
rect 2142 12486 2172 12538
rect 2196 12486 2206 12538
rect 2206 12486 2252 12538
rect 1956 12484 2012 12486
rect 2036 12484 2092 12486
rect 2116 12484 2172 12486
rect 2196 12484 2252 12486
rect 1956 11450 2012 11452
rect 2036 11450 2092 11452
rect 2116 11450 2172 11452
rect 2196 11450 2252 11452
rect 1956 11398 2002 11450
rect 2002 11398 2012 11450
rect 2036 11398 2066 11450
rect 2066 11398 2078 11450
rect 2078 11398 2092 11450
rect 2116 11398 2130 11450
rect 2130 11398 2142 11450
rect 2142 11398 2172 11450
rect 2196 11398 2206 11450
rect 2206 11398 2252 11450
rect 1956 11396 2012 11398
rect 2036 11396 2092 11398
rect 2116 11396 2172 11398
rect 2196 11396 2252 11398
rect 1956 10362 2012 10364
rect 2036 10362 2092 10364
rect 2116 10362 2172 10364
rect 2196 10362 2252 10364
rect 1956 10310 2002 10362
rect 2002 10310 2012 10362
rect 2036 10310 2066 10362
rect 2066 10310 2078 10362
rect 2078 10310 2092 10362
rect 2116 10310 2130 10362
rect 2130 10310 2142 10362
rect 2142 10310 2172 10362
rect 2196 10310 2206 10362
rect 2206 10310 2252 10362
rect 1956 10308 2012 10310
rect 2036 10308 2092 10310
rect 2116 10308 2172 10310
rect 2196 10308 2252 10310
rect 1956 9274 2012 9276
rect 2036 9274 2092 9276
rect 2116 9274 2172 9276
rect 2196 9274 2252 9276
rect 1956 9222 2002 9274
rect 2002 9222 2012 9274
rect 2036 9222 2066 9274
rect 2066 9222 2078 9274
rect 2078 9222 2092 9274
rect 2116 9222 2130 9274
rect 2130 9222 2142 9274
rect 2142 9222 2172 9274
rect 2196 9222 2206 9274
rect 2206 9222 2252 9274
rect 1956 9220 2012 9222
rect 2036 9220 2092 9222
rect 2116 9220 2172 9222
rect 2196 9220 2252 9222
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 2616 44634 2672 44636
rect 2696 44634 2752 44636
rect 2776 44634 2832 44636
rect 2856 44634 2912 44636
rect 2616 44582 2662 44634
rect 2662 44582 2672 44634
rect 2696 44582 2726 44634
rect 2726 44582 2738 44634
rect 2738 44582 2752 44634
rect 2776 44582 2790 44634
rect 2790 44582 2802 44634
rect 2802 44582 2832 44634
rect 2856 44582 2866 44634
rect 2866 44582 2912 44634
rect 2616 44580 2672 44582
rect 2696 44580 2752 44582
rect 2776 44580 2832 44582
rect 2856 44580 2912 44582
rect 2616 43546 2672 43548
rect 2696 43546 2752 43548
rect 2776 43546 2832 43548
rect 2856 43546 2912 43548
rect 2616 43494 2662 43546
rect 2662 43494 2672 43546
rect 2696 43494 2726 43546
rect 2726 43494 2738 43546
rect 2738 43494 2752 43546
rect 2776 43494 2790 43546
rect 2790 43494 2802 43546
rect 2802 43494 2832 43546
rect 2856 43494 2866 43546
rect 2866 43494 2912 43546
rect 2616 43492 2672 43494
rect 2696 43492 2752 43494
rect 2776 43492 2832 43494
rect 2856 43492 2912 43494
rect 2616 42458 2672 42460
rect 2696 42458 2752 42460
rect 2776 42458 2832 42460
rect 2856 42458 2912 42460
rect 2616 42406 2662 42458
rect 2662 42406 2672 42458
rect 2696 42406 2726 42458
rect 2726 42406 2738 42458
rect 2738 42406 2752 42458
rect 2776 42406 2790 42458
rect 2790 42406 2802 42458
rect 2802 42406 2832 42458
rect 2856 42406 2866 42458
rect 2866 42406 2912 42458
rect 2616 42404 2672 42406
rect 2696 42404 2752 42406
rect 2776 42404 2832 42406
rect 2856 42404 2912 42406
rect 2616 41370 2672 41372
rect 2696 41370 2752 41372
rect 2776 41370 2832 41372
rect 2856 41370 2912 41372
rect 2616 41318 2662 41370
rect 2662 41318 2672 41370
rect 2696 41318 2726 41370
rect 2726 41318 2738 41370
rect 2738 41318 2752 41370
rect 2776 41318 2790 41370
rect 2790 41318 2802 41370
rect 2802 41318 2832 41370
rect 2856 41318 2866 41370
rect 2866 41318 2912 41370
rect 2616 41316 2672 41318
rect 2696 41316 2752 41318
rect 2776 41316 2832 41318
rect 2856 41316 2912 41318
rect 2616 40282 2672 40284
rect 2696 40282 2752 40284
rect 2776 40282 2832 40284
rect 2856 40282 2912 40284
rect 2616 40230 2662 40282
rect 2662 40230 2672 40282
rect 2696 40230 2726 40282
rect 2726 40230 2738 40282
rect 2738 40230 2752 40282
rect 2776 40230 2790 40282
rect 2790 40230 2802 40282
rect 2802 40230 2832 40282
rect 2856 40230 2866 40282
rect 2866 40230 2912 40282
rect 2616 40228 2672 40230
rect 2696 40228 2752 40230
rect 2776 40228 2832 40230
rect 2856 40228 2912 40230
rect 2616 39194 2672 39196
rect 2696 39194 2752 39196
rect 2776 39194 2832 39196
rect 2856 39194 2912 39196
rect 2616 39142 2662 39194
rect 2662 39142 2672 39194
rect 2696 39142 2726 39194
rect 2726 39142 2738 39194
rect 2738 39142 2752 39194
rect 2776 39142 2790 39194
rect 2790 39142 2802 39194
rect 2802 39142 2832 39194
rect 2856 39142 2866 39194
rect 2866 39142 2912 39194
rect 2616 39140 2672 39142
rect 2696 39140 2752 39142
rect 2776 39140 2832 39142
rect 2856 39140 2912 39142
rect 2616 38106 2672 38108
rect 2696 38106 2752 38108
rect 2776 38106 2832 38108
rect 2856 38106 2912 38108
rect 2616 38054 2662 38106
rect 2662 38054 2672 38106
rect 2696 38054 2726 38106
rect 2726 38054 2738 38106
rect 2738 38054 2752 38106
rect 2776 38054 2790 38106
rect 2790 38054 2802 38106
rect 2802 38054 2832 38106
rect 2856 38054 2866 38106
rect 2866 38054 2912 38106
rect 2616 38052 2672 38054
rect 2696 38052 2752 38054
rect 2776 38052 2832 38054
rect 2856 38052 2912 38054
rect 2616 37018 2672 37020
rect 2696 37018 2752 37020
rect 2776 37018 2832 37020
rect 2856 37018 2912 37020
rect 2616 36966 2662 37018
rect 2662 36966 2672 37018
rect 2696 36966 2726 37018
rect 2726 36966 2738 37018
rect 2738 36966 2752 37018
rect 2776 36966 2790 37018
rect 2790 36966 2802 37018
rect 2802 36966 2832 37018
rect 2856 36966 2866 37018
rect 2866 36966 2912 37018
rect 2616 36964 2672 36966
rect 2696 36964 2752 36966
rect 2776 36964 2832 36966
rect 2856 36964 2912 36966
rect 2616 35930 2672 35932
rect 2696 35930 2752 35932
rect 2776 35930 2832 35932
rect 2856 35930 2912 35932
rect 2616 35878 2662 35930
rect 2662 35878 2672 35930
rect 2696 35878 2726 35930
rect 2726 35878 2738 35930
rect 2738 35878 2752 35930
rect 2776 35878 2790 35930
rect 2790 35878 2802 35930
rect 2802 35878 2832 35930
rect 2856 35878 2866 35930
rect 2866 35878 2912 35930
rect 2616 35876 2672 35878
rect 2696 35876 2752 35878
rect 2776 35876 2832 35878
rect 2856 35876 2912 35878
rect 2616 34842 2672 34844
rect 2696 34842 2752 34844
rect 2776 34842 2832 34844
rect 2856 34842 2912 34844
rect 2616 34790 2662 34842
rect 2662 34790 2672 34842
rect 2696 34790 2726 34842
rect 2726 34790 2738 34842
rect 2738 34790 2752 34842
rect 2776 34790 2790 34842
rect 2790 34790 2802 34842
rect 2802 34790 2832 34842
rect 2856 34790 2866 34842
rect 2866 34790 2912 34842
rect 2616 34788 2672 34790
rect 2696 34788 2752 34790
rect 2776 34788 2832 34790
rect 2856 34788 2912 34790
rect 2616 33754 2672 33756
rect 2696 33754 2752 33756
rect 2776 33754 2832 33756
rect 2856 33754 2912 33756
rect 2616 33702 2662 33754
rect 2662 33702 2672 33754
rect 2696 33702 2726 33754
rect 2726 33702 2738 33754
rect 2738 33702 2752 33754
rect 2776 33702 2790 33754
rect 2790 33702 2802 33754
rect 2802 33702 2832 33754
rect 2856 33702 2866 33754
rect 2866 33702 2912 33754
rect 2616 33700 2672 33702
rect 2696 33700 2752 33702
rect 2776 33700 2832 33702
rect 2856 33700 2912 33702
rect 2616 32666 2672 32668
rect 2696 32666 2752 32668
rect 2776 32666 2832 32668
rect 2856 32666 2912 32668
rect 2616 32614 2662 32666
rect 2662 32614 2672 32666
rect 2696 32614 2726 32666
rect 2726 32614 2738 32666
rect 2738 32614 2752 32666
rect 2776 32614 2790 32666
rect 2790 32614 2802 32666
rect 2802 32614 2832 32666
rect 2856 32614 2866 32666
rect 2866 32614 2912 32666
rect 2616 32612 2672 32614
rect 2696 32612 2752 32614
rect 2776 32612 2832 32614
rect 2856 32612 2912 32614
rect 2616 31578 2672 31580
rect 2696 31578 2752 31580
rect 2776 31578 2832 31580
rect 2856 31578 2912 31580
rect 2616 31526 2662 31578
rect 2662 31526 2672 31578
rect 2696 31526 2726 31578
rect 2726 31526 2738 31578
rect 2738 31526 2752 31578
rect 2776 31526 2790 31578
rect 2790 31526 2802 31578
rect 2802 31526 2832 31578
rect 2856 31526 2866 31578
rect 2866 31526 2912 31578
rect 2616 31524 2672 31526
rect 2696 31524 2752 31526
rect 2776 31524 2832 31526
rect 2856 31524 2912 31526
rect 2616 30490 2672 30492
rect 2696 30490 2752 30492
rect 2776 30490 2832 30492
rect 2856 30490 2912 30492
rect 2616 30438 2662 30490
rect 2662 30438 2672 30490
rect 2696 30438 2726 30490
rect 2726 30438 2738 30490
rect 2738 30438 2752 30490
rect 2776 30438 2790 30490
rect 2790 30438 2802 30490
rect 2802 30438 2832 30490
rect 2856 30438 2866 30490
rect 2866 30438 2912 30490
rect 2616 30436 2672 30438
rect 2696 30436 2752 30438
rect 2776 30436 2832 30438
rect 2856 30436 2912 30438
rect 2616 29402 2672 29404
rect 2696 29402 2752 29404
rect 2776 29402 2832 29404
rect 2856 29402 2912 29404
rect 2616 29350 2662 29402
rect 2662 29350 2672 29402
rect 2696 29350 2726 29402
rect 2726 29350 2738 29402
rect 2738 29350 2752 29402
rect 2776 29350 2790 29402
rect 2790 29350 2802 29402
rect 2802 29350 2832 29402
rect 2856 29350 2866 29402
rect 2866 29350 2912 29402
rect 2616 29348 2672 29350
rect 2696 29348 2752 29350
rect 2776 29348 2832 29350
rect 2856 29348 2912 29350
rect 2616 28314 2672 28316
rect 2696 28314 2752 28316
rect 2776 28314 2832 28316
rect 2856 28314 2912 28316
rect 2616 28262 2662 28314
rect 2662 28262 2672 28314
rect 2696 28262 2726 28314
rect 2726 28262 2738 28314
rect 2738 28262 2752 28314
rect 2776 28262 2790 28314
rect 2790 28262 2802 28314
rect 2802 28262 2832 28314
rect 2856 28262 2866 28314
rect 2866 28262 2912 28314
rect 2616 28260 2672 28262
rect 2696 28260 2752 28262
rect 2776 28260 2832 28262
rect 2856 28260 2912 28262
rect 2616 27226 2672 27228
rect 2696 27226 2752 27228
rect 2776 27226 2832 27228
rect 2856 27226 2912 27228
rect 2616 27174 2662 27226
rect 2662 27174 2672 27226
rect 2696 27174 2726 27226
rect 2726 27174 2738 27226
rect 2738 27174 2752 27226
rect 2776 27174 2790 27226
rect 2790 27174 2802 27226
rect 2802 27174 2832 27226
rect 2856 27174 2866 27226
rect 2866 27174 2912 27226
rect 2616 27172 2672 27174
rect 2696 27172 2752 27174
rect 2776 27172 2832 27174
rect 2856 27172 2912 27174
rect 2616 26138 2672 26140
rect 2696 26138 2752 26140
rect 2776 26138 2832 26140
rect 2856 26138 2912 26140
rect 2616 26086 2662 26138
rect 2662 26086 2672 26138
rect 2696 26086 2726 26138
rect 2726 26086 2738 26138
rect 2738 26086 2752 26138
rect 2776 26086 2790 26138
rect 2790 26086 2802 26138
rect 2802 26086 2832 26138
rect 2856 26086 2866 26138
rect 2866 26086 2912 26138
rect 2616 26084 2672 26086
rect 2696 26084 2752 26086
rect 2776 26084 2832 26086
rect 2856 26084 2912 26086
rect 2616 25050 2672 25052
rect 2696 25050 2752 25052
rect 2776 25050 2832 25052
rect 2856 25050 2912 25052
rect 2616 24998 2662 25050
rect 2662 24998 2672 25050
rect 2696 24998 2726 25050
rect 2726 24998 2738 25050
rect 2738 24998 2752 25050
rect 2776 24998 2790 25050
rect 2790 24998 2802 25050
rect 2802 24998 2832 25050
rect 2856 24998 2866 25050
rect 2866 24998 2912 25050
rect 2616 24996 2672 24998
rect 2696 24996 2752 24998
rect 2776 24996 2832 24998
rect 2856 24996 2912 24998
rect 2616 23962 2672 23964
rect 2696 23962 2752 23964
rect 2776 23962 2832 23964
rect 2856 23962 2912 23964
rect 2616 23910 2662 23962
rect 2662 23910 2672 23962
rect 2696 23910 2726 23962
rect 2726 23910 2738 23962
rect 2738 23910 2752 23962
rect 2776 23910 2790 23962
rect 2790 23910 2802 23962
rect 2802 23910 2832 23962
rect 2856 23910 2866 23962
rect 2866 23910 2912 23962
rect 2616 23908 2672 23910
rect 2696 23908 2752 23910
rect 2776 23908 2832 23910
rect 2856 23908 2912 23910
rect 2616 22874 2672 22876
rect 2696 22874 2752 22876
rect 2776 22874 2832 22876
rect 2856 22874 2912 22876
rect 2616 22822 2662 22874
rect 2662 22822 2672 22874
rect 2696 22822 2726 22874
rect 2726 22822 2738 22874
rect 2738 22822 2752 22874
rect 2776 22822 2790 22874
rect 2790 22822 2802 22874
rect 2802 22822 2832 22874
rect 2856 22822 2866 22874
rect 2866 22822 2912 22874
rect 2616 22820 2672 22822
rect 2696 22820 2752 22822
rect 2776 22820 2832 22822
rect 2856 22820 2912 22822
rect 2616 21786 2672 21788
rect 2696 21786 2752 21788
rect 2776 21786 2832 21788
rect 2856 21786 2912 21788
rect 2616 21734 2662 21786
rect 2662 21734 2672 21786
rect 2696 21734 2726 21786
rect 2726 21734 2738 21786
rect 2738 21734 2752 21786
rect 2776 21734 2790 21786
rect 2790 21734 2802 21786
rect 2802 21734 2832 21786
rect 2856 21734 2866 21786
rect 2866 21734 2912 21786
rect 2616 21732 2672 21734
rect 2696 21732 2752 21734
rect 2776 21732 2832 21734
rect 2856 21732 2912 21734
rect 2616 20698 2672 20700
rect 2696 20698 2752 20700
rect 2776 20698 2832 20700
rect 2856 20698 2912 20700
rect 2616 20646 2662 20698
rect 2662 20646 2672 20698
rect 2696 20646 2726 20698
rect 2726 20646 2738 20698
rect 2738 20646 2752 20698
rect 2776 20646 2790 20698
rect 2790 20646 2802 20698
rect 2802 20646 2832 20698
rect 2856 20646 2866 20698
rect 2866 20646 2912 20698
rect 2616 20644 2672 20646
rect 2696 20644 2752 20646
rect 2776 20644 2832 20646
rect 2856 20644 2912 20646
rect 2616 19610 2672 19612
rect 2696 19610 2752 19612
rect 2776 19610 2832 19612
rect 2856 19610 2912 19612
rect 2616 19558 2662 19610
rect 2662 19558 2672 19610
rect 2696 19558 2726 19610
rect 2726 19558 2738 19610
rect 2738 19558 2752 19610
rect 2776 19558 2790 19610
rect 2790 19558 2802 19610
rect 2802 19558 2832 19610
rect 2856 19558 2866 19610
rect 2866 19558 2912 19610
rect 2616 19556 2672 19558
rect 2696 19556 2752 19558
rect 2776 19556 2832 19558
rect 2856 19556 2912 19558
rect 2616 18522 2672 18524
rect 2696 18522 2752 18524
rect 2776 18522 2832 18524
rect 2856 18522 2912 18524
rect 2616 18470 2662 18522
rect 2662 18470 2672 18522
rect 2696 18470 2726 18522
rect 2726 18470 2738 18522
rect 2738 18470 2752 18522
rect 2776 18470 2790 18522
rect 2790 18470 2802 18522
rect 2802 18470 2832 18522
rect 2856 18470 2866 18522
rect 2866 18470 2912 18522
rect 2616 18468 2672 18470
rect 2696 18468 2752 18470
rect 2776 18468 2832 18470
rect 2856 18468 2912 18470
rect 2616 17434 2672 17436
rect 2696 17434 2752 17436
rect 2776 17434 2832 17436
rect 2856 17434 2912 17436
rect 2616 17382 2662 17434
rect 2662 17382 2672 17434
rect 2696 17382 2726 17434
rect 2726 17382 2738 17434
rect 2738 17382 2752 17434
rect 2776 17382 2790 17434
rect 2790 17382 2802 17434
rect 2802 17382 2832 17434
rect 2856 17382 2866 17434
rect 2866 17382 2912 17434
rect 2616 17380 2672 17382
rect 2696 17380 2752 17382
rect 2776 17380 2832 17382
rect 2856 17380 2912 17382
rect 2616 16346 2672 16348
rect 2696 16346 2752 16348
rect 2776 16346 2832 16348
rect 2856 16346 2912 16348
rect 2616 16294 2662 16346
rect 2662 16294 2672 16346
rect 2696 16294 2726 16346
rect 2726 16294 2738 16346
rect 2738 16294 2752 16346
rect 2776 16294 2790 16346
rect 2790 16294 2802 16346
rect 2802 16294 2832 16346
rect 2856 16294 2866 16346
rect 2866 16294 2912 16346
rect 2616 16292 2672 16294
rect 2696 16292 2752 16294
rect 2776 16292 2832 16294
rect 2856 16292 2912 16294
rect 2616 15258 2672 15260
rect 2696 15258 2752 15260
rect 2776 15258 2832 15260
rect 2856 15258 2912 15260
rect 2616 15206 2662 15258
rect 2662 15206 2672 15258
rect 2696 15206 2726 15258
rect 2726 15206 2738 15258
rect 2738 15206 2752 15258
rect 2776 15206 2790 15258
rect 2790 15206 2802 15258
rect 2802 15206 2832 15258
rect 2856 15206 2866 15258
rect 2866 15206 2912 15258
rect 2616 15204 2672 15206
rect 2696 15204 2752 15206
rect 2776 15204 2832 15206
rect 2856 15204 2912 15206
rect 2616 14170 2672 14172
rect 2696 14170 2752 14172
rect 2776 14170 2832 14172
rect 2856 14170 2912 14172
rect 2616 14118 2662 14170
rect 2662 14118 2672 14170
rect 2696 14118 2726 14170
rect 2726 14118 2738 14170
rect 2738 14118 2752 14170
rect 2776 14118 2790 14170
rect 2790 14118 2802 14170
rect 2802 14118 2832 14170
rect 2856 14118 2866 14170
rect 2866 14118 2912 14170
rect 2616 14116 2672 14118
rect 2696 14116 2752 14118
rect 2776 14116 2832 14118
rect 2856 14116 2912 14118
rect 2616 13082 2672 13084
rect 2696 13082 2752 13084
rect 2776 13082 2832 13084
rect 2856 13082 2912 13084
rect 2616 13030 2662 13082
rect 2662 13030 2672 13082
rect 2696 13030 2726 13082
rect 2726 13030 2738 13082
rect 2738 13030 2752 13082
rect 2776 13030 2790 13082
rect 2790 13030 2802 13082
rect 2802 13030 2832 13082
rect 2856 13030 2866 13082
rect 2866 13030 2912 13082
rect 2616 13028 2672 13030
rect 2696 13028 2752 13030
rect 2776 13028 2832 13030
rect 2856 13028 2912 13030
rect 2616 11994 2672 11996
rect 2696 11994 2752 11996
rect 2776 11994 2832 11996
rect 2856 11994 2912 11996
rect 2616 11942 2662 11994
rect 2662 11942 2672 11994
rect 2696 11942 2726 11994
rect 2726 11942 2738 11994
rect 2738 11942 2752 11994
rect 2776 11942 2790 11994
rect 2790 11942 2802 11994
rect 2802 11942 2832 11994
rect 2856 11942 2866 11994
rect 2866 11942 2912 11994
rect 2616 11940 2672 11942
rect 2696 11940 2752 11942
rect 2776 11940 2832 11942
rect 2856 11940 2912 11942
rect 2616 10906 2672 10908
rect 2696 10906 2752 10908
rect 2776 10906 2832 10908
rect 2856 10906 2912 10908
rect 2616 10854 2662 10906
rect 2662 10854 2672 10906
rect 2696 10854 2726 10906
rect 2726 10854 2738 10906
rect 2738 10854 2752 10906
rect 2776 10854 2790 10906
rect 2790 10854 2802 10906
rect 2802 10854 2832 10906
rect 2856 10854 2866 10906
rect 2866 10854 2912 10906
rect 2616 10852 2672 10854
rect 2696 10852 2752 10854
rect 2776 10852 2832 10854
rect 2856 10852 2912 10854
rect 2616 9818 2672 9820
rect 2696 9818 2752 9820
rect 2776 9818 2832 9820
rect 2856 9818 2912 9820
rect 2616 9766 2662 9818
rect 2662 9766 2672 9818
rect 2696 9766 2726 9818
rect 2726 9766 2738 9818
rect 2738 9766 2752 9818
rect 2776 9766 2790 9818
rect 2790 9766 2802 9818
rect 2802 9766 2832 9818
rect 2856 9766 2866 9818
rect 2866 9766 2912 9818
rect 2616 9764 2672 9766
rect 2696 9764 2752 9766
rect 2776 9764 2832 9766
rect 2856 9764 2912 9766
rect 2616 8730 2672 8732
rect 2696 8730 2752 8732
rect 2776 8730 2832 8732
rect 2856 8730 2912 8732
rect 2616 8678 2662 8730
rect 2662 8678 2672 8730
rect 2696 8678 2726 8730
rect 2726 8678 2738 8730
rect 2738 8678 2752 8730
rect 2776 8678 2790 8730
rect 2790 8678 2802 8730
rect 2802 8678 2832 8730
rect 2856 8678 2866 8730
rect 2866 8678 2912 8730
rect 2616 8676 2672 8678
rect 2696 8676 2752 8678
rect 2776 8676 2832 8678
rect 2856 8676 2912 8678
rect 2616 7642 2672 7644
rect 2696 7642 2752 7644
rect 2776 7642 2832 7644
rect 2856 7642 2912 7644
rect 2616 7590 2662 7642
rect 2662 7590 2672 7642
rect 2696 7590 2726 7642
rect 2726 7590 2738 7642
rect 2738 7590 2752 7642
rect 2776 7590 2790 7642
rect 2790 7590 2802 7642
rect 2802 7590 2832 7642
rect 2856 7590 2866 7642
rect 2866 7590 2912 7642
rect 2616 7588 2672 7590
rect 2696 7588 2752 7590
rect 2776 7588 2832 7590
rect 2856 7588 2912 7590
rect 2616 6554 2672 6556
rect 2696 6554 2752 6556
rect 2776 6554 2832 6556
rect 2856 6554 2912 6556
rect 2616 6502 2662 6554
rect 2662 6502 2672 6554
rect 2696 6502 2726 6554
rect 2726 6502 2738 6554
rect 2738 6502 2752 6554
rect 2776 6502 2790 6554
rect 2790 6502 2802 6554
rect 2802 6502 2832 6554
rect 2856 6502 2866 6554
rect 2866 6502 2912 6554
rect 2616 6500 2672 6502
rect 2696 6500 2752 6502
rect 2776 6500 2832 6502
rect 2856 6500 2912 6502
rect 2616 5466 2672 5468
rect 2696 5466 2752 5468
rect 2776 5466 2832 5468
rect 2856 5466 2912 5468
rect 2616 5414 2662 5466
rect 2662 5414 2672 5466
rect 2696 5414 2726 5466
rect 2726 5414 2738 5466
rect 2738 5414 2752 5466
rect 2776 5414 2790 5466
rect 2790 5414 2802 5466
rect 2802 5414 2832 5466
rect 2856 5414 2866 5466
rect 2866 5414 2912 5466
rect 2616 5412 2672 5414
rect 2696 5412 2752 5414
rect 2776 5412 2832 5414
rect 2856 5412 2912 5414
rect 2616 4378 2672 4380
rect 2696 4378 2752 4380
rect 2776 4378 2832 4380
rect 2856 4378 2912 4380
rect 2616 4326 2662 4378
rect 2662 4326 2672 4378
rect 2696 4326 2726 4378
rect 2726 4326 2738 4378
rect 2738 4326 2752 4378
rect 2776 4326 2790 4378
rect 2790 4326 2802 4378
rect 2802 4326 2832 4378
rect 2856 4326 2866 4378
rect 2866 4326 2912 4378
rect 2616 4324 2672 4326
rect 2696 4324 2752 4326
rect 2776 4324 2832 4326
rect 2856 4324 2912 4326
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 6956 68026 7012 68028
rect 7036 68026 7092 68028
rect 7116 68026 7172 68028
rect 7196 68026 7252 68028
rect 6956 67974 7002 68026
rect 7002 67974 7012 68026
rect 7036 67974 7066 68026
rect 7066 67974 7078 68026
rect 7078 67974 7092 68026
rect 7116 67974 7130 68026
rect 7130 67974 7142 68026
rect 7142 67974 7172 68026
rect 7196 67974 7206 68026
rect 7206 67974 7252 68026
rect 6956 67972 7012 67974
rect 7036 67972 7092 67974
rect 7116 67972 7172 67974
rect 7196 67972 7252 67974
rect 6956 66938 7012 66940
rect 7036 66938 7092 66940
rect 7116 66938 7172 66940
rect 7196 66938 7252 66940
rect 6956 66886 7002 66938
rect 7002 66886 7012 66938
rect 7036 66886 7066 66938
rect 7066 66886 7078 66938
rect 7078 66886 7092 66938
rect 7116 66886 7130 66938
rect 7130 66886 7142 66938
rect 7142 66886 7172 66938
rect 7196 66886 7206 66938
rect 7206 66886 7252 66938
rect 6956 66884 7012 66886
rect 7036 66884 7092 66886
rect 7116 66884 7172 66886
rect 7196 66884 7252 66886
rect 6956 65850 7012 65852
rect 7036 65850 7092 65852
rect 7116 65850 7172 65852
rect 7196 65850 7252 65852
rect 6956 65798 7002 65850
rect 7002 65798 7012 65850
rect 7036 65798 7066 65850
rect 7066 65798 7078 65850
rect 7078 65798 7092 65850
rect 7116 65798 7130 65850
rect 7130 65798 7142 65850
rect 7142 65798 7172 65850
rect 7196 65798 7206 65850
rect 7206 65798 7252 65850
rect 6956 65796 7012 65798
rect 7036 65796 7092 65798
rect 7116 65796 7172 65798
rect 7196 65796 7252 65798
rect 6956 64762 7012 64764
rect 7036 64762 7092 64764
rect 7116 64762 7172 64764
rect 7196 64762 7252 64764
rect 6956 64710 7002 64762
rect 7002 64710 7012 64762
rect 7036 64710 7066 64762
rect 7066 64710 7078 64762
rect 7078 64710 7092 64762
rect 7116 64710 7130 64762
rect 7130 64710 7142 64762
rect 7142 64710 7172 64762
rect 7196 64710 7206 64762
rect 7206 64710 7252 64762
rect 6956 64708 7012 64710
rect 7036 64708 7092 64710
rect 7116 64708 7172 64710
rect 7196 64708 7252 64710
rect 6956 63674 7012 63676
rect 7036 63674 7092 63676
rect 7116 63674 7172 63676
rect 7196 63674 7252 63676
rect 6956 63622 7002 63674
rect 7002 63622 7012 63674
rect 7036 63622 7066 63674
rect 7066 63622 7078 63674
rect 7078 63622 7092 63674
rect 7116 63622 7130 63674
rect 7130 63622 7142 63674
rect 7142 63622 7172 63674
rect 7196 63622 7206 63674
rect 7206 63622 7252 63674
rect 6956 63620 7012 63622
rect 7036 63620 7092 63622
rect 7116 63620 7172 63622
rect 7196 63620 7252 63622
rect 6956 62586 7012 62588
rect 7036 62586 7092 62588
rect 7116 62586 7172 62588
rect 7196 62586 7252 62588
rect 6956 62534 7002 62586
rect 7002 62534 7012 62586
rect 7036 62534 7066 62586
rect 7066 62534 7078 62586
rect 7078 62534 7092 62586
rect 7116 62534 7130 62586
rect 7130 62534 7142 62586
rect 7142 62534 7172 62586
rect 7196 62534 7206 62586
rect 7206 62534 7252 62586
rect 6956 62532 7012 62534
rect 7036 62532 7092 62534
rect 7116 62532 7172 62534
rect 7196 62532 7252 62534
rect 6956 61498 7012 61500
rect 7036 61498 7092 61500
rect 7116 61498 7172 61500
rect 7196 61498 7252 61500
rect 6956 61446 7002 61498
rect 7002 61446 7012 61498
rect 7036 61446 7066 61498
rect 7066 61446 7078 61498
rect 7078 61446 7092 61498
rect 7116 61446 7130 61498
rect 7130 61446 7142 61498
rect 7142 61446 7172 61498
rect 7196 61446 7206 61498
rect 7206 61446 7252 61498
rect 6956 61444 7012 61446
rect 7036 61444 7092 61446
rect 7116 61444 7172 61446
rect 7196 61444 7252 61446
rect 6956 60410 7012 60412
rect 7036 60410 7092 60412
rect 7116 60410 7172 60412
rect 7196 60410 7252 60412
rect 6956 60358 7002 60410
rect 7002 60358 7012 60410
rect 7036 60358 7066 60410
rect 7066 60358 7078 60410
rect 7078 60358 7092 60410
rect 7116 60358 7130 60410
rect 7130 60358 7142 60410
rect 7142 60358 7172 60410
rect 7196 60358 7206 60410
rect 7206 60358 7252 60410
rect 6956 60356 7012 60358
rect 7036 60356 7092 60358
rect 7116 60356 7172 60358
rect 7196 60356 7252 60358
rect 6956 59322 7012 59324
rect 7036 59322 7092 59324
rect 7116 59322 7172 59324
rect 7196 59322 7252 59324
rect 6956 59270 7002 59322
rect 7002 59270 7012 59322
rect 7036 59270 7066 59322
rect 7066 59270 7078 59322
rect 7078 59270 7092 59322
rect 7116 59270 7130 59322
rect 7130 59270 7142 59322
rect 7142 59270 7172 59322
rect 7196 59270 7206 59322
rect 7206 59270 7252 59322
rect 6956 59268 7012 59270
rect 7036 59268 7092 59270
rect 7116 59268 7172 59270
rect 7196 59268 7252 59270
rect 6956 58234 7012 58236
rect 7036 58234 7092 58236
rect 7116 58234 7172 58236
rect 7196 58234 7252 58236
rect 6956 58182 7002 58234
rect 7002 58182 7012 58234
rect 7036 58182 7066 58234
rect 7066 58182 7078 58234
rect 7078 58182 7092 58234
rect 7116 58182 7130 58234
rect 7130 58182 7142 58234
rect 7142 58182 7172 58234
rect 7196 58182 7206 58234
rect 7206 58182 7252 58234
rect 6956 58180 7012 58182
rect 7036 58180 7092 58182
rect 7116 58180 7172 58182
rect 7196 58180 7252 58182
rect 6956 57146 7012 57148
rect 7036 57146 7092 57148
rect 7116 57146 7172 57148
rect 7196 57146 7252 57148
rect 6956 57094 7002 57146
rect 7002 57094 7012 57146
rect 7036 57094 7066 57146
rect 7066 57094 7078 57146
rect 7078 57094 7092 57146
rect 7116 57094 7130 57146
rect 7130 57094 7142 57146
rect 7142 57094 7172 57146
rect 7196 57094 7206 57146
rect 7206 57094 7252 57146
rect 6956 57092 7012 57094
rect 7036 57092 7092 57094
rect 7116 57092 7172 57094
rect 7196 57092 7252 57094
rect 6956 56058 7012 56060
rect 7036 56058 7092 56060
rect 7116 56058 7172 56060
rect 7196 56058 7252 56060
rect 6956 56006 7002 56058
rect 7002 56006 7012 56058
rect 7036 56006 7066 56058
rect 7066 56006 7078 56058
rect 7078 56006 7092 56058
rect 7116 56006 7130 56058
rect 7130 56006 7142 56058
rect 7142 56006 7172 56058
rect 7196 56006 7206 56058
rect 7206 56006 7252 56058
rect 6956 56004 7012 56006
rect 7036 56004 7092 56006
rect 7116 56004 7172 56006
rect 7196 56004 7252 56006
rect 3238 22636 3294 22672
rect 3238 22616 3240 22636
rect 3240 22616 3292 22636
rect 3292 22616 3294 22636
rect 2616 3290 2672 3292
rect 2696 3290 2752 3292
rect 2776 3290 2832 3292
rect 2856 3290 2912 3292
rect 2616 3238 2662 3290
rect 2662 3238 2672 3290
rect 2696 3238 2726 3290
rect 2726 3238 2738 3290
rect 2738 3238 2752 3290
rect 2776 3238 2790 3290
rect 2790 3238 2802 3290
rect 2802 3238 2832 3290
rect 2856 3238 2866 3290
rect 2866 3238 2912 3290
rect 2616 3236 2672 3238
rect 2696 3236 2752 3238
rect 2776 3236 2832 3238
rect 2856 3236 2912 3238
rect 6956 54970 7012 54972
rect 7036 54970 7092 54972
rect 7116 54970 7172 54972
rect 7196 54970 7252 54972
rect 6956 54918 7002 54970
rect 7002 54918 7012 54970
rect 7036 54918 7066 54970
rect 7066 54918 7078 54970
rect 7078 54918 7092 54970
rect 7116 54918 7130 54970
rect 7130 54918 7142 54970
rect 7142 54918 7172 54970
rect 7196 54918 7206 54970
rect 7206 54918 7252 54970
rect 6956 54916 7012 54918
rect 7036 54916 7092 54918
rect 7116 54916 7172 54918
rect 7196 54916 7252 54918
rect 6956 53882 7012 53884
rect 7036 53882 7092 53884
rect 7116 53882 7172 53884
rect 7196 53882 7252 53884
rect 6956 53830 7002 53882
rect 7002 53830 7012 53882
rect 7036 53830 7066 53882
rect 7066 53830 7078 53882
rect 7078 53830 7092 53882
rect 7116 53830 7130 53882
rect 7130 53830 7142 53882
rect 7142 53830 7172 53882
rect 7196 53830 7206 53882
rect 7206 53830 7252 53882
rect 6956 53828 7012 53830
rect 7036 53828 7092 53830
rect 7116 53828 7172 53830
rect 7196 53828 7252 53830
rect 6956 52794 7012 52796
rect 7036 52794 7092 52796
rect 7116 52794 7172 52796
rect 7196 52794 7252 52796
rect 6956 52742 7002 52794
rect 7002 52742 7012 52794
rect 7036 52742 7066 52794
rect 7066 52742 7078 52794
rect 7078 52742 7092 52794
rect 7116 52742 7130 52794
rect 7130 52742 7142 52794
rect 7142 52742 7172 52794
rect 7196 52742 7206 52794
rect 7206 52742 7252 52794
rect 6956 52740 7012 52742
rect 7036 52740 7092 52742
rect 7116 52740 7172 52742
rect 7196 52740 7252 52742
rect 6956 51706 7012 51708
rect 7036 51706 7092 51708
rect 7116 51706 7172 51708
rect 7196 51706 7252 51708
rect 6956 51654 7002 51706
rect 7002 51654 7012 51706
rect 7036 51654 7066 51706
rect 7066 51654 7078 51706
rect 7078 51654 7092 51706
rect 7116 51654 7130 51706
rect 7130 51654 7142 51706
rect 7142 51654 7172 51706
rect 7196 51654 7206 51706
rect 7206 51654 7252 51706
rect 6956 51652 7012 51654
rect 7036 51652 7092 51654
rect 7116 51652 7172 51654
rect 7196 51652 7252 51654
rect 6956 50618 7012 50620
rect 7036 50618 7092 50620
rect 7116 50618 7172 50620
rect 7196 50618 7252 50620
rect 6956 50566 7002 50618
rect 7002 50566 7012 50618
rect 7036 50566 7066 50618
rect 7066 50566 7078 50618
rect 7078 50566 7092 50618
rect 7116 50566 7130 50618
rect 7130 50566 7142 50618
rect 7142 50566 7172 50618
rect 7196 50566 7206 50618
rect 7206 50566 7252 50618
rect 6956 50564 7012 50566
rect 7036 50564 7092 50566
rect 7116 50564 7172 50566
rect 7196 50564 7252 50566
rect 6956 49530 7012 49532
rect 7036 49530 7092 49532
rect 7116 49530 7172 49532
rect 7196 49530 7252 49532
rect 6956 49478 7002 49530
rect 7002 49478 7012 49530
rect 7036 49478 7066 49530
rect 7066 49478 7078 49530
rect 7078 49478 7092 49530
rect 7116 49478 7130 49530
rect 7130 49478 7142 49530
rect 7142 49478 7172 49530
rect 7196 49478 7206 49530
rect 7206 49478 7252 49530
rect 6956 49476 7012 49478
rect 7036 49476 7092 49478
rect 7116 49476 7172 49478
rect 7196 49476 7252 49478
rect 6956 48442 7012 48444
rect 7036 48442 7092 48444
rect 7116 48442 7172 48444
rect 7196 48442 7252 48444
rect 6956 48390 7002 48442
rect 7002 48390 7012 48442
rect 7036 48390 7066 48442
rect 7066 48390 7078 48442
rect 7078 48390 7092 48442
rect 7116 48390 7130 48442
rect 7130 48390 7142 48442
rect 7142 48390 7172 48442
rect 7196 48390 7206 48442
rect 7206 48390 7252 48442
rect 6956 48388 7012 48390
rect 7036 48388 7092 48390
rect 7116 48388 7172 48390
rect 7196 48388 7252 48390
rect 6956 47354 7012 47356
rect 7036 47354 7092 47356
rect 7116 47354 7172 47356
rect 7196 47354 7252 47356
rect 6956 47302 7002 47354
rect 7002 47302 7012 47354
rect 7036 47302 7066 47354
rect 7066 47302 7078 47354
rect 7078 47302 7092 47354
rect 7116 47302 7130 47354
rect 7130 47302 7142 47354
rect 7142 47302 7172 47354
rect 7196 47302 7206 47354
rect 7206 47302 7252 47354
rect 6956 47300 7012 47302
rect 7036 47300 7092 47302
rect 7116 47300 7172 47302
rect 7196 47300 7252 47302
rect 6956 46266 7012 46268
rect 7036 46266 7092 46268
rect 7116 46266 7172 46268
rect 7196 46266 7252 46268
rect 6956 46214 7002 46266
rect 7002 46214 7012 46266
rect 7036 46214 7066 46266
rect 7066 46214 7078 46266
rect 7078 46214 7092 46266
rect 7116 46214 7130 46266
rect 7130 46214 7142 46266
rect 7142 46214 7172 46266
rect 7196 46214 7206 46266
rect 7206 46214 7252 46266
rect 6956 46212 7012 46214
rect 7036 46212 7092 46214
rect 7116 46212 7172 46214
rect 7196 46212 7252 46214
rect 6956 45178 7012 45180
rect 7036 45178 7092 45180
rect 7116 45178 7172 45180
rect 7196 45178 7252 45180
rect 6956 45126 7002 45178
rect 7002 45126 7012 45178
rect 7036 45126 7066 45178
rect 7066 45126 7078 45178
rect 7078 45126 7092 45178
rect 7116 45126 7130 45178
rect 7130 45126 7142 45178
rect 7142 45126 7172 45178
rect 7196 45126 7206 45178
rect 7206 45126 7252 45178
rect 6956 45124 7012 45126
rect 7036 45124 7092 45126
rect 7116 45124 7172 45126
rect 7196 45124 7252 45126
rect 6956 44090 7012 44092
rect 7036 44090 7092 44092
rect 7116 44090 7172 44092
rect 7196 44090 7252 44092
rect 6956 44038 7002 44090
rect 7002 44038 7012 44090
rect 7036 44038 7066 44090
rect 7066 44038 7078 44090
rect 7078 44038 7092 44090
rect 7116 44038 7130 44090
rect 7130 44038 7142 44090
rect 7142 44038 7172 44090
rect 7196 44038 7206 44090
rect 7206 44038 7252 44090
rect 6956 44036 7012 44038
rect 7036 44036 7092 44038
rect 7116 44036 7172 44038
rect 7196 44036 7252 44038
rect 6956 43002 7012 43004
rect 7036 43002 7092 43004
rect 7116 43002 7172 43004
rect 7196 43002 7252 43004
rect 6956 42950 7002 43002
rect 7002 42950 7012 43002
rect 7036 42950 7066 43002
rect 7066 42950 7078 43002
rect 7078 42950 7092 43002
rect 7116 42950 7130 43002
rect 7130 42950 7142 43002
rect 7142 42950 7172 43002
rect 7196 42950 7206 43002
rect 7206 42950 7252 43002
rect 6956 42948 7012 42950
rect 7036 42948 7092 42950
rect 7116 42948 7172 42950
rect 7196 42948 7252 42950
rect 6956 41914 7012 41916
rect 7036 41914 7092 41916
rect 7116 41914 7172 41916
rect 7196 41914 7252 41916
rect 6956 41862 7002 41914
rect 7002 41862 7012 41914
rect 7036 41862 7066 41914
rect 7066 41862 7078 41914
rect 7078 41862 7092 41914
rect 7116 41862 7130 41914
rect 7130 41862 7142 41914
rect 7142 41862 7172 41914
rect 7196 41862 7206 41914
rect 7206 41862 7252 41914
rect 6956 41860 7012 41862
rect 7036 41860 7092 41862
rect 7116 41860 7172 41862
rect 7196 41860 7252 41862
rect 6956 40826 7012 40828
rect 7036 40826 7092 40828
rect 7116 40826 7172 40828
rect 7196 40826 7252 40828
rect 6956 40774 7002 40826
rect 7002 40774 7012 40826
rect 7036 40774 7066 40826
rect 7066 40774 7078 40826
rect 7078 40774 7092 40826
rect 7116 40774 7130 40826
rect 7130 40774 7142 40826
rect 7142 40774 7172 40826
rect 7196 40774 7206 40826
rect 7206 40774 7252 40826
rect 6956 40772 7012 40774
rect 7036 40772 7092 40774
rect 7116 40772 7172 40774
rect 7196 40772 7252 40774
rect 6956 39738 7012 39740
rect 7036 39738 7092 39740
rect 7116 39738 7172 39740
rect 7196 39738 7252 39740
rect 6956 39686 7002 39738
rect 7002 39686 7012 39738
rect 7036 39686 7066 39738
rect 7066 39686 7078 39738
rect 7078 39686 7092 39738
rect 7116 39686 7130 39738
rect 7130 39686 7142 39738
rect 7142 39686 7172 39738
rect 7196 39686 7206 39738
rect 7206 39686 7252 39738
rect 6956 39684 7012 39686
rect 7036 39684 7092 39686
rect 7116 39684 7172 39686
rect 7196 39684 7252 39686
rect 6956 38650 7012 38652
rect 7036 38650 7092 38652
rect 7116 38650 7172 38652
rect 7196 38650 7252 38652
rect 6956 38598 7002 38650
rect 7002 38598 7012 38650
rect 7036 38598 7066 38650
rect 7066 38598 7078 38650
rect 7078 38598 7092 38650
rect 7116 38598 7130 38650
rect 7130 38598 7142 38650
rect 7142 38598 7172 38650
rect 7196 38598 7206 38650
rect 7206 38598 7252 38650
rect 6956 38596 7012 38598
rect 7036 38596 7092 38598
rect 7116 38596 7172 38598
rect 7196 38596 7252 38598
rect 6956 37562 7012 37564
rect 7036 37562 7092 37564
rect 7116 37562 7172 37564
rect 7196 37562 7252 37564
rect 6956 37510 7002 37562
rect 7002 37510 7012 37562
rect 7036 37510 7066 37562
rect 7066 37510 7078 37562
rect 7078 37510 7092 37562
rect 7116 37510 7130 37562
rect 7130 37510 7142 37562
rect 7142 37510 7172 37562
rect 7196 37510 7206 37562
rect 7206 37510 7252 37562
rect 6956 37508 7012 37510
rect 7036 37508 7092 37510
rect 7116 37508 7172 37510
rect 7196 37508 7252 37510
rect 6956 36474 7012 36476
rect 7036 36474 7092 36476
rect 7116 36474 7172 36476
rect 7196 36474 7252 36476
rect 6956 36422 7002 36474
rect 7002 36422 7012 36474
rect 7036 36422 7066 36474
rect 7066 36422 7078 36474
rect 7078 36422 7092 36474
rect 7116 36422 7130 36474
rect 7130 36422 7142 36474
rect 7142 36422 7172 36474
rect 7196 36422 7206 36474
rect 7206 36422 7252 36474
rect 6956 36420 7012 36422
rect 7036 36420 7092 36422
rect 7116 36420 7172 36422
rect 7196 36420 7252 36422
rect 6956 35386 7012 35388
rect 7036 35386 7092 35388
rect 7116 35386 7172 35388
rect 7196 35386 7252 35388
rect 6956 35334 7002 35386
rect 7002 35334 7012 35386
rect 7036 35334 7066 35386
rect 7066 35334 7078 35386
rect 7078 35334 7092 35386
rect 7116 35334 7130 35386
rect 7130 35334 7142 35386
rect 7142 35334 7172 35386
rect 7196 35334 7206 35386
rect 7206 35334 7252 35386
rect 6956 35332 7012 35334
rect 7036 35332 7092 35334
rect 7116 35332 7172 35334
rect 7196 35332 7252 35334
rect 6956 34298 7012 34300
rect 7036 34298 7092 34300
rect 7116 34298 7172 34300
rect 7196 34298 7252 34300
rect 6956 34246 7002 34298
rect 7002 34246 7012 34298
rect 7036 34246 7066 34298
rect 7066 34246 7078 34298
rect 7078 34246 7092 34298
rect 7116 34246 7130 34298
rect 7130 34246 7142 34298
rect 7142 34246 7172 34298
rect 7196 34246 7206 34298
rect 7206 34246 7252 34298
rect 6956 34244 7012 34246
rect 7036 34244 7092 34246
rect 7116 34244 7172 34246
rect 7196 34244 7252 34246
rect 6956 33210 7012 33212
rect 7036 33210 7092 33212
rect 7116 33210 7172 33212
rect 7196 33210 7252 33212
rect 6956 33158 7002 33210
rect 7002 33158 7012 33210
rect 7036 33158 7066 33210
rect 7066 33158 7078 33210
rect 7078 33158 7092 33210
rect 7116 33158 7130 33210
rect 7130 33158 7142 33210
rect 7142 33158 7172 33210
rect 7196 33158 7206 33210
rect 7206 33158 7252 33210
rect 6956 33156 7012 33158
rect 7036 33156 7092 33158
rect 7116 33156 7172 33158
rect 7196 33156 7252 33158
rect 6956 32122 7012 32124
rect 7036 32122 7092 32124
rect 7116 32122 7172 32124
rect 7196 32122 7252 32124
rect 6956 32070 7002 32122
rect 7002 32070 7012 32122
rect 7036 32070 7066 32122
rect 7066 32070 7078 32122
rect 7078 32070 7092 32122
rect 7116 32070 7130 32122
rect 7130 32070 7142 32122
rect 7142 32070 7172 32122
rect 7196 32070 7206 32122
rect 7206 32070 7252 32122
rect 6956 32068 7012 32070
rect 7036 32068 7092 32070
rect 7116 32068 7172 32070
rect 7196 32068 7252 32070
rect 6956 31034 7012 31036
rect 7036 31034 7092 31036
rect 7116 31034 7172 31036
rect 7196 31034 7252 31036
rect 6956 30982 7002 31034
rect 7002 30982 7012 31034
rect 7036 30982 7066 31034
rect 7066 30982 7078 31034
rect 7078 30982 7092 31034
rect 7116 30982 7130 31034
rect 7130 30982 7142 31034
rect 7142 30982 7172 31034
rect 7196 30982 7206 31034
rect 7206 30982 7252 31034
rect 6956 30980 7012 30982
rect 7036 30980 7092 30982
rect 7116 30980 7172 30982
rect 7196 30980 7252 30982
rect 6956 29946 7012 29948
rect 7036 29946 7092 29948
rect 7116 29946 7172 29948
rect 7196 29946 7252 29948
rect 6956 29894 7002 29946
rect 7002 29894 7012 29946
rect 7036 29894 7066 29946
rect 7066 29894 7078 29946
rect 7078 29894 7092 29946
rect 7116 29894 7130 29946
rect 7130 29894 7142 29946
rect 7142 29894 7172 29946
rect 7196 29894 7206 29946
rect 7206 29894 7252 29946
rect 6956 29892 7012 29894
rect 7036 29892 7092 29894
rect 7116 29892 7172 29894
rect 7196 29892 7252 29894
rect 6956 28858 7012 28860
rect 7036 28858 7092 28860
rect 7116 28858 7172 28860
rect 7196 28858 7252 28860
rect 6956 28806 7002 28858
rect 7002 28806 7012 28858
rect 7036 28806 7066 28858
rect 7066 28806 7078 28858
rect 7078 28806 7092 28858
rect 7116 28806 7130 28858
rect 7130 28806 7142 28858
rect 7142 28806 7172 28858
rect 7196 28806 7206 28858
rect 7206 28806 7252 28858
rect 6956 28804 7012 28806
rect 7036 28804 7092 28806
rect 7116 28804 7172 28806
rect 7196 28804 7252 28806
rect 6956 27770 7012 27772
rect 7036 27770 7092 27772
rect 7116 27770 7172 27772
rect 7196 27770 7252 27772
rect 6956 27718 7002 27770
rect 7002 27718 7012 27770
rect 7036 27718 7066 27770
rect 7066 27718 7078 27770
rect 7078 27718 7092 27770
rect 7116 27718 7130 27770
rect 7130 27718 7142 27770
rect 7142 27718 7172 27770
rect 7196 27718 7206 27770
rect 7206 27718 7252 27770
rect 6956 27716 7012 27718
rect 7036 27716 7092 27718
rect 7116 27716 7172 27718
rect 7196 27716 7252 27718
rect 6956 26682 7012 26684
rect 7036 26682 7092 26684
rect 7116 26682 7172 26684
rect 7196 26682 7252 26684
rect 6956 26630 7002 26682
rect 7002 26630 7012 26682
rect 7036 26630 7066 26682
rect 7066 26630 7078 26682
rect 7078 26630 7092 26682
rect 7116 26630 7130 26682
rect 7130 26630 7142 26682
rect 7142 26630 7172 26682
rect 7196 26630 7206 26682
rect 7206 26630 7252 26682
rect 6956 26628 7012 26630
rect 7036 26628 7092 26630
rect 7116 26628 7172 26630
rect 7196 26628 7252 26630
rect 6956 25594 7012 25596
rect 7036 25594 7092 25596
rect 7116 25594 7172 25596
rect 7196 25594 7252 25596
rect 6956 25542 7002 25594
rect 7002 25542 7012 25594
rect 7036 25542 7066 25594
rect 7066 25542 7078 25594
rect 7078 25542 7092 25594
rect 7116 25542 7130 25594
rect 7130 25542 7142 25594
rect 7142 25542 7172 25594
rect 7196 25542 7206 25594
rect 7206 25542 7252 25594
rect 6956 25540 7012 25542
rect 7036 25540 7092 25542
rect 7116 25540 7172 25542
rect 7196 25540 7252 25542
rect 6956 24506 7012 24508
rect 7036 24506 7092 24508
rect 7116 24506 7172 24508
rect 7196 24506 7252 24508
rect 6956 24454 7002 24506
rect 7002 24454 7012 24506
rect 7036 24454 7066 24506
rect 7066 24454 7078 24506
rect 7078 24454 7092 24506
rect 7116 24454 7130 24506
rect 7130 24454 7142 24506
rect 7142 24454 7172 24506
rect 7196 24454 7206 24506
rect 7206 24454 7252 24506
rect 6956 24452 7012 24454
rect 7036 24452 7092 24454
rect 7116 24452 7172 24454
rect 7196 24452 7252 24454
rect 6956 23418 7012 23420
rect 7036 23418 7092 23420
rect 7116 23418 7172 23420
rect 7196 23418 7252 23420
rect 6956 23366 7002 23418
rect 7002 23366 7012 23418
rect 7036 23366 7066 23418
rect 7066 23366 7078 23418
rect 7078 23366 7092 23418
rect 7116 23366 7130 23418
rect 7130 23366 7142 23418
rect 7142 23366 7172 23418
rect 7196 23366 7206 23418
rect 7206 23366 7252 23418
rect 6956 23364 7012 23366
rect 7036 23364 7092 23366
rect 7116 23364 7172 23366
rect 7196 23364 7252 23366
rect 7616 67482 7672 67484
rect 7696 67482 7752 67484
rect 7776 67482 7832 67484
rect 7856 67482 7912 67484
rect 7616 67430 7662 67482
rect 7662 67430 7672 67482
rect 7696 67430 7726 67482
rect 7726 67430 7738 67482
rect 7738 67430 7752 67482
rect 7776 67430 7790 67482
rect 7790 67430 7802 67482
rect 7802 67430 7832 67482
rect 7856 67430 7866 67482
rect 7866 67430 7912 67482
rect 7616 67428 7672 67430
rect 7696 67428 7752 67430
rect 7776 67428 7832 67430
rect 7856 67428 7912 67430
rect 7616 66394 7672 66396
rect 7696 66394 7752 66396
rect 7776 66394 7832 66396
rect 7856 66394 7912 66396
rect 7616 66342 7662 66394
rect 7662 66342 7672 66394
rect 7696 66342 7726 66394
rect 7726 66342 7738 66394
rect 7738 66342 7752 66394
rect 7776 66342 7790 66394
rect 7790 66342 7802 66394
rect 7802 66342 7832 66394
rect 7856 66342 7866 66394
rect 7866 66342 7912 66394
rect 7616 66340 7672 66342
rect 7696 66340 7752 66342
rect 7776 66340 7832 66342
rect 7856 66340 7912 66342
rect 7616 65306 7672 65308
rect 7696 65306 7752 65308
rect 7776 65306 7832 65308
rect 7856 65306 7912 65308
rect 7616 65254 7662 65306
rect 7662 65254 7672 65306
rect 7696 65254 7726 65306
rect 7726 65254 7738 65306
rect 7738 65254 7752 65306
rect 7776 65254 7790 65306
rect 7790 65254 7802 65306
rect 7802 65254 7832 65306
rect 7856 65254 7866 65306
rect 7866 65254 7912 65306
rect 7616 65252 7672 65254
rect 7696 65252 7752 65254
rect 7776 65252 7832 65254
rect 7856 65252 7912 65254
rect 7616 64218 7672 64220
rect 7696 64218 7752 64220
rect 7776 64218 7832 64220
rect 7856 64218 7912 64220
rect 7616 64166 7662 64218
rect 7662 64166 7672 64218
rect 7696 64166 7726 64218
rect 7726 64166 7738 64218
rect 7738 64166 7752 64218
rect 7776 64166 7790 64218
rect 7790 64166 7802 64218
rect 7802 64166 7832 64218
rect 7856 64166 7866 64218
rect 7866 64166 7912 64218
rect 7616 64164 7672 64166
rect 7696 64164 7752 64166
rect 7776 64164 7832 64166
rect 7856 64164 7912 64166
rect 7616 63130 7672 63132
rect 7696 63130 7752 63132
rect 7776 63130 7832 63132
rect 7856 63130 7912 63132
rect 7616 63078 7662 63130
rect 7662 63078 7672 63130
rect 7696 63078 7726 63130
rect 7726 63078 7738 63130
rect 7738 63078 7752 63130
rect 7776 63078 7790 63130
rect 7790 63078 7802 63130
rect 7802 63078 7832 63130
rect 7856 63078 7866 63130
rect 7866 63078 7912 63130
rect 7616 63076 7672 63078
rect 7696 63076 7752 63078
rect 7776 63076 7832 63078
rect 7856 63076 7912 63078
rect 7616 62042 7672 62044
rect 7696 62042 7752 62044
rect 7776 62042 7832 62044
rect 7856 62042 7912 62044
rect 7616 61990 7662 62042
rect 7662 61990 7672 62042
rect 7696 61990 7726 62042
rect 7726 61990 7738 62042
rect 7738 61990 7752 62042
rect 7776 61990 7790 62042
rect 7790 61990 7802 62042
rect 7802 61990 7832 62042
rect 7856 61990 7866 62042
rect 7866 61990 7912 62042
rect 7616 61988 7672 61990
rect 7696 61988 7752 61990
rect 7776 61988 7832 61990
rect 7856 61988 7912 61990
rect 7616 60954 7672 60956
rect 7696 60954 7752 60956
rect 7776 60954 7832 60956
rect 7856 60954 7912 60956
rect 7616 60902 7662 60954
rect 7662 60902 7672 60954
rect 7696 60902 7726 60954
rect 7726 60902 7738 60954
rect 7738 60902 7752 60954
rect 7776 60902 7790 60954
rect 7790 60902 7802 60954
rect 7802 60902 7832 60954
rect 7856 60902 7866 60954
rect 7866 60902 7912 60954
rect 7616 60900 7672 60902
rect 7696 60900 7752 60902
rect 7776 60900 7832 60902
rect 7856 60900 7912 60902
rect 7616 59866 7672 59868
rect 7696 59866 7752 59868
rect 7776 59866 7832 59868
rect 7856 59866 7912 59868
rect 7616 59814 7662 59866
rect 7662 59814 7672 59866
rect 7696 59814 7726 59866
rect 7726 59814 7738 59866
rect 7738 59814 7752 59866
rect 7776 59814 7790 59866
rect 7790 59814 7802 59866
rect 7802 59814 7832 59866
rect 7856 59814 7866 59866
rect 7866 59814 7912 59866
rect 7616 59812 7672 59814
rect 7696 59812 7752 59814
rect 7776 59812 7832 59814
rect 7856 59812 7912 59814
rect 7616 58778 7672 58780
rect 7696 58778 7752 58780
rect 7776 58778 7832 58780
rect 7856 58778 7912 58780
rect 7616 58726 7662 58778
rect 7662 58726 7672 58778
rect 7696 58726 7726 58778
rect 7726 58726 7738 58778
rect 7738 58726 7752 58778
rect 7776 58726 7790 58778
rect 7790 58726 7802 58778
rect 7802 58726 7832 58778
rect 7856 58726 7866 58778
rect 7866 58726 7912 58778
rect 7616 58724 7672 58726
rect 7696 58724 7752 58726
rect 7776 58724 7832 58726
rect 7856 58724 7912 58726
rect 7616 57690 7672 57692
rect 7696 57690 7752 57692
rect 7776 57690 7832 57692
rect 7856 57690 7912 57692
rect 7616 57638 7662 57690
rect 7662 57638 7672 57690
rect 7696 57638 7726 57690
rect 7726 57638 7738 57690
rect 7738 57638 7752 57690
rect 7776 57638 7790 57690
rect 7790 57638 7802 57690
rect 7802 57638 7832 57690
rect 7856 57638 7866 57690
rect 7866 57638 7912 57690
rect 7616 57636 7672 57638
rect 7696 57636 7752 57638
rect 7776 57636 7832 57638
rect 7856 57636 7912 57638
rect 7616 56602 7672 56604
rect 7696 56602 7752 56604
rect 7776 56602 7832 56604
rect 7856 56602 7912 56604
rect 7616 56550 7662 56602
rect 7662 56550 7672 56602
rect 7696 56550 7726 56602
rect 7726 56550 7738 56602
rect 7738 56550 7752 56602
rect 7776 56550 7790 56602
rect 7790 56550 7802 56602
rect 7802 56550 7832 56602
rect 7856 56550 7866 56602
rect 7866 56550 7912 56602
rect 7616 56548 7672 56550
rect 7696 56548 7752 56550
rect 7776 56548 7832 56550
rect 7856 56548 7912 56550
rect 7616 55514 7672 55516
rect 7696 55514 7752 55516
rect 7776 55514 7832 55516
rect 7856 55514 7912 55516
rect 7616 55462 7662 55514
rect 7662 55462 7672 55514
rect 7696 55462 7726 55514
rect 7726 55462 7738 55514
rect 7738 55462 7752 55514
rect 7776 55462 7790 55514
rect 7790 55462 7802 55514
rect 7802 55462 7832 55514
rect 7856 55462 7866 55514
rect 7866 55462 7912 55514
rect 7616 55460 7672 55462
rect 7696 55460 7752 55462
rect 7776 55460 7832 55462
rect 7856 55460 7912 55462
rect 7616 54426 7672 54428
rect 7696 54426 7752 54428
rect 7776 54426 7832 54428
rect 7856 54426 7912 54428
rect 7616 54374 7662 54426
rect 7662 54374 7672 54426
rect 7696 54374 7726 54426
rect 7726 54374 7738 54426
rect 7738 54374 7752 54426
rect 7776 54374 7790 54426
rect 7790 54374 7802 54426
rect 7802 54374 7832 54426
rect 7856 54374 7866 54426
rect 7866 54374 7912 54426
rect 7616 54372 7672 54374
rect 7696 54372 7752 54374
rect 7776 54372 7832 54374
rect 7856 54372 7912 54374
rect 7616 53338 7672 53340
rect 7696 53338 7752 53340
rect 7776 53338 7832 53340
rect 7856 53338 7912 53340
rect 7616 53286 7662 53338
rect 7662 53286 7672 53338
rect 7696 53286 7726 53338
rect 7726 53286 7738 53338
rect 7738 53286 7752 53338
rect 7776 53286 7790 53338
rect 7790 53286 7802 53338
rect 7802 53286 7832 53338
rect 7856 53286 7866 53338
rect 7866 53286 7912 53338
rect 7616 53284 7672 53286
rect 7696 53284 7752 53286
rect 7776 53284 7832 53286
rect 7856 53284 7912 53286
rect 7616 52250 7672 52252
rect 7696 52250 7752 52252
rect 7776 52250 7832 52252
rect 7856 52250 7912 52252
rect 7616 52198 7662 52250
rect 7662 52198 7672 52250
rect 7696 52198 7726 52250
rect 7726 52198 7738 52250
rect 7738 52198 7752 52250
rect 7776 52198 7790 52250
rect 7790 52198 7802 52250
rect 7802 52198 7832 52250
rect 7856 52198 7866 52250
rect 7866 52198 7912 52250
rect 7616 52196 7672 52198
rect 7696 52196 7752 52198
rect 7776 52196 7832 52198
rect 7856 52196 7912 52198
rect 7616 51162 7672 51164
rect 7696 51162 7752 51164
rect 7776 51162 7832 51164
rect 7856 51162 7912 51164
rect 7616 51110 7662 51162
rect 7662 51110 7672 51162
rect 7696 51110 7726 51162
rect 7726 51110 7738 51162
rect 7738 51110 7752 51162
rect 7776 51110 7790 51162
rect 7790 51110 7802 51162
rect 7802 51110 7832 51162
rect 7856 51110 7866 51162
rect 7866 51110 7912 51162
rect 7616 51108 7672 51110
rect 7696 51108 7752 51110
rect 7776 51108 7832 51110
rect 7856 51108 7912 51110
rect 7616 50074 7672 50076
rect 7696 50074 7752 50076
rect 7776 50074 7832 50076
rect 7856 50074 7912 50076
rect 7616 50022 7662 50074
rect 7662 50022 7672 50074
rect 7696 50022 7726 50074
rect 7726 50022 7738 50074
rect 7738 50022 7752 50074
rect 7776 50022 7790 50074
rect 7790 50022 7802 50074
rect 7802 50022 7832 50074
rect 7856 50022 7866 50074
rect 7866 50022 7912 50074
rect 7616 50020 7672 50022
rect 7696 50020 7752 50022
rect 7776 50020 7832 50022
rect 7856 50020 7912 50022
rect 7616 48986 7672 48988
rect 7696 48986 7752 48988
rect 7776 48986 7832 48988
rect 7856 48986 7912 48988
rect 7616 48934 7662 48986
rect 7662 48934 7672 48986
rect 7696 48934 7726 48986
rect 7726 48934 7738 48986
rect 7738 48934 7752 48986
rect 7776 48934 7790 48986
rect 7790 48934 7802 48986
rect 7802 48934 7832 48986
rect 7856 48934 7866 48986
rect 7866 48934 7912 48986
rect 7616 48932 7672 48934
rect 7696 48932 7752 48934
rect 7776 48932 7832 48934
rect 7856 48932 7912 48934
rect 7616 47898 7672 47900
rect 7696 47898 7752 47900
rect 7776 47898 7832 47900
rect 7856 47898 7912 47900
rect 7616 47846 7662 47898
rect 7662 47846 7672 47898
rect 7696 47846 7726 47898
rect 7726 47846 7738 47898
rect 7738 47846 7752 47898
rect 7776 47846 7790 47898
rect 7790 47846 7802 47898
rect 7802 47846 7832 47898
rect 7856 47846 7866 47898
rect 7866 47846 7912 47898
rect 7616 47844 7672 47846
rect 7696 47844 7752 47846
rect 7776 47844 7832 47846
rect 7856 47844 7912 47846
rect 7616 46810 7672 46812
rect 7696 46810 7752 46812
rect 7776 46810 7832 46812
rect 7856 46810 7912 46812
rect 7616 46758 7662 46810
rect 7662 46758 7672 46810
rect 7696 46758 7726 46810
rect 7726 46758 7738 46810
rect 7738 46758 7752 46810
rect 7776 46758 7790 46810
rect 7790 46758 7802 46810
rect 7802 46758 7832 46810
rect 7856 46758 7866 46810
rect 7866 46758 7912 46810
rect 7616 46756 7672 46758
rect 7696 46756 7752 46758
rect 7776 46756 7832 46758
rect 7856 46756 7912 46758
rect 7616 45722 7672 45724
rect 7696 45722 7752 45724
rect 7776 45722 7832 45724
rect 7856 45722 7912 45724
rect 7616 45670 7662 45722
rect 7662 45670 7672 45722
rect 7696 45670 7726 45722
rect 7726 45670 7738 45722
rect 7738 45670 7752 45722
rect 7776 45670 7790 45722
rect 7790 45670 7802 45722
rect 7802 45670 7832 45722
rect 7856 45670 7866 45722
rect 7866 45670 7912 45722
rect 7616 45668 7672 45670
rect 7696 45668 7752 45670
rect 7776 45668 7832 45670
rect 7856 45668 7912 45670
rect 7616 44634 7672 44636
rect 7696 44634 7752 44636
rect 7776 44634 7832 44636
rect 7856 44634 7912 44636
rect 7616 44582 7662 44634
rect 7662 44582 7672 44634
rect 7696 44582 7726 44634
rect 7726 44582 7738 44634
rect 7738 44582 7752 44634
rect 7776 44582 7790 44634
rect 7790 44582 7802 44634
rect 7802 44582 7832 44634
rect 7856 44582 7866 44634
rect 7866 44582 7912 44634
rect 7616 44580 7672 44582
rect 7696 44580 7752 44582
rect 7776 44580 7832 44582
rect 7856 44580 7912 44582
rect 7616 43546 7672 43548
rect 7696 43546 7752 43548
rect 7776 43546 7832 43548
rect 7856 43546 7912 43548
rect 7616 43494 7662 43546
rect 7662 43494 7672 43546
rect 7696 43494 7726 43546
rect 7726 43494 7738 43546
rect 7738 43494 7752 43546
rect 7776 43494 7790 43546
rect 7790 43494 7802 43546
rect 7802 43494 7832 43546
rect 7856 43494 7866 43546
rect 7866 43494 7912 43546
rect 7616 43492 7672 43494
rect 7696 43492 7752 43494
rect 7776 43492 7832 43494
rect 7856 43492 7912 43494
rect 7616 42458 7672 42460
rect 7696 42458 7752 42460
rect 7776 42458 7832 42460
rect 7856 42458 7912 42460
rect 7616 42406 7662 42458
rect 7662 42406 7672 42458
rect 7696 42406 7726 42458
rect 7726 42406 7738 42458
rect 7738 42406 7752 42458
rect 7776 42406 7790 42458
rect 7790 42406 7802 42458
rect 7802 42406 7832 42458
rect 7856 42406 7866 42458
rect 7866 42406 7912 42458
rect 7616 42404 7672 42406
rect 7696 42404 7752 42406
rect 7776 42404 7832 42406
rect 7856 42404 7912 42406
rect 7616 41370 7672 41372
rect 7696 41370 7752 41372
rect 7776 41370 7832 41372
rect 7856 41370 7912 41372
rect 7616 41318 7662 41370
rect 7662 41318 7672 41370
rect 7696 41318 7726 41370
rect 7726 41318 7738 41370
rect 7738 41318 7752 41370
rect 7776 41318 7790 41370
rect 7790 41318 7802 41370
rect 7802 41318 7832 41370
rect 7856 41318 7866 41370
rect 7866 41318 7912 41370
rect 7616 41316 7672 41318
rect 7696 41316 7752 41318
rect 7776 41316 7832 41318
rect 7856 41316 7912 41318
rect 6918 22616 6974 22672
rect 6956 22330 7012 22332
rect 7036 22330 7092 22332
rect 7116 22330 7172 22332
rect 7196 22330 7252 22332
rect 6956 22278 7002 22330
rect 7002 22278 7012 22330
rect 7036 22278 7066 22330
rect 7066 22278 7078 22330
rect 7078 22278 7092 22330
rect 7116 22278 7130 22330
rect 7130 22278 7142 22330
rect 7142 22278 7172 22330
rect 7196 22278 7206 22330
rect 7206 22278 7252 22330
rect 6956 22276 7012 22278
rect 7036 22276 7092 22278
rect 7116 22276 7172 22278
rect 7196 22276 7252 22278
rect 6956 21242 7012 21244
rect 7036 21242 7092 21244
rect 7116 21242 7172 21244
rect 7196 21242 7252 21244
rect 6956 21190 7002 21242
rect 7002 21190 7012 21242
rect 7036 21190 7066 21242
rect 7066 21190 7078 21242
rect 7078 21190 7092 21242
rect 7116 21190 7130 21242
rect 7130 21190 7142 21242
rect 7142 21190 7172 21242
rect 7196 21190 7206 21242
rect 7206 21190 7252 21242
rect 6956 21188 7012 21190
rect 7036 21188 7092 21190
rect 7116 21188 7172 21190
rect 7196 21188 7252 21190
rect 6956 20154 7012 20156
rect 7036 20154 7092 20156
rect 7116 20154 7172 20156
rect 7196 20154 7252 20156
rect 6956 20102 7002 20154
rect 7002 20102 7012 20154
rect 7036 20102 7066 20154
rect 7066 20102 7078 20154
rect 7078 20102 7092 20154
rect 7116 20102 7130 20154
rect 7130 20102 7142 20154
rect 7142 20102 7172 20154
rect 7196 20102 7206 20154
rect 7206 20102 7252 20154
rect 6956 20100 7012 20102
rect 7036 20100 7092 20102
rect 7116 20100 7172 20102
rect 7196 20100 7252 20102
rect 6956 19066 7012 19068
rect 7036 19066 7092 19068
rect 7116 19066 7172 19068
rect 7196 19066 7252 19068
rect 6956 19014 7002 19066
rect 7002 19014 7012 19066
rect 7036 19014 7066 19066
rect 7066 19014 7078 19066
rect 7078 19014 7092 19066
rect 7116 19014 7130 19066
rect 7130 19014 7142 19066
rect 7142 19014 7172 19066
rect 7196 19014 7206 19066
rect 7206 19014 7252 19066
rect 6956 19012 7012 19014
rect 7036 19012 7092 19014
rect 7116 19012 7172 19014
rect 7196 19012 7252 19014
rect 6956 17978 7012 17980
rect 7036 17978 7092 17980
rect 7116 17978 7172 17980
rect 7196 17978 7252 17980
rect 6956 17926 7002 17978
rect 7002 17926 7012 17978
rect 7036 17926 7066 17978
rect 7066 17926 7078 17978
rect 7078 17926 7092 17978
rect 7116 17926 7130 17978
rect 7130 17926 7142 17978
rect 7142 17926 7172 17978
rect 7196 17926 7206 17978
rect 7206 17926 7252 17978
rect 6956 17924 7012 17926
rect 7036 17924 7092 17926
rect 7116 17924 7172 17926
rect 7196 17924 7252 17926
rect 6956 16890 7012 16892
rect 7036 16890 7092 16892
rect 7116 16890 7172 16892
rect 7196 16890 7252 16892
rect 6956 16838 7002 16890
rect 7002 16838 7012 16890
rect 7036 16838 7066 16890
rect 7066 16838 7078 16890
rect 7078 16838 7092 16890
rect 7116 16838 7130 16890
rect 7130 16838 7142 16890
rect 7142 16838 7172 16890
rect 7196 16838 7206 16890
rect 7206 16838 7252 16890
rect 6956 16836 7012 16838
rect 7036 16836 7092 16838
rect 7116 16836 7172 16838
rect 7196 16836 7252 16838
rect 6956 15802 7012 15804
rect 7036 15802 7092 15804
rect 7116 15802 7172 15804
rect 7196 15802 7252 15804
rect 6956 15750 7002 15802
rect 7002 15750 7012 15802
rect 7036 15750 7066 15802
rect 7066 15750 7078 15802
rect 7078 15750 7092 15802
rect 7116 15750 7130 15802
rect 7130 15750 7142 15802
rect 7142 15750 7172 15802
rect 7196 15750 7206 15802
rect 7206 15750 7252 15802
rect 6956 15748 7012 15750
rect 7036 15748 7092 15750
rect 7116 15748 7172 15750
rect 7196 15748 7252 15750
rect 6956 14714 7012 14716
rect 7036 14714 7092 14716
rect 7116 14714 7172 14716
rect 7196 14714 7252 14716
rect 6956 14662 7002 14714
rect 7002 14662 7012 14714
rect 7036 14662 7066 14714
rect 7066 14662 7078 14714
rect 7078 14662 7092 14714
rect 7116 14662 7130 14714
rect 7130 14662 7142 14714
rect 7142 14662 7172 14714
rect 7196 14662 7206 14714
rect 7206 14662 7252 14714
rect 6956 14660 7012 14662
rect 7036 14660 7092 14662
rect 7116 14660 7172 14662
rect 7196 14660 7252 14662
rect 6956 13626 7012 13628
rect 7036 13626 7092 13628
rect 7116 13626 7172 13628
rect 7196 13626 7252 13628
rect 6956 13574 7002 13626
rect 7002 13574 7012 13626
rect 7036 13574 7066 13626
rect 7066 13574 7078 13626
rect 7078 13574 7092 13626
rect 7116 13574 7130 13626
rect 7130 13574 7142 13626
rect 7142 13574 7172 13626
rect 7196 13574 7206 13626
rect 7206 13574 7252 13626
rect 6956 13572 7012 13574
rect 7036 13572 7092 13574
rect 7116 13572 7172 13574
rect 7196 13572 7252 13574
rect 6956 12538 7012 12540
rect 7036 12538 7092 12540
rect 7116 12538 7172 12540
rect 7196 12538 7252 12540
rect 6956 12486 7002 12538
rect 7002 12486 7012 12538
rect 7036 12486 7066 12538
rect 7066 12486 7078 12538
rect 7078 12486 7092 12538
rect 7116 12486 7130 12538
rect 7130 12486 7142 12538
rect 7142 12486 7172 12538
rect 7196 12486 7206 12538
rect 7206 12486 7252 12538
rect 6956 12484 7012 12486
rect 7036 12484 7092 12486
rect 7116 12484 7172 12486
rect 7196 12484 7252 12486
rect 6956 11450 7012 11452
rect 7036 11450 7092 11452
rect 7116 11450 7172 11452
rect 7196 11450 7252 11452
rect 6956 11398 7002 11450
rect 7002 11398 7012 11450
rect 7036 11398 7066 11450
rect 7066 11398 7078 11450
rect 7078 11398 7092 11450
rect 7116 11398 7130 11450
rect 7130 11398 7142 11450
rect 7142 11398 7172 11450
rect 7196 11398 7206 11450
rect 7206 11398 7252 11450
rect 6956 11396 7012 11398
rect 7036 11396 7092 11398
rect 7116 11396 7172 11398
rect 7196 11396 7252 11398
rect 6956 10362 7012 10364
rect 7036 10362 7092 10364
rect 7116 10362 7172 10364
rect 7196 10362 7252 10364
rect 6956 10310 7002 10362
rect 7002 10310 7012 10362
rect 7036 10310 7066 10362
rect 7066 10310 7078 10362
rect 7078 10310 7092 10362
rect 7116 10310 7130 10362
rect 7130 10310 7142 10362
rect 7142 10310 7172 10362
rect 7196 10310 7206 10362
rect 7206 10310 7252 10362
rect 6956 10308 7012 10310
rect 7036 10308 7092 10310
rect 7116 10308 7172 10310
rect 7196 10308 7252 10310
rect 6956 9274 7012 9276
rect 7036 9274 7092 9276
rect 7116 9274 7172 9276
rect 7196 9274 7252 9276
rect 6956 9222 7002 9274
rect 7002 9222 7012 9274
rect 7036 9222 7066 9274
rect 7066 9222 7078 9274
rect 7078 9222 7092 9274
rect 7116 9222 7130 9274
rect 7130 9222 7142 9274
rect 7142 9222 7172 9274
rect 7196 9222 7206 9274
rect 7206 9222 7252 9274
rect 6956 9220 7012 9222
rect 7036 9220 7092 9222
rect 7116 9220 7172 9222
rect 7196 9220 7252 9222
rect 6956 8186 7012 8188
rect 7036 8186 7092 8188
rect 7116 8186 7172 8188
rect 7196 8186 7252 8188
rect 6956 8134 7002 8186
rect 7002 8134 7012 8186
rect 7036 8134 7066 8186
rect 7066 8134 7078 8186
rect 7078 8134 7092 8186
rect 7116 8134 7130 8186
rect 7130 8134 7142 8186
rect 7142 8134 7172 8186
rect 7196 8134 7206 8186
rect 7206 8134 7252 8186
rect 6956 8132 7012 8134
rect 7036 8132 7092 8134
rect 7116 8132 7172 8134
rect 7196 8132 7252 8134
rect 6956 7098 7012 7100
rect 7036 7098 7092 7100
rect 7116 7098 7172 7100
rect 7196 7098 7252 7100
rect 6956 7046 7002 7098
rect 7002 7046 7012 7098
rect 7036 7046 7066 7098
rect 7066 7046 7078 7098
rect 7078 7046 7092 7098
rect 7116 7046 7130 7098
rect 7130 7046 7142 7098
rect 7142 7046 7172 7098
rect 7196 7046 7206 7098
rect 7206 7046 7252 7098
rect 6956 7044 7012 7046
rect 7036 7044 7092 7046
rect 7116 7044 7172 7046
rect 7196 7044 7252 7046
rect 6956 6010 7012 6012
rect 7036 6010 7092 6012
rect 7116 6010 7172 6012
rect 7196 6010 7252 6012
rect 6956 5958 7002 6010
rect 7002 5958 7012 6010
rect 7036 5958 7066 6010
rect 7066 5958 7078 6010
rect 7078 5958 7092 6010
rect 7116 5958 7130 6010
rect 7130 5958 7142 6010
rect 7142 5958 7172 6010
rect 7196 5958 7206 6010
rect 7206 5958 7252 6010
rect 6956 5956 7012 5958
rect 7036 5956 7092 5958
rect 7116 5956 7172 5958
rect 7196 5956 7252 5958
rect 6956 4922 7012 4924
rect 7036 4922 7092 4924
rect 7116 4922 7172 4924
rect 7196 4922 7252 4924
rect 6956 4870 7002 4922
rect 7002 4870 7012 4922
rect 7036 4870 7066 4922
rect 7066 4870 7078 4922
rect 7078 4870 7092 4922
rect 7116 4870 7130 4922
rect 7130 4870 7142 4922
rect 7142 4870 7172 4922
rect 7196 4870 7206 4922
rect 7206 4870 7252 4922
rect 6956 4868 7012 4870
rect 7036 4868 7092 4870
rect 7116 4868 7172 4870
rect 7196 4868 7252 4870
rect 6956 3834 7012 3836
rect 7036 3834 7092 3836
rect 7116 3834 7172 3836
rect 7196 3834 7252 3836
rect 6956 3782 7002 3834
rect 7002 3782 7012 3834
rect 7036 3782 7066 3834
rect 7066 3782 7078 3834
rect 7078 3782 7092 3834
rect 7116 3782 7130 3834
rect 7130 3782 7142 3834
rect 7142 3782 7172 3834
rect 7196 3782 7206 3834
rect 7206 3782 7252 3834
rect 6956 3780 7012 3782
rect 7036 3780 7092 3782
rect 7116 3780 7172 3782
rect 7196 3780 7252 3782
rect 7616 40282 7672 40284
rect 7696 40282 7752 40284
rect 7776 40282 7832 40284
rect 7856 40282 7912 40284
rect 7616 40230 7662 40282
rect 7662 40230 7672 40282
rect 7696 40230 7726 40282
rect 7726 40230 7738 40282
rect 7738 40230 7752 40282
rect 7776 40230 7790 40282
rect 7790 40230 7802 40282
rect 7802 40230 7832 40282
rect 7856 40230 7866 40282
rect 7866 40230 7912 40282
rect 7616 40228 7672 40230
rect 7696 40228 7752 40230
rect 7776 40228 7832 40230
rect 7856 40228 7912 40230
rect 7616 39194 7672 39196
rect 7696 39194 7752 39196
rect 7776 39194 7832 39196
rect 7856 39194 7912 39196
rect 7616 39142 7662 39194
rect 7662 39142 7672 39194
rect 7696 39142 7726 39194
rect 7726 39142 7738 39194
rect 7738 39142 7752 39194
rect 7776 39142 7790 39194
rect 7790 39142 7802 39194
rect 7802 39142 7832 39194
rect 7856 39142 7866 39194
rect 7866 39142 7912 39194
rect 7616 39140 7672 39142
rect 7696 39140 7752 39142
rect 7776 39140 7832 39142
rect 7856 39140 7912 39142
rect 7616 38106 7672 38108
rect 7696 38106 7752 38108
rect 7776 38106 7832 38108
rect 7856 38106 7912 38108
rect 7616 38054 7662 38106
rect 7662 38054 7672 38106
rect 7696 38054 7726 38106
rect 7726 38054 7738 38106
rect 7738 38054 7752 38106
rect 7776 38054 7790 38106
rect 7790 38054 7802 38106
rect 7802 38054 7832 38106
rect 7856 38054 7866 38106
rect 7866 38054 7912 38106
rect 7616 38052 7672 38054
rect 7696 38052 7752 38054
rect 7776 38052 7832 38054
rect 7856 38052 7912 38054
rect 7616 37018 7672 37020
rect 7696 37018 7752 37020
rect 7776 37018 7832 37020
rect 7856 37018 7912 37020
rect 7616 36966 7662 37018
rect 7662 36966 7672 37018
rect 7696 36966 7726 37018
rect 7726 36966 7738 37018
rect 7738 36966 7752 37018
rect 7776 36966 7790 37018
rect 7790 36966 7802 37018
rect 7802 36966 7832 37018
rect 7856 36966 7866 37018
rect 7866 36966 7912 37018
rect 7616 36964 7672 36966
rect 7696 36964 7752 36966
rect 7776 36964 7832 36966
rect 7856 36964 7912 36966
rect 7616 35930 7672 35932
rect 7696 35930 7752 35932
rect 7776 35930 7832 35932
rect 7856 35930 7912 35932
rect 7616 35878 7662 35930
rect 7662 35878 7672 35930
rect 7696 35878 7726 35930
rect 7726 35878 7738 35930
rect 7738 35878 7752 35930
rect 7776 35878 7790 35930
rect 7790 35878 7802 35930
rect 7802 35878 7832 35930
rect 7856 35878 7866 35930
rect 7866 35878 7912 35930
rect 7616 35876 7672 35878
rect 7696 35876 7752 35878
rect 7776 35876 7832 35878
rect 7856 35876 7912 35878
rect 7616 34842 7672 34844
rect 7696 34842 7752 34844
rect 7776 34842 7832 34844
rect 7856 34842 7912 34844
rect 7616 34790 7662 34842
rect 7662 34790 7672 34842
rect 7696 34790 7726 34842
rect 7726 34790 7738 34842
rect 7738 34790 7752 34842
rect 7776 34790 7790 34842
rect 7790 34790 7802 34842
rect 7802 34790 7832 34842
rect 7856 34790 7866 34842
rect 7866 34790 7912 34842
rect 7616 34788 7672 34790
rect 7696 34788 7752 34790
rect 7776 34788 7832 34790
rect 7856 34788 7912 34790
rect 7616 33754 7672 33756
rect 7696 33754 7752 33756
rect 7776 33754 7832 33756
rect 7856 33754 7912 33756
rect 7616 33702 7662 33754
rect 7662 33702 7672 33754
rect 7696 33702 7726 33754
rect 7726 33702 7738 33754
rect 7738 33702 7752 33754
rect 7776 33702 7790 33754
rect 7790 33702 7802 33754
rect 7802 33702 7832 33754
rect 7856 33702 7866 33754
rect 7866 33702 7912 33754
rect 7616 33700 7672 33702
rect 7696 33700 7752 33702
rect 7776 33700 7832 33702
rect 7856 33700 7912 33702
rect 7616 32666 7672 32668
rect 7696 32666 7752 32668
rect 7776 32666 7832 32668
rect 7856 32666 7912 32668
rect 7616 32614 7662 32666
rect 7662 32614 7672 32666
rect 7696 32614 7726 32666
rect 7726 32614 7738 32666
rect 7738 32614 7752 32666
rect 7776 32614 7790 32666
rect 7790 32614 7802 32666
rect 7802 32614 7832 32666
rect 7856 32614 7866 32666
rect 7866 32614 7912 32666
rect 7616 32612 7672 32614
rect 7696 32612 7752 32614
rect 7776 32612 7832 32614
rect 7856 32612 7912 32614
rect 7616 31578 7672 31580
rect 7696 31578 7752 31580
rect 7776 31578 7832 31580
rect 7856 31578 7912 31580
rect 7616 31526 7662 31578
rect 7662 31526 7672 31578
rect 7696 31526 7726 31578
rect 7726 31526 7738 31578
rect 7738 31526 7752 31578
rect 7776 31526 7790 31578
rect 7790 31526 7802 31578
rect 7802 31526 7832 31578
rect 7856 31526 7866 31578
rect 7866 31526 7912 31578
rect 7616 31524 7672 31526
rect 7696 31524 7752 31526
rect 7776 31524 7832 31526
rect 7856 31524 7912 31526
rect 7616 30490 7672 30492
rect 7696 30490 7752 30492
rect 7776 30490 7832 30492
rect 7856 30490 7912 30492
rect 7616 30438 7662 30490
rect 7662 30438 7672 30490
rect 7696 30438 7726 30490
rect 7726 30438 7738 30490
rect 7738 30438 7752 30490
rect 7776 30438 7790 30490
rect 7790 30438 7802 30490
rect 7802 30438 7832 30490
rect 7856 30438 7866 30490
rect 7866 30438 7912 30490
rect 7616 30436 7672 30438
rect 7696 30436 7752 30438
rect 7776 30436 7832 30438
rect 7856 30436 7912 30438
rect 7616 29402 7672 29404
rect 7696 29402 7752 29404
rect 7776 29402 7832 29404
rect 7856 29402 7912 29404
rect 7616 29350 7662 29402
rect 7662 29350 7672 29402
rect 7696 29350 7726 29402
rect 7726 29350 7738 29402
rect 7738 29350 7752 29402
rect 7776 29350 7790 29402
rect 7790 29350 7802 29402
rect 7802 29350 7832 29402
rect 7856 29350 7866 29402
rect 7866 29350 7912 29402
rect 7616 29348 7672 29350
rect 7696 29348 7752 29350
rect 7776 29348 7832 29350
rect 7856 29348 7912 29350
rect 7616 28314 7672 28316
rect 7696 28314 7752 28316
rect 7776 28314 7832 28316
rect 7856 28314 7912 28316
rect 7616 28262 7662 28314
rect 7662 28262 7672 28314
rect 7696 28262 7726 28314
rect 7726 28262 7738 28314
rect 7738 28262 7752 28314
rect 7776 28262 7790 28314
rect 7790 28262 7802 28314
rect 7802 28262 7832 28314
rect 7856 28262 7866 28314
rect 7866 28262 7912 28314
rect 7616 28260 7672 28262
rect 7696 28260 7752 28262
rect 7776 28260 7832 28262
rect 7856 28260 7912 28262
rect 7616 27226 7672 27228
rect 7696 27226 7752 27228
rect 7776 27226 7832 27228
rect 7856 27226 7912 27228
rect 7616 27174 7662 27226
rect 7662 27174 7672 27226
rect 7696 27174 7726 27226
rect 7726 27174 7738 27226
rect 7738 27174 7752 27226
rect 7776 27174 7790 27226
rect 7790 27174 7802 27226
rect 7802 27174 7832 27226
rect 7856 27174 7866 27226
rect 7866 27174 7912 27226
rect 7616 27172 7672 27174
rect 7696 27172 7752 27174
rect 7776 27172 7832 27174
rect 7856 27172 7912 27174
rect 7616 26138 7672 26140
rect 7696 26138 7752 26140
rect 7776 26138 7832 26140
rect 7856 26138 7912 26140
rect 7616 26086 7662 26138
rect 7662 26086 7672 26138
rect 7696 26086 7726 26138
rect 7726 26086 7738 26138
rect 7738 26086 7752 26138
rect 7776 26086 7790 26138
rect 7790 26086 7802 26138
rect 7802 26086 7832 26138
rect 7856 26086 7866 26138
rect 7866 26086 7912 26138
rect 7616 26084 7672 26086
rect 7696 26084 7752 26086
rect 7776 26084 7832 26086
rect 7856 26084 7912 26086
rect 7616 25050 7672 25052
rect 7696 25050 7752 25052
rect 7776 25050 7832 25052
rect 7856 25050 7912 25052
rect 7616 24998 7662 25050
rect 7662 24998 7672 25050
rect 7696 24998 7726 25050
rect 7726 24998 7738 25050
rect 7738 24998 7752 25050
rect 7776 24998 7790 25050
rect 7790 24998 7802 25050
rect 7802 24998 7832 25050
rect 7856 24998 7866 25050
rect 7866 24998 7912 25050
rect 7616 24996 7672 24998
rect 7696 24996 7752 24998
rect 7776 24996 7832 24998
rect 7856 24996 7912 24998
rect 7616 23962 7672 23964
rect 7696 23962 7752 23964
rect 7776 23962 7832 23964
rect 7856 23962 7912 23964
rect 7616 23910 7662 23962
rect 7662 23910 7672 23962
rect 7696 23910 7726 23962
rect 7726 23910 7738 23962
rect 7738 23910 7752 23962
rect 7776 23910 7790 23962
rect 7790 23910 7802 23962
rect 7802 23910 7832 23962
rect 7856 23910 7866 23962
rect 7866 23910 7912 23962
rect 7616 23908 7672 23910
rect 7696 23908 7752 23910
rect 7776 23908 7832 23910
rect 7856 23908 7912 23910
rect 7616 22874 7672 22876
rect 7696 22874 7752 22876
rect 7776 22874 7832 22876
rect 7856 22874 7912 22876
rect 7616 22822 7662 22874
rect 7662 22822 7672 22874
rect 7696 22822 7726 22874
rect 7726 22822 7738 22874
rect 7738 22822 7752 22874
rect 7776 22822 7790 22874
rect 7790 22822 7802 22874
rect 7802 22822 7832 22874
rect 7856 22822 7866 22874
rect 7866 22822 7912 22874
rect 7616 22820 7672 22822
rect 7696 22820 7752 22822
rect 7776 22820 7832 22822
rect 7856 22820 7912 22822
rect 7616 21786 7672 21788
rect 7696 21786 7752 21788
rect 7776 21786 7832 21788
rect 7856 21786 7912 21788
rect 7616 21734 7662 21786
rect 7662 21734 7672 21786
rect 7696 21734 7726 21786
rect 7726 21734 7738 21786
rect 7738 21734 7752 21786
rect 7776 21734 7790 21786
rect 7790 21734 7802 21786
rect 7802 21734 7832 21786
rect 7856 21734 7866 21786
rect 7866 21734 7912 21786
rect 7616 21732 7672 21734
rect 7696 21732 7752 21734
rect 7776 21732 7832 21734
rect 7856 21732 7912 21734
rect 7616 20698 7672 20700
rect 7696 20698 7752 20700
rect 7776 20698 7832 20700
rect 7856 20698 7912 20700
rect 7616 20646 7662 20698
rect 7662 20646 7672 20698
rect 7696 20646 7726 20698
rect 7726 20646 7738 20698
rect 7738 20646 7752 20698
rect 7776 20646 7790 20698
rect 7790 20646 7802 20698
rect 7802 20646 7832 20698
rect 7856 20646 7866 20698
rect 7866 20646 7912 20698
rect 7616 20644 7672 20646
rect 7696 20644 7752 20646
rect 7776 20644 7832 20646
rect 7856 20644 7912 20646
rect 7616 19610 7672 19612
rect 7696 19610 7752 19612
rect 7776 19610 7832 19612
rect 7856 19610 7912 19612
rect 7616 19558 7662 19610
rect 7662 19558 7672 19610
rect 7696 19558 7726 19610
rect 7726 19558 7738 19610
rect 7738 19558 7752 19610
rect 7776 19558 7790 19610
rect 7790 19558 7802 19610
rect 7802 19558 7832 19610
rect 7856 19558 7866 19610
rect 7866 19558 7912 19610
rect 7616 19556 7672 19558
rect 7696 19556 7752 19558
rect 7776 19556 7832 19558
rect 7856 19556 7912 19558
rect 7616 18522 7672 18524
rect 7696 18522 7752 18524
rect 7776 18522 7832 18524
rect 7856 18522 7912 18524
rect 7616 18470 7662 18522
rect 7662 18470 7672 18522
rect 7696 18470 7726 18522
rect 7726 18470 7738 18522
rect 7738 18470 7752 18522
rect 7776 18470 7790 18522
rect 7790 18470 7802 18522
rect 7802 18470 7832 18522
rect 7856 18470 7866 18522
rect 7866 18470 7912 18522
rect 7616 18468 7672 18470
rect 7696 18468 7752 18470
rect 7776 18468 7832 18470
rect 7856 18468 7912 18470
rect 7616 17434 7672 17436
rect 7696 17434 7752 17436
rect 7776 17434 7832 17436
rect 7856 17434 7912 17436
rect 7616 17382 7662 17434
rect 7662 17382 7672 17434
rect 7696 17382 7726 17434
rect 7726 17382 7738 17434
rect 7738 17382 7752 17434
rect 7776 17382 7790 17434
rect 7790 17382 7802 17434
rect 7802 17382 7832 17434
rect 7856 17382 7866 17434
rect 7866 17382 7912 17434
rect 7616 17380 7672 17382
rect 7696 17380 7752 17382
rect 7776 17380 7832 17382
rect 7856 17380 7912 17382
rect 7616 16346 7672 16348
rect 7696 16346 7752 16348
rect 7776 16346 7832 16348
rect 7856 16346 7912 16348
rect 7616 16294 7662 16346
rect 7662 16294 7672 16346
rect 7696 16294 7726 16346
rect 7726 16294 7738 16346
rect 7738 16294 7752 16346
rect 7776 16294 7790 16346
rect 7790 16294 7802 16346
rect 7802 16294 7832 16346
rect 7856 16294 7866 16346
rect 7866 16294 7912 16346
rect 7616 16292 7672 16294
rect 7696 16292 7752 16294
rect 7776 16292 7832 16294
rect 7856 16292 7912 16294
rect 7616 15258 7672 15260
rect 7696 15258 7752 15260
rect 7776 15258 7832 15260
rect 7856 15258 7912 15260
rect 7616 15206 7662 15258
rect 7662 15206 7672 15258
rect 7696 15206 7726 15258
rect 7726 15206 7738 15258
rect 7738 15206 7752 15258
rect 7776 15206 7790 15258
rect 7790 15206 7802 15258
rect 7802 15206 7832 15258
rect 7856 15206 7866 15258
rect 7866 15206 7912 15258
rect 7616 15204 7672 15206
rect 7696 15204 7752 15206
rect 7776 15204 7832 15206
rect 7856 15204 7912 15206
rect 7616 14170 7672 14172
rect 7696 14170 7752 14172
rect 7776 14170 7832 14172
rect 7856 14170 7912 14172
rect 7616 14118 7662 14170
rect 7662 14118 7672 14170
rect 7696 14118 7726 14170
rect 7726 14118 7738 14170
rect 7738 14118 7752 14170
rect 7776 14118 7790 14170
rect 7790 14118 7802 14170
rect 7802 14118 7832 14170
rect 7856 14118 7866 14170
rect 7866 14118 7912 14170
rect 7616 14116 7672 14118
rect 7696 14116 7752 14118
rect 7776 14116 7832 14118
rect 7856 14116 7912 14118
rect 7616 13082 7672 13084
rect 7696 13082 7752 13084
rect 7776 13082 7832 13084
rect 7856 13082 7912 13084
rect 7616 13030 7662 13082
rect 7662 13030 7672 13082
rect 7696 13030 7726 13082
rect 7726 13030 7738 13082
rect 7738 13030 7752 13082
rect 7776 13030 7790 13082
rect 7790 13030 7802 13082
rect 7802 13030 7832 13082
rect 7856 13030 7866 13082
rect 7866 13030 7912 13082
rect 7616 13028 7672 13030
rect 7696 13028 7752 13030
rect 7776 13028 7832 13030
rect 7856 13028 7912 13030
rect 7616 11994 7672 11996
rect 7696 11994 7752 11996
rect 7776 11994 7832 11996
rect 7856 11994 7912 11996
rect 7616 11942 7662 11994
rect 7662 11942 7672 11994
rect 7696 11942 7726 11994
rect 7726 11942 7738 11994
rect 7738 11942 7752 11994
rect 7776 11942 7790 11994
rect 7790 11942 7802 11994
rect 7802 11942 7832 11994
rect 7856 11942 7866 11994
rect 7866 11942 7912 11994
rect 7616 11940 7672 11942
rect 7696 11940 7752 11942
rect 7776 11940 7832 11942
rect 7856 11940 7912 11942
rect 7616 10906 7672 10908
rect 7696 10906 7752 10908
rect 7776 10906 7832 10908
rect 7856 10906 7912 10908
rect 7616 10854 7662 10906
rect 7662 10854 7672 10906
rect 7696 10854 7726 10906
rect 7726 10854 7738 10906
rect 7738 10854 7752 10906
rect 7776 10854 7790 10906
rect 7790 10854 7802 10906
rect 7802 10854 7832 10906
rect 7856 10854 7866 10906
rect 7866 10854 7912 10906
rect 7616 10852 7672 10854
rect 7696 10852 7752 10854
rect 7776 10852 7832 10854
rect 7856 10852 7912 10854
rect 7616 9818 7672 9820
rect 7696 9818 7752 9820
rect 7776 9818 7832 9820
rect 7856 9818 7912 9820
rect 7616 9766 7662 9818
rect 7662 9766 7672 9818
rect 7696 9766 7726 9818
rect 7726 9766 7738 9818
rect 7738 9766 7752 9818
rect 7776 9766 7790 9818
rect 7790 9766 7802 9818
rect 7802 9766 7832 9818
rect 7856 9766 7866 9818
rect 7866 9766 7912 9818
rect 7616 9764 7672 9766
rect 7696 9764 7752 9766
rect 7776 9764 7832 9766
rect 7856 9764 7912 9766
rect 7562 9596 7564 9616
rect 7564 9596 7616 9616
rect 7616 9596 7618 9616
rect 7562 9560 7618 9596
rect 7616 8730 7672 8732
rect 7696 8730 7752 8732
rect 7776 8730 7832 8732
rect 7856 8730 7912 8732
rect 7616 8678 7662 8730
rect 7662 8678 7672 8730
rect 7696 8678 7726 8730
rect 7726 8678 7738 8730
rect 7738 8678 7752 8730
rect 7776 8678 7790 8730
rect 7790 8678 7802 8730
rect 7802 8678 7832 8730
rect 7856 8678 7866 8730
rect 7866 8678 7912 8730
rect 7616 8676 7672 8678
rect 7696 8676 7752 8678
rect 7776 8676 7832 8678
rect 7856 8676 7912 8678
rect 7616 7642 7672 7644
rect 7696 7642 7752 7644
rect 7776 7642 7832 7644
rect 7856 7642 7912 7644
rect 7616 7590 7662 7642
rect 7662 7590 7672 7642
rect 7696 7590 7726 7642
rect 7726 7590 7738 7642
rect 7738 7590 7752 7642
rect 7776 7590 7790 7642
rect 7790 7590 7802 7642
rect 7802 7590 7832 7642
rect 7856 7590 7866 7642
rect 7866 7590 7912 7642
rect 7616 7588 7672 7590
rect 7696 7588 7752 7590
rect 7776 7588 7832 7590
rect 7856 7588 7912 7590
rect 7616 6554 7672 6556
rect 7696 6554 7752 6556
rect 7776 6554 7832 6556
rect 7856 6554 7912 6556
rect 7616 6502 7662 6554
rect 7662 6502 7672 6554
rect 7696 6502 7726 6554
rect 7726 6502 7738 6554
rect 7738 6502 7752 6554
rect 7776 6502 7790 6554
rect 7790 6502 7802 6554
rect 7802 6502 7832 6554
rect 7856 6502 7866 6554
rect 7866 6502 7912 6554
rect 7616 6500 7672 6502
rect 7696 6500 7752 6502
rect 7776 6500 7832 6502
rect 7856 6500 7912 6502
rect 7616 5466 7672 5468
rect 7696 5466 7752 5468
rect 7776 5466 7832 5468
rect 7856 5466 7912 5468
rect 7616 5414 7662 5466
rect 7662 5414 7672 5466
rect 7696 5414 7726 5466
rect 7726 5414 7738 5466
rect 7738 5414 7752 5466
rect 7776 5414 7790 5466
rect 7790 5414 7802 5466
rect 7802 5414 7832 5466
rect 7856 5414 7866 5466
rect 7866 5414 7912 5466
rect 7616 5412 7672 5414
rect 7696 5412 7752 5414
rect 7776 5412 7832 5414
rect 7856 5412 7912 5414
rect 7616 4378 7672 4380
rect 7696 4378 7752 4380
rect 7776 4378 7832 4380
rect 7856 4378 7912 4380
rect 7616 4326 7662 4378
rect 7662 4326 7672 4378
rect 7696 4326 7726 4378
rect 7726 4326 7738 4378
rect 7738 4326 7752 4378
rect 7776 4326 7790 4378
rect 7790 4326 7802 4378
rect 7802 4326 7832 4378
rect 7856 4326 7866 4378
rect 7866 4326 7912 4378
rect 7616 4324 7672 4326
rect 7696 4324 7752 4326
rect 7776 4324 7832 4326
rect 7856 4324 7912 4326
rect 7616 3290 7672 3292
rect 7696 3290 7752 3292
rect 7776 3290 7832 3292
rect 7856 3290 7912 3292
rect 7616 3238 7662 3290
rect 7662 3238 7672 3290
rect 7696 3238 7726 3290
rect 7726 3238 7738 3290
rect 7738 3238 7752 3290
rect 7776 3238 7790 3290
rect 7790 3238 7802 3290
rect 7802 3238 7832 3290
rect 7856 3238 7866 3290
rect 7866 3238 7912 3290
rect 7616 3236 7672 3238
rect 7696 3236 7752 3238
rect 7776 3236 7832 3238
rect 7856 3236 7912 3238
rect 11956 69114 12012 69116
rect 12036 69114 12092 69116
rect 12116 69114 12172 69116
rect 12196 69114 12252 69116
rect 11956 69062 12002 69114
rect 12002 69062 12012 69114
rect 12036 69062 12066 69114
rect 12066 69062 12078 69114
rect 12078 69062 12092 69114
rect 12116 69062 12130 69114
rect 12130 69062 12142 69114
rect 12142 69062 12172 69114
rect 12196 69062 12206 69114
rect 12206 69062 12252 69114
rect 11956 69060 12012 69062
rect 12036 69060 12092 69062
rect 12116 69060 12172 69062
rect 12196 69060 12252 69062
rect 12616 68570 12672 68572
rect 12696 68570 12752 68572
rect 12776 68570 12832 68572
rect 12856 68570 12912 68572
rect 12616 68518 12662 68570
rect 12662 68518 12672 68570
rect 12696 68518 12726 68570
rect 12726 68518 12738 68570
rect 12738 68518 12752 68570
rect 12776 68518 12790 68570
rect 12790 68518 12802 68570
rect 12802 68518 12832 68570
rect 12856 68518 12866 68570
rect 12866 68518 12912 68570
rect 12616 68516 12672 68518
rect 12696 68516 12752 68518
rect 12776 68516 12832 68518
rect 12856 68516 12912 68518
rect 9034 30640 9090 30696
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 6956 2746 7012 2748
rect 7036 2746 7092 2748
rect 7116 2746 7172 2748
rect 7196 2746 7252 2748
rect 6956 2694 7002 2746
rect 7002 2694 7012 2746
rect 7036 2694 7066 2746
rect 7066 2694 7078 2746
rect 7078 2694 7092 2746
rect 7116 2694 7130 2746
rect 7130 2694 7142 2746
rect 7142 2694 7172 2746
rect 7196 2694 7206 2746
rect 7206 2694 7252 2746
rect 6956 2692 7012 2694
rect 7036 2692 7092 2694
rect 7116 2692 7172 2694
rect 7196 2692 7252 2694
rect 11956 68026 12012 68028
rect 12036 68026 12092 68028
rect 12116 68026 12172 68028
rect 12196 68026 12252 68028
rect 11956 67974 12002 68026
rect 12002 67974 12012 68026
rect 12036 67974 12066 68026
rect 12066 67974 12078 68026
rect 12078 67974 12092 68026
rect 12116 67974 12130 68026
rect 12130 67974 12142 68026
rect 12142 67974 12172 68026
rect 12196 67974 12206 68026
rect 12206 67974 12252 68026
rect 11956 67972 12012 67974
rect 12036 67972 12092 67974
rect 12116 67972 12172 67974
rect 12196 67972 12252 67974
rect 12616 67482 12672 67484
rect 12696 67482 12752 67484
rect 12776 67482 12832 67484
rect 12856 67482 12912 67484
rect 12616 67430 12662 67482
rect 12662 67430 12672 67482
rect 12696 67430 12726 67482
rect 12726 67430 12738 67482
rect 12738 67430 12752 67482
rect 12776 67430 12790 67482
rect 12790 67430 12802 67482
rect 12802 67430 12832 67482
rect 12856 67430 12866 67482
rect 12866 67430 12912 67482
rect 12616 67428 12672 67430
rect 12696 67428 12752 67430
rect 12776 67428 12832 67430
rect 12856 67428 12912 67430
rect 11956 66938 12012 66940
rect 12036 66938 12092 66940
rect 12116 66938 12172 66940
rect 12196 66938 12252 66940
rect 11956 66886 12002 66938
rect 12002 66886 12012 66938
rect 12036 66886 12066 66938
rect 12066 66886 12078 66938
rect 12078 66886 12092 66938
rect 12116 66886 12130 66938
rect 12130 66886 12142 66938
rect 12142 66886 12172 66938
rect 12196 66886 12206 66938
rect 12206 66886 12252 66938
rect 11956 66884 12012 66886
rect 12036 66884 12092 66886
rect 12116 66884 12172 66886
rect 12196 66884 12252 66886
rect 12616 66394 12672 66396
rect 12696 66394 12752 66396
rect 12776 66394 12832 66396
rect 12856 66394 12912 66396
rect 12616 66342 12662 66394
rect 12662 66342 12672 66394
rect 12696 66342 12726 66394
rect 12726 66342 12738 66394
rect 12738 66342 12752 66394
rect 12776 66342 12790 66394
rect 12790 66342 12802 66394
rect 12802 66342 12832 66394
rect 12856 66342 12866 66394
rect 12866 66342 12912 66394
rect 12616 66340 12672 66342
rect 12696 66340 12752 66342
rect 12776 66340 12832 66342
rect 12856 66340 12912 66342
rect 11956 65850 12012 65852
rect 12036 65850 12092 65852
rect 12116 65850 12172 65852
rect 12196 65850 12252 65852
rect 11956 65798 12002 65850
rect 12002 65798 12012 65850
rect 12036 65798 12066 65850
rect 12066 65798 12078 65850
rect 12078 65798 12092 65850
rect 12116 65798 12130 65850
rect 12130 65798 12142 65850
rect 12142 65798 12172 65850
rect 12196 65798 12206 65850
rect 12206 65798 12252 65850
rect 11956 65796 12012 65798
rect 12036 65796 12092 65798
rect 12116 65796 12172 65798
rect 12196 65796 12252 65798
rect 12616 65306 12672 65308
rect 12696 65306 12752 65308
rect 12776 65306 12832 65308
rect 12856 65306 12912 65308
rect 12616 65254 12662 65306
rect 12662 65254 12672 65306
rect 12696 65254 12726 65306
rect 12726 65254 12738 65306
rect 12738 65254 12752 65306
rect 12776 65254 12790 65306
rect 12790 65254 12802 65306
rect 12802 65254 12832 65306
rect 12856 65254 12866 65306
rect 12866 65254 12912 65306
rect 12616 65252 12672 65254
rect 12696 65252 12752 65254
rect 12776 65252 12832 65254
rect 12856 65252 12912 65254
rect 11956 64762 12012 64764
rect 12036 64762 12092 64764
rect 12116 64762 12172 64764
rect 12196 64762 12252 64764
rect 11956 64710 12002 64762
rect 12002 64710 12012 64762
rect 12036 64710 12066 64762
rect 12066 64710 12078 64762
rect 12078 64710 12092 64762
rect 12116 64710 12130 64762
rect 12130 64710 12142 64762
rect 12142 64710 12172 64762
rect 12196 64710 12206 64762
rect 12206 64710 12252 64762
rect 11956 64708 12012 64710
rect 12036 64708 12092 64710
rect 12116 64708 12172 64710
rect 12196 64708 12252 64710
rect 11956 63674 12012 63676
rect 12036 63674 12092 63676
rect 12116 63674 12172 63676
rect 12196 63674 12252 63676
rect 11956 63622 12002 63674
rect 12002 63622 12012 63674
rect 12036 63622 12066 63674
rect 12066 63622 12078 63674
rect 12078 63622 12092 63674
rect 12116 63622 12130 63674
rect 12130 63622 12142 63674
rect 12142 63622 12172 63674
rect 12196 63622 12206 63674
rect 12206 63622 12252 63674
rect 11956 63620 12012 63622
rect 12036 63620 12092 63622
rect 12116 63620 12172 63622
rect 12196 63620 12252 63622
rect 11956 62586 12012 62588
rect 12036 62586 12092 62588
rect 12116 62586 12172 62588
rect 12196 62586 12252 62588
rect 11956 62534 12002 62586
rect 12002 62534 12012 62586
rect 12036 62534 12066 62586
rect 12066 62534 12078 62586
rect 12078 62534 12092 62586
rect 12116 62534 12130 62586
rect 12130 62534 12142 62586
rect 12142 62534 12172 62586
rect 12196 62534 12206 62586
rect 12206 62534 12252 62586
rect 11956 62532 12012 62534
rect 12036 62532 12092 62534
rect 12116 62532 12172 62534
rect 12196 62532 12252 62534
rect 11956 61498 12012 61500
rect 12036 61498 12092 61500
rect 12116 61498 12172 61500
rect 12196 61498 12252 61500
rect 11956 61446 12002 61498
rect 12002 61446 12012 61498
rect 12036 61446 12066 61498
rect 12066 61446 12078 61498
rect 12078 61446 12092 61498
rect 12116 61446 12130 61498
rect 12130 61446 12142 61498
rect 12142 61446 12172 61498
rect 12196 61446 12206 61498
rect 12206 61446 12252 61498
rect 11956 61444 12012 61446
rect 12036 61444 12092 61446
rect 12116 61444 12172 61446
rect 12196 61444 12252 61446
rect 11956 60410 12012 60412
rect 12036 60410 12092 60412
rect 12116 60410 12172 60412
rect 12196 60410 12252 60412
rect 11956 60358 12002 60410
rect 12002 60358 12012 60410
rect 12036 60358 12066 60410
rect 12066 60358 12078 60410
rect 12078 60358 12092 60410
rect 12116 60358 12130 60410
rect 12130 60358 12142 60410
rect 12142 60358 12172 60410
rect 12196 60358 12206 60410
rect 12206 60358 12252 60410
rect 11956 60356 12012 60358
rect 12036 60356 12092 60358
rect 12116 60356 12172 60358
rect 12196 60356 12252 60358
rect 11956 59322 12012 59324
rect 12036 59322 12092 59324
rect 12116 59322 12172 59324
rect 12196 59322 12252 59324
rect 11956 59270 12002 59322
rect 12002 59270 12012 59322
rect 12036 59270 12066 59322
rect 12066 59270 12078 59322
rect 12078 59270 12092 59322
rect 12116 59270 12130 59322
rect 12130 59270 12142 59322
rect 12142 59270 12172 59322
rect 12196 59270 12206 59322
rect 12206 59270 12252 59322
rect 11956 59268 12012 59270
rect 12036 59268 12092 59270
rect 12116 59268 12172 59270
rect 12196 59268 12252 59270
rect 11956 58234 12012 58236
rect 12036 58234 12092 58236
rect 12116 58234 12172 58236
rect 12196 58234 12252 58236
rect 11956 58182 12002 58234
rect 12002 58182 12012 58234
rect 12036 58182 12066 58234
rect 12066 58182 12078 58234
rect 12078 58182 12092 58234
rect 12116 58182 12130 58234
rect 12130 58182 12142 58234
rect 12142 58182 12172 58234
rect 12196 58182 12206 58234
rect 12206 58182 12252 58234
rect 11956 58180 12012 58182
rect 12036 58180 12092 58182
rect 12116 58180 12172 58182
rect 12196 58180 12252 58182
rect 11956 57146 12012 57148
rect 12036 57146 12092 57148
rect 12116 57146 12172 57148
rect 12196 57146 12252 57148
rect 11956 57094 12002 57146
rect 12002 57094 12012 57146
rect 12036 57094 12066 57146
rect 12066 57094 12078 57146
rect 12078 57094 12092 57146
rect 12116 57094 12130 57146
rect 12130 57094 12142 57146
rect 12142 57094 12172 57146
rect 12196 57094 12206 57146
rect 12206 57094 12252 57146
rect 11956 57092 12012 57094
rect 12036 57092 12092 57094
rect 12116 57092 12172 57094
rect 12196 57092 12252 57094
rect 11956 56058 12012 56060
rect 12036 56058 12092 56060
rect 12116 56058 12172 56060
rect 12196 56058 12252 56060
rect 11956 56006 12002 56058
rect 12002 56006 12012 56058
rect 12036 56006 12066 56058
rect 12066 56006 12078 56058
rect 12078 56006 12092 56058
rect 12116 56006 12130 56058
rect 12130 56006 12142 56058
rect 12142 56006 12172 56058
rect 12196 56006 12206 56058
rect 12206 56006 12252 56058
rect 11956 56004 12012 56006
rect 12036 56004 12092 56006
rect 12116 56004 12172 56006
rect 12196 56004 12252 56006
rect 12616 64218 12672 64220
rect 12696 64218 12752 64220
rect 12776 64218 12832 64220
rect 12856 64218 12912 64220
rect 12616 64166 12662 64218
rect 12662 64166 12672 64218
rect 12696 64166 12726 64218
rect 12726 64166 12738 64218
rect 12738 64166 12752 64218
rect 12776 64166 12790 64218
rect 12790 64166 12802 64218
rect 12802 64166 12832 64218
rect 12856 64166 12866 64218
rect 12866 64166 12912 64218
rect 12616 64164 12672 64166
rect 12696 64164 12752 64166
rect 12776 64164 12832 64166
rect 12856 64164 12912 64166
rect 12616 63130 12672 63132
rect 12696 63130 12752 63132
rect 12776 63130 12832 63132
rect 12856 63130 12912 63132
rect 12616 63078 12662 63130
rect 12662 63078 12672 63130
rect 12696 63078 12726 63130
rect 12726 63078 12738 63130
rect 12738 63078 12752 63130
rect 12776 63078 12790 63130
rect 12790 63078 12802 63130
rect 12802 63078 12832 63130
rect 12856 63078 12866 63130
rect 12866 63078 12912 63130
rect 12616 63076 12672 63078
rect 12696 63076 12752 63078
rect 12776 63076 12832 63078
rect 12856 63076 12912 63078
rect 12616 62042 12672 62044
rect 12696 62042 12752 62044
rect 12776 62042 12832 62044
rect 12856 62042 12912 62044
rect 12616 61990 12662 62042
rect 12662 61990 12672 62042
rect 12696 61990 12726 62042
rect 12726 61990 12738 62042
rect 12738 61990 12752 62042
rect 12776 61990 12790 62042
rect 12790 61990 12802 62042
rect 12802 61990 12832 62042
rect 12856 61990 12866 62042
rect 12866 61990 12912 62042
rect 12616 61988 12672 61990
rect 12696 61988 12752 61990
rect 12776 61988 12832 61990
rect 12856 61988 12912 61990
rect 12616 60954 12672 60956
rect 12696 60954 12752 60956
rect 12776 60954 12832 60956
rect 12856 60954 12912 60956
rect 12616 60902 12662 60954
rect 12662 60902 12672 60954
rect 12696 60902 12726 60954
rect 12726 60902 12738 60954
rect 12738 60902 12752 60954
rect 12776 60902 12790 60954
rect 12790 60902 12802 60954
rect 12802 60902 12832 60954
rect 12856 60902 12866 60954
rect 12866 60902 12912 60954
rect 12616 60900 12672 60902
rect 12696 60900 12752 60902
rect 12776 60900 12832 60902
rect 12856 60900 12912 60902
rect 12616 59866 12672 59868
rect 12696 59866 12752 59868
rect 12776 59866 12832 59868
rect 12856 59866 12912 59868
rect 12616 59814 12662 59866
rect 12662 59814 12672 59866
rect 12696 59814 12726 59866
rect 12726 59814 12738 59866
rect 12738 59814 12752 59866
rect 12776 59814 12790 59866
rect 12790 59814 12802 59866
rect 12802 59814 12832 59866
rect 12856 59814 12866 59866
rect 12866 59814 12912 59866
rect 12616 59812 12672 59814
rect 12696 59812 12752 59814
rect 12776 59812 12832 59814
rect 12856 59812 12912 59814
rect 12616 58778 12672 58780
rect 12696 58778 12752 58780
rect 12776 58778 12832 58780
rect 12856 58778 12912 58780
rect 12616 58726 12662 58778
rect 12662 58726 12672 58778
rect 12696 58726 12726 58778
rect 12726 58726 12738 58778
rect 12738 58726 12752 58778
rect 12776 58726 12790 58778
rect 12790 58726 12802 58778
rect 12802 58726 12832 58778
rect 12856 58726 12866 58778
rect 12866 58726 12912 58778
rect 12616 58724 12672 58726
rect 12696 58724 12752 58726
rect 12776 58724 12832 58726
rect 12856 58724 12912 58726
rect 12616 57690 12672 57692
rect 12696 57690 12752 57692
rect 12776 57690 12832 57692
rect 12856 57690 12912 57692
rect 12616 57638 12662 57690
rect 12662 57638 12672 57690
rect 12696 57638 12726 57690
rect 12726 57638 12738 57690
rect 12738 57638 12752 57690
rect 12776 57638 12790 57690
rect 12790 57638 12802 57690
rect 12802 57638 12832 57690
rect 12856 57638 12866 57690
rect 12866 57638 12912 57690
rect 12616 57636 12672 57638
rect 12696 57636 12752 57638
rect 12776 57636 12832 57638
rect 12856 57636 12912 57638
rect 12616 56602 12672 56604
rect 12696 56602 12752 56604
rect 12776 56602 12832 56604
rect 12856 56602 12912 56604
rect 12616 56550 12662 56602
rect 12662 56550 12672 56602
rect 12696 56550 12726 56602
rect 12726 56550 12738 56602
rect 12738 56550 12752 56602
rect 12776 56550 12790 56602
rect 12790 56550 12802 56602
rect 12802 56550 12832 56602
rect 12856 56550 12866 56602
rect 12866 56550 12912 56602
rect 12616 56548 12672 56550
rect 12696 56548 12752 56550
rect 12776 56548 12832 56550
rect 12856 56548 12912 56550
rect 12616 55514 12672 55516
rect 12696 55514 12752 55516
rect 12776 55514 12832 55516
rect 12856 55514 12912 55516
rect 12616 55462 12662 55514
rect 12662 55462 12672 55514
rect 12696 55462 12726 55514
rect 12726 55462 12738 55514
rect 12738 55462 12752 55514
rect 12776 55462 12790 55514
rect 12790 55462 12802 55514
rect 12802 55462 12832 55514
rect 12856 55462 12866 55514
rect 12866 55462 12912 55514
rect 12616 55460 12672 55462
rect 12696 55460 12752 55462
rect 12776 55460 12832 55462
rect 12856 55460 12912 55462
rect 11956 54970 12012 54972
rect 12036 54970 12092 54972
rect 12116 54970 12172 54972
rect 12196 54970 12252 54972
rect 11956 54918 12002 54970
rect 12002 54918 12012 54970
rect 12036 54918 12066 54970
rect 12066 54918 12078 54970
rect 12078 54918 12092 54970
rect 12116 54918 12130 54970
rect 12130 54918 12142 54970
rect 12142 54918 12172 54970
rect 12196 54918 12206 54970
rect 12206 54918 12252 54970
rect 11956 54916 12012 54918
rect 12036 54916 12092 54918
rect 12116 54916 12172 54918
rect 12196 54916 12252 54918
rect 12616 54426 12672 54428
rect 12696 54426 12752 54428
rect 12776 54426 12832 54428
rect 12856 54426 12912 54428
rect 12616 54374 12662 54426
rect 12662 54374 12672 54426
rect 12696 54374 12726 54426
rect 12726 54374 12738 54426
rect 12738 54374 12752 54426
rect 12776 54374 12790 54426
rect 12790 54374 12802 54426
rect 12802 54374 12832 54426
rect 12856 54374 12866 54426
rect 12866 54374 12912 54426
rect 12616 54372 12672 54374
rect 12696 54372 12752 54374
rect 12776 54372 12832 54374
rect 12856 54372 12912 54374
rect 11956 53882 12012 53884
rect 12036 53882 12092 53884
rect 12116 53882 12172 53884
rect 12196 53882 12252 53884
rect 11956 53830 12002 53882
rect 12002 53830 12012 53882
rect 12036 53830 12066 53882
rect 12066 53830 12078 53882
rect 12078 53830 12092 53882
rect 12116 53830 12130 53882
rect 12130 53830 12142 53882
rect 12142 53830 12172 53882
rect 12196 53830 12206 53882
rect 12206 53830 12252 53882
rect 11956 53828 12012 53830
rect 12036 53828 12092 53830
rect 12116 53828 12172 53830
rect 12196 53828 12252 53830
rect 12616 53338 12672 53340
rect 12696 53338 12752 53340
rect 12776 53338 12832 53340
rect 12856 53338 12912 53340
rect 12616 53286 12662 53338
rect 12662 53286 12672 53338
rect 12696 53286 12726 53338
rect 12726 53286 12738 53338
rect 12738 53286 12752 53338
rect 12776 53286 12790 53338
rect 12790 53286 12802 53338
rect 12802 53286 12832 53338
rect 12856 53286 12866 53338
rect 12866 53286 12912 53338
rect 12616 53284 12672 53286
rect 12696 53284 12752 53286
rect 12776 53284 12832 53286
rect 12856 53284 12912 53286
rect 11956 52794 12012 52796
rect 12036 52794 12092 52796
rect 12116 52794 12172 52796
rect 12196 52794 12252 52796
rect 11956 52742 12002 52794
rect 12002 52742 12012 52794
rect 12036 52742 12066 52794
rect 12066 52742 12078 52794
rect 12078 52742 12092 52794
rect 12116 52742 12130 52794
rect 12130 52742 12142 52794
rect 12142 52742 12172 52794
rect 12196 52742 12206 52794
rect 12206 52742 12252 52794
rect 11956 52740 12012 52742
rect 12036 52740 12092 52742
rect 12116 52740 12172 52742
rect 12196 52740 12252 52742
rect 12616 52250 12672 52252
rect 12696 52250 12752 52252
rect 12776 52250 12832 52252
rect 12856 52250 12912 52252
rect 12616 52198 12662 52250
rect 12662 52198 12672 52250
rect 12696 52198 12726 52250
rect 12726 52198 12738 52250
rect 12738 52198 12752 52250
rect 12776 52198 12790 52250
rect 12790 52198 12802 52250
rect 12802 52198 12832 52250
rect 12856 52198 12866 52250
rect 12866 52198 12912 52250
rect 12616 52196 12672 52198
rect 12696 52196 12752 52198
rect 12776 52196 12832 52198
rect 12856 52196 12912 52198
rect 11956 51706 12012 51708
rect 12036 51706 12092 51708
rect 12116 51706 12172 51708
rect 12196 51706 12252 51708
rect 11956 51654 12002 51706
rect 12002 51654 12012 51706
rect 12036 51654 12066 51706
rect 12066 51654 12078 51706
rect 12078 51654 12092 51706
rect 12116 51654 12130 51706
rect 12130 51654 12142 51706
rect 12142 51654 12172 51706
rect 12196 51654 12206 51706
rect 12206 51654 12252 51706
rect 11956 51652 12012 51654
rect 12036 51652 12092 51654
rect 12116 51652 12172 51654
rect 12196 51652 12252 51654
rect 11956 50618 12012 50620
rect 12036 50618 12092 50620
rect 12116 50618 12172 50620
rect 12196 50618 12252 50620
rect 11956 50566 12002 50618
rect 12002 50566 12012 50618
rect 12036 50566 12066 50618
rect 12066 50566 12078 50618
rect 12078 50566 12092 50618
rect 12116 50566 12130 50618
rect 12130 50566 12142 50618
rect 12142 50566 12172 50618
rect 12196 50566 12206 50618
rect 12206 50566 12252 50618
rect 11956 50564 12012 50566
rect 12036 50564 12092 50566
rect 12116 50564 12172 50566
rect 12196 50564 12252 50566
rect 11956 49530 12012 49532
rect 12036 49530 12092 49532
rect 12116 49530 12172 49532
rect 12196 49530 12252 49532
rect 11956 49478 12002 49530
rect 12002 49478 12012 49530
rect 12036 49478 12066 49530
rect 12066 49478 12078 49530
rect 12078 49478 12092 49530
rect 12116 49478 12130 49530
rect 12130 49478 12142 49530
rect 12142 49478 12172 49530
rect 12196 49478 12206 49530
rect 12206 49478 12252 49530
rect 11956 49476 12012 49478
rect 12036 49476 12092 49478
rect 12116 49476 12172 49478
rect 12196 49476 12252 49478
rect 11956 48442 12012 48444
rect 12036 48442 12092 48444
rect 12116 48442 12172 48444
rect 12196 48442 12252 48444
rect 11956 48390 12002 48442
rect 12002 48390 12012 48442
rect 12036 48390 12066 48442
rect 12066 48390 12078 48442
rect 12078 48390 12092 48442
rect 12116 48390 12130 48442
rect 12130 48390 12142 48442
rect 12142 48390 12172 48442
rect 12196 48390 12206 48442
rect 12206 48390 12252 48442
rect 11956 48388 12012 48390
rect 12036 48388 12092 48390
rect 12116 48388 12172 48390
rect 12196 48388 12252 48390
rect 11956 47354 12012 47356
rect 12036 47354 12092 47356
rect 12116 47354 12172 47356
rect 12196 47354 12252 47356
rect 11956 47302 12002 47354
rect 12002 47302 12012 47354
rect 12036 47302 12066 47354
rect 12066 47302 12078 47354
rect 12078 47302 12092 47354
rect 12116 47302 12130 47354
rect 12130 47302 12142 47354
rect 12142 47302 12172 47354
rect 12196 47302 12206 47354
rect 12206 47302 12252 47354
rect 11956 47300 12012 47302
rect 12036 47300 12092 47302
rect 12116 47300 12172 47302
rect 12196 47300 12252 47302
rect 11956 46266 12012 46268
rect 12036 46266 12092 46268
rect 12116 46266 12172 46268
rect 12196 46266 12252 46268
rect 11956 46214 12002 46266
rect 12002 46214 12012 46266
rect 12036 46214 12066 46266
rect 12066 46214 12078 46266
rect 12078 46214 12092 46266
rect 12116 46214 12130 46266
rect 12130 46214 12142 46266
rect 12142 46214 12172 46266
rect 12196 46214 12206 46266
rect 12206 46214 12252 46266
rect 11956 46212 12012 46214
rect 12036 46212 12092 46214
rect 12116 46212 12172 46214
rect 12196 46212 12252 46214
rect 11956 45178 12012 45180
rect 12036 45178 12092 45180
rect 12116 45178 12172 45180
rect 12196 45178 12252 45180
rect 11956 45126 12002 45178
rect 12002 45126 12012 45178
rect 12036 45126 12066 45178
rect 12066 45126 12078 45178
rect 12078 45126 12092 45178
rect 12116 45126 12130 45178
rect 12130 45126 12142 45178
rect 12142 45126 12172 45178
rect 12196 45126 12206 45178
rect 12206 45126 12252 45178
rect 11956 45124 12012 45126
rect 12036 45124 12092 45126
rect 12116 45124 12172 45126
rect 12196 45124 12252 45126
rect 11956 44090 12012 44092
rect 12036 44090 12092 44092
rect 12116 44090 12172 44092
rect 12196 44090 12252 44092
rect 11956 44038 12002 44090
rect 12002 44038 12012 44090
rect 12036 44038 12066 44090
rect 12066 44038 12078 44090
rect 12078 44038 12092 44090
rect 12116 44038 12130 44090
rect 12130 44038 12142 44090
rect 12142 44038 12172 44090
rect 12196 44038 12206 44090
rect 12206 44038 12252 44090
rect 11956 44036 12012 44038
rect 12036 44036 12092 44038
rect 12116 44036 12172 44038
rect 12196 44036 12252 44038
rect 11956 43002 12012 43004
rect 12036 43002 12092 43004
rect 12116 43002 12172 43004
rect 12196 43002 12252 43004
rect 11956 42950 12002 43002
rect 12002 42950 12012 43002
rect 12036 42950 12066 43002
rect 12066 42950 12078 43002
rect 12078 42950 12092 43002
rect 12116 42950 12130 43002
rect 12130 42950 12142 43002
rect 12142 42950 12172 43002
rect 12196 42950 12206 43002
rect 12206 42950 12252 43002
rect 11956 42948 12012 42950
rect 12036 42948 12092 42950
rect 12116 42948 12172 42950
rect 12196 42948 12252 42950
rect 11956 41914 12012 41916
rect 12036 41914 12092 41916
rect 12116 41914 12172 41916
rect 12196 41914 12252 41916
rect 11956 41862 12002 41914
rect 12002 41862 12012 41914
rect 12036 41862 12066 41914
rect 12066 41862 12078 41914
rect 12078 41862 12092 41914
rect 12116 41862 12130 41914
rect 12130 41862 12142 41914
rect 12142 41862 12172 41914
rect 12196 41862 12206 41914
rect 12206 41862 12252 41914
rect 11956 41860 12012 41862
rect 12036 41860 12092 41862
rect 12116 41860 12172 41862
rect 12196 41860 12252 41862
rect 11956 40826 12012 40828
rect 12036 40826 12092 40828
rect 12116 40826 12172 40828
rect 12196 40826 12252 40828
rect 11956 40774 12002 40826
rect 12002 40774 12012 40826
rect 12036 40774 12066 40826
rect 12066 40774 12078 40826
rect 12078 40774 12092 40826
rect 12116 40774 12130 40826
rect 12130 40774 12142 40826
rect 12142 40774 12172 40826
rect 12196 40774 12206 40826
rect 12206 40774 12252 40826
rect 11956 40772 12012 40774
rect 12036 40772 12092 40774
rect 12116 40772 12172 40774
rect 12196 40772 12252 40774
rect 11956 39738 12012 39740
rect 12036 39738 12092 39740
rect 12116 39738 12172 39740
rect 12196 39738 12252 39740
rect 11956 39686 12002 39738
rect 12002 39686 12012 39738
rect 12036 39686 12066 39738
rect 12066 39686 12078 39738
rect 12078 39686 12092 39738
rect 12116 39686 12130 39738
rect 12130 39686 12142 39738
rect 12142 39686 12172 39738
rect 12196 39686 12206 39738
rect 12206 39686 12252 39738
rect 11956 39684 12012 39686
rect 12036 39684 12092 39686
rect 12116 39684 12172 39686
rect 12196 39684 12252 39686
rect 11956 38650 12012 38652
rect 12036 38650 12092 38652
rect 12116 38650 12172 38652
rect 12196 38650 12252 38652
rect 11956 38598 12002 38650
rect 12002 38598 12012 38650
rect 12036 38598 12066 38650
rect 12066 38598 12078 38650
rect 12078 38598 12092 38650
rect 12116 38598 12130 38650
rect 12130 38598 12142 38650
rect 12142 38598 12172 38650
rect 12196 38598 12206 38650
rect 12206 38598 12252 38650
rect 11956 38596 12012 38598
rect 12036 38596 12092 38598
rect 12116 38596 12172 38598
rect 12196 38596 12252 38598
rect 11956 37562 12012 37564
rect 12036 37562 12092 37564
rect 12116 37562 12172 37564
rect 12196 37562 12252 37564
rect 11956 37510 12002 37562
rect 12002 37510 12012 37562
rect 12036 37510 12066 37562
rect 12066 37510 12078 37562
rect 12078 37510 12092 37562
rect 12116 37510 12130 37562
rect 12130 37510 12142 37562
rect 12142 37510 12172 37562
rect 12196 37510 12206 37562
rect 12206 37510 12252 37562
rect 11956 37508 12012 37510
rect 12036 37508 12092 37510
rect 12116 37508 12172 37510
rect 12196 37508 12252 37510
rect 11956 36474 12012 36476
rect 12036 36474 12092 36476
rect 12116 36474 12172 36476
rect 12196 36474 12252 36476
rect 11956 36422 12002 36474
rect 12002 36422 12012 36474
rect 12036 36422 12066 36474
rect 12066 36422 12078 36474
rect 12078 36422 12092 36474
rect 12116 36422 12130 36474
rect 12130 36422 12142 36474
rect 12142 36422 12172 36474
rect 12196 36422 12206 36474
rect 12206 36422 12252 36474
rect 11956 36420 12012 36422
rect 12036 36420 12092 36422
rect 12116 36420 12172 36422
rect 12196 36420 12252 36422
rect 11956 35386 12012 35388
rect 12036 35386 12092 35388
rect 12116 35386 12172 35388
rect 12196 35386 12252 35388
rect 11956 35334 12002 35386
rect 12002 35334 12012 35386
rect 12036 35334 12066 35386
rect 12066 35334 12078 35386
rect 12078 35334 12092 35386
rect 12116 35334 12130 35386
rect 12130 35334 12142 35386
rect 12142 35334 12172 35386
rect 12196 35334 12206 35386
rect 12206 35334 12252 35386
rect 11956 35332 12012 35334
rect 12036 35332 12092 35334
rect 12116 35332 12172 35334
rect 12196 35332 12252 35334
rect 11956 34298 12012 34300
rect 12036 34298 12092 34300
rect 12116 34298 12172 34300
rect 12196 34298 12252 34300
rect 11956 34246 12002 34298
rect 12002 34246 12012 34298
rect 12036 34246 12066 34298
rect 12066 34246 12078 34298
rect 12078 34246 12092 34298
rect 12116 34246 12130 34298
rect 12130 34246 12142 34298
rect 12142 34246 12172 34298
rect 12196 34246 12206 34298
rect 12206 34246 12252 34298
rect 11956 34244 12012 34246
rect 12036 34244 12092 34246
rect 12116 34244 12172 34246
rect 12196 34244 12252 34246
rect 11956 33210 12012 33212
rect 12036 33210 12092 33212
rect 12116 33210 12172 33212
rect 12196 33210 12252 33212
rect 11956 33158 12002 33210
rect 12002 33158 12012 33210
rect 12036 33158 12066 33210
rect 12066 33158 12078 33210
rect 12078 33158 12092 33210
rect 12116 33158 12130 33210
rect 12130 33158 12142 33210
rect 12142 33158 12172 33210
rect 12196 33158 12206 33210
rect 12206 33158 12252 33210
rect 11956 33156 12012 33158
rect 12036 33156 12092 33158
rect 12116 33156 12172 33158
rect 12196 33156 12252 33158
rect 11956 32122 12012 32124
rect 12036 32122 12092 32124
rect 12116 32122 12172 32124
rect 12196 32122 12252 32124
rect 11956 32070 12002 32122
rect 12002 32070 12012 32122
rect 12036 32070 12066 32122
rect 12066 32070 12078 32122
rect 12078 32070 12092 32122
rect 12116 32070 12130 32122
rect 12130 32070 12142 32122
rect 12142 32070 12172 32122
rect 12196 32070 12206 32122
rect 12206 32070 12252 32122
rect 11956 32068 12012 32070
rect 12036 32068 12092 32070
rect 12116 32068 12172 32070
rect 12196 32068 12252 32070
rect 12616 51162 12672 51164
rect 12696 51162 12752 51164
rect 12776 51162 12832 51164
rect 12856 51162 12912 51164
rect 12616 51110 12662 51162
rect 12662 51110 12672 51162
rect 12696 51110 12726 51162
rect 12726 51110 12738 51162
rect 12738 51110 12752 51162
rect 12776 51110 12790 51162
rect 12790 51110 12802 51162
rect 12802 51110 12832 51162
rect 12856 51110 12866 51162
rect 12866 51110 12912 51162
rect 12616 51108 12672 51110
rect 12696 51108 12752 51110
rect 12776 51108 12832 51110
rect 12856 51108 12912 51110
rect 12616 50074 12672 50076
rect 12696 50074 12752 50076
rect 12776 50074 12832 50076
rect 12856 50074 12912 50076
rect 12616 50022 12662 50074
rect 12662 50022 12672 50074
rect 12696 50022 12726 50074
rect 12726 50022 12738 50074
rect 12738 50022 12752 50074
rect 12776 50022 12790 50074
rect 12790 50022 12802 50074
rect 12802 50022 12832 50074
rect 12856 50022 12866 50074
rect 12866 50022 12912 50074
rect 12616 50020 12672 50022
rect 12696 50020 12752 50022
rect 12776 50020 12832 50022
rect 12856 50020 12912 50022
rect 12616 48986 12672 48988
rect 12696 48986 12752 48988
rect 12776 48986 12832 48988
rect 12856 48986 12912 48988
rect 12616 48934 12662 48986
rect 12662 48934 12672 48986
rect 12696 48934 12726 48986
rect 12726 48934 12738 48986
rect 12738 48934 12752 48986
rect 12776 48934 12790 48986
rect 12790 48934 12802 48986
rect 12802 48934 12832 48986
rect 12856 48934 12866 48986
rect 12866 48934 12912 48986
rect 12616 48932 12672 48934
rect 12696 48932 12752 48934
rect 12776 48932 12832 48934
rect 12856 48932 12912 48934
rect 12616 47898 12672 47900
rect 12696 47898 12752 47900
rect 12776 47898 12832 47900
rect 12856 47898 12912 47900
rect 12616 47846 12662 47898
rect 12662 47846 12672 47898
rect 12696 47846 12726 47898
rect 12726 47846 12738 47898
rect 12738 47846 12752 47898
rect 12776 47846 12790 47898
rect 12790 47846 12802 47898
rect 12802 47846 12832 47898
rect 12856 47846 12866 47898
rect 12866 47846 12912 47898
rect 12616 47844 12672 47846
rect 12696 47844 12752 47846
rect 12776 47844 12832 47846
rect 12856 47844 12912 47846
rect 12616 46810 12672 46812
rect 12696 46810 12752 46812
rect 12776 46810 12832 46812
rect 12856 46810 12912 46812
rect 12616 46758 12662 46810
rect 12662 46758 12672 46810
rect 12696 46758 12726 46810
rect 12726 46758 12738 46810
rect 12738 46758 12752 46810
rect 12776 46758 12790 46810
rect 12790 46758 12802 46810
rect 12802 46758 12832 46810
rect 12856 46758 12866 46810
rect 12866 46758 12912 46810
rect 12616 46756 12672 46758
rect 12696 46756 12752 46758
rect 12776 46756 12832 46758
rect 12856 46756 12912 46758
rect 12616 45722 12672 45724
rect 12696 45722 12752 45724
rect 12776 45722 12832 45724
rect 12856 45722 12912 45724
rect 12616 45670 12662 45722
rect 12662 45670 12672 45722
rect 12696 45670 12726 45722
rect 12726 45670 12738 45722
rect 12738 45670 12752 45722
rect 12776 45670 12790 45722
rect 12790 45670 12802 45722
rect 12802 45670 12832 45722
rect 12856 45670 12866 45722
rect 12866 45670 12912 45722
rect 12616 45668 12672 45670
rect 12696 45668 12752 45670
rect 12776 45668 12832 45670
rect 12856 45668 12912 45670
rect 12616 44634 12672 44636
rect 12696 44634 12752 44636
rect 12776 44634 12832 44636
rect 12856 44634 12912 44636
rect 12616 44582 12662 44634
rect 12662 44582 12672 44634
rect 12696 44582 12726 44634
rect 12726 44582 12738 44634
rect 12738 44582 12752 44634
rect 12776 44582 12790 44634
rect 12790 44582 12802 44634
rect 12802 44582 12832 44634
rect 12856 44582 12866 44634
rect 12866 44582 12912 44634
rect 12616 44580 12672 44582
rect 12696 44580 12752 44582
rect 12776 44580 12832 44582
rect 12856 44580 12912 44582
rect 12616 43546 12672 43548
rect 12696 43546 12752 43548
rect 12776 43546 12832 43548
rect 12856 43546 12912 43548
rect 12616 43494 12662 43546
rect 12662 43494 12672 43546
rect 12696 43494 12726 43546
rect 12726 43494 12738 43546
rect 12738 43494 12752 43546
rect 12776 43494 12790 43546
rect 12790 43494 12802 43546
rect 12802 43494 12832 43546
rect 12856 43494 12866 43546
rect 12866 43494 12912 43546
rect 12616 43492 12672 43494
rect 12696 43492 12752 43494
rect 12776 43492 12832 43494
rect 12856 43492 12912 43494
rect 12616 42458 12672 42460
rect 12696 42458 12752 42460
rect 12776 42458 12832 42460
rect 12856 42458 12912 42460
rect 12616 42406 12662 42458
rect 12662 42406 12672 42458
rect 12696 42406 12726 42458
rect 12726 42406 12738 42458
rect 12738 42406 12752 42458
rect 12776 42406 12790 42458
rect 12790 42406 12802 42458
rect 12802 42406 12832 42458
rect 12856 42406 12866 42458
rect 12866 42406 12912 42458
rect 12616 42404 12672 42406
rect 12696 42404 12752 42406
rect 12776 42404 12832 42406
rect 12856 42404 12912 42406
rect 12616 41370 12672 41372
rect 12696 41370 12752 41372
rect 12776 41370 12832 41372
rect 12856 41370 12912 41372
rect 12616 41318 12662 41370
rect 12662 41318 12672 41370
rect 12696 41318 12726 41370
rect 12726 41318 12738 41370
rect 12738 41318 12752 41370
rect 12776 41318 12790 41370
rect 12790 41318 12802 41370
rect 12802 41318 12832 41370
rect 12856 41318 12866 41370
rect 12866 41318 12912 41370
rect 12616 41316 12672 41318
rect 12696 41316 12752 41318
rect 12776 41316 12832 41318
rect 12856 41316 12912 41318
rect 12616 40282 12672 40284
rect 12696 40282 12752 40284
rect 12776 40282 12832 40284
rect 12856 40282 12912 40284
rect 12616 40230 12662 40282
rect 12662 40230 12672 40282
rect 12696 40230 12726 40282
rect 12726 40230 12738 40282
rect 12738 40230 12752 40282
rect 12776 40230 12790 40282
rect 12790 40230 12802 40282
rect 12802 40230 12832 40282
rect 12856 40230 12866 40282
rect 12866 40230 12912 40282
rect 12616 40228 12672 40230
rect 12696 40228 12752 40230
rect 12776 40228 12832 40230
rect 12856 40228 12912 40230
rect 12616 39194 12672 39196
rect 12696 39194 12752 39196
rect 12776 39194 12832 39196
rect 12856 39194 12912 39196
rect 12616 39142 12662 39194
rect 12662 39142 12672 39194
rect 12696 39142 12726 39194
rect 12726 39142 12738 39194
rect 12738 39142 12752 39194
rect 12776 39142 12790 39194
rect 12790 39142 12802 39194
rect 12802 39142 12832 39194
rect 12856 39142 12866 39194
rect 12866 39142 12912 39194
rect 12616 39140 12672 39142
rect 12696 39140 12752 39142
rect 12776 39140 12832 39142
rect 12856 39140 12912 39142
rect 12616 38106 12672 38108
rect 12696 38106 12752 38108
rect 12776 38106 12832 38108
rect 12856 38106 12912 38108
rect 12616 38054 12662 38106
rect 12662 38054 12672 38106
rect 12696 38054 12726 38106
rect 12726 38054 12738 38106
rect 12738 38054 12752 38106
rect 12776 38054 12790 38106
rect 12790 38054 12802 38106
rect 12802 38054 12832 38106
rect 12856 38054 12866 38106
rect 12866 38054 12912 38106
rect 12616 38052 12672 38054
rect 12696 38052 12752 38054
rect 12776 38052 12832 38054
rect 12856 38052 12912 38054
rect 12616 37018 12672 37020
rect 12696 37018 12752 37020
rect 12776 37018 12832 37020
rect 12856 37018 12912 37020
rect 12616 36966 12662 37018
rect 12662 36966 12672 37018
rect 12696 36966 12726 37018
rect 12726 36966 12738 37018
rect 12738 36966 12752 37018
rect 12776 36966 12790 37018
rect 12790 36966 12802 37018
rect 12802 36966 12832 37018
rect 12856 36966 12866 37018
rect 12866 36966 12912 37018
rect 12616 36964 12672 36966
rect 12696 36964 12752 36966
rect 12776 36964 12832 36966
rect 12856 36964 12912 36966
rect 12616 35930 12672 35932
rect 12696 35930 12752 35932
rect 12776 35930 12832 35932
rect 12856 35930 12912 35932
rect 12616 35878 12662 35930
rect 12662 35878 12672 35930
rect 12696 35878 12726 35930
rect 12726 35878 12738 35930
rect 12738 35878 12752 35930
rect 12776 35878 12790 35930
rect 12790 35878 12802 35930
rect 12802 35878 12832 35930
rect 12856 35878 12866 35930
rect 12866 35878 12912 35930
rect 12616 35876 12672 35878
rect 12696 35876 12752 35878
rect 12776 35876 12832 35878
rect 12856 35876 12912 35878
rect 12616 34842 12672 34844
rect 12696 34842 12752 34844
rect 12776 34842 12832 34844
rect 12856 34842 12912 34844
rect 12616 34790 12662 34842
rect 12662 34790 12672 34842
rect 12696 34790 12726 34842
rect 12726 34790 12738 34842
rect 12738 34790 12752 34842
rect 12776 34790 12790 34842
rect 12790 34790 12802 34842
rect 12802 34790 12832 34842
rect 12856 34790 12866 34842
rect 12866 34790 12912 34842
rect 12616 34788 12672 34790
rect 12696 34788 12752 34790
rect 12776 34788 12832 34790
rect 12856 34788 12912 34790
rect 12616 33754 12672 33756
rect 12696 33754 12752 33756
rect 12776 33754 12832 33756
rect 12856 33754 12912 33756
rect 12616 33702 12662 33754
rect 12662 33702 12672 33754
rect 12696 33702 12726 33754
rect 12726 33702 12738 33754
rect 12738 33702 12752 33754
rect 12776 33702 12790 33754
rect 12790 33702 12802 33754
rect 12802 33702 12832 33754
rect 12856 33702 12866 33754
rect 12866 33702 12912 33754
rect 12616 33700 12672 33702
rect 12696 33700 12752 33702
rect 12776 33700 12832 33702
rect 12856 33700 12912 33702
rect 12616 32666 12672 32668
rect 12696 32666 12752 32668
rect 12776 32666 12832 32668
rect 12856 32666 12912 32668
rect 12616 32614 12662 32666
rect 12662 32614 12672 32666
rect 12696 32614 12726 32666
rect 12726 32614 12738 32666
rect 12738 32614 12752 32666
rect 12776 32614 12790 32666
rect 12790 32614 12802 32666
rect 12802 32614 12832 32666
rect 12856 32614 12866 32666
rect 12866 32614 12912 32666
rect 12616 32612 12672 32614
rect 12696 32612 12752 32614
rect 12776 32612 12832 32614
rect 12856 32612 12912 32614
rect 11956 31034 12012 31036
rect 12036 31034 12092 31036
rect 12116 31034 12172 31036
rect 12196 31034 12252 31036
rect 11956 30982 12002 31034
rect 12002 30982 12012 31034
rect 12036 30982 12066 31034
rect 12066 30982 12078 31034
rect 12078 30982 12092 31034
rect 12116 30982 12130 31034
rect 12130 30982 12142 31034
rect 12142 30982 12172 31034
rect 12196 30982 12206 31034
rect 12206 30982 12252 31034
rect 11956 30980 12012 30982
rect 12036 30980 12092 30982
rect 12116 30980 12172 30982
rect 12196 30980 12252 30982
rect 11956 29946 12012 29948
rect 12036 29946 12092 29948
rect 12116 29946 12172 29948
rect 12196 29946 12252 29948
rect 11956 29894 12002 29946
rect 12002 29894 12012 29946
rect 12036 29894 12066 29946
rect 12066 29894 12078 29946
rect 12078 29894 12092 29946
rect 12116 29894 12130 29946
rect 12130 29894 12142 29946
rect 12142 29894 12172 29946
rect 12196 29894 12206 29946
rect 12206 29894 12252 29946
rect 11956 29892 12012 29894
rect 12036 29892 12092 29894
rect 12116 29892 12172 29894
rect 12196 29892 12252 29894
rect 11956 28858 12012 28860
rect 12036 28858 12092 28860
rect 12116 28858 12172 28860
rect 12196 28858 12252 28860
rect 11956 28806 12002 28858
rect 12002 28806 12012 28858
rect 12036 28806 12066 28858
rect 12066 28806 12078 28858
rect 12078 28806 12092 28858
rect 12116 28806 12130 28858
rect 12130 28806 12142 28858
rect 12142 28806 12172 28858
rect 12196 28806 12206 28858
rect 12206 28806 12252 28858
rect 11956 28804 12012 28806
rect 12036 28804 12092 28806
rect 12116 28804 12172 28806
rect 12196 28804 12252 28806
rect 11956 27770 12012 27772
rect 12036 27770 12092 27772
rect 12116 27770 12172 27772
rect 12196 27770 12252 27772
rect 11956 27718 12002 27770
rect 12002 27718 12012 27770
rect 12036 27718 12066 27770
rect 12066 27718 12078 27770
rect 12078 27718 12092 27770
rect 12116 27718 12130 27770
rect 12130 27718 12142 27770
rect 12142 27718 12172 27770
rect 12196 27718 12206 27770
rect 12206 27718 12252 27770
rect 11956 27716 12012 27718
rect 12036 27716 12092 27718
rect 12116 27716 12172 27718
rect 12196 27716 12252 27718
rect 12616 31578 12672 31580
rect 12696 31578 12752 31580
rect 12776 31578 12832 31580
rect 12856 31578 12912 31580
rect 12616 31526 12662 31578
rect 12662 31526 12672 31578
rect 12696 31526 12726 31578
rect 12726 31526 12738 31578
rect 12738 31526 12752 31578
rect 12776 31526 12790 31578
rect 12790 31526 12802 31578
rect 12802 31526 12832 31578
rect 12856 31526 12866 31578
rect 12866 31526 12912 31578
rect 12616 31524 12672 31526
rect 12696 31524 12752 31526
rect 12776 31524 12832 31526
rect 12856 31524 12912 31526
rect 12616 30490 12672 30492
rect 12696 30490 12752 30492
rect 12776 30490 12832 30492
rect 12856 30490 12912 30492
rect 12616 30438 12662 30490
rect 12662 30438 12672 30490
rect 12696 30438 12726 30490
rect 12726 30438 12738 30490
rect 12738 30438 12752 30490
rect 12776 30438 12790 30490
rect 12790 30438 12802 30490
rect 12802 30438 12832 30490
rect 12856 30438 12866 30490
rect 12866 30438 12912 30490
rect 12616 30436 12672 30438
rect 12696 30436 12752 30438
rect 12776 30436 12832 30438
rect 12856 30436 12912 30438
rect 12616 29402 12672 29404
rect 12696 29402 12752 29404
rect 12776 29402 12832 29404
rect 12856 29402 12912 29404
rect 12616 29350 12662 29402
rect 12662 29350 12672 29402
rect 12696 29350 12726 29402
rect 12726 29350 12738 29402
rect 12738 29350 12752 29402
rect 12776 29350 12790 29402
rect 12790 29350 12802 29402
rect 12802 29350 12832 29402
rect 12856 29350 12866 29402
rect 12866 29350 12912 29402
rect 12616 29348 12672 29350
rect 12696 29348 12752 29350
rect 12776 29348 12832 29350
rect 12856 29348 12912 29350
rect 12616 28314 12672 28316
rect 12696 28314 12752 28316
rect 12776 28314 12832 28316
rect 12856 28314 12912 28316
rect 12616 28262 12662 28314
rect 12662 28262 12672 28314
rect 12696 28262 12726 28314
rect 12726 28262 12738 28314
rect 12738 28262 12752 28314
rect 12776 28262 12790 28314
rect 12790 28262 12802 28314
rect 12802 28262 12832 28314
rect 12856 28262 12866 28314
rect 12866 28262 12912 28314
rect 12616 28260 12672 28262
rect 12696 28260 12752 28262
rect 12776 28260 12832 28262
rect 12856 28260 12912 28262
rect 11956 26682 12012 26684
rect 12036 26682 12092 26684
rect 12116 26682 12172 26684
rect 12196 26682 12252 26684
rect 11956 26630 12002 26682
rect 12002 26630 12012 26682
rect 12036 26630 12066 26682
rect 12066 26630 12078 26682
rect 12078 26630 12092 26682
rect 12116 26630 12130 26682
rect 12130 26630 12142 26682
rect 12142 26630 12172 26682
rect 12196 26630 12206 26682
rect 12206 26630 12252 26682
rect 11956 26628 12012 26630
rect 12036 26628 12092 26630
rect 12116 26628 12172 26630
rect 12196 26628 12252 26630
rect 11956 25594 12012 25596
rect 12036 25594 12092 25596
rect 12116 25594 12172 25596
rect 12196 25594 12252 25596
rect 11956 25542 12002 25594
rect 12002 25542 12012 25594
rect 12036 25542 12066 25594
rect 12066 25542 12078 25594
rect 12078 25542 12092 25594
rect 12116 25542 12130 25594
rect 12130 25542 12142 25594
rect 12142 25542 12172 25594
rect 12196 25542 12206 25594
rect 12206 25542 12252 25594
rect 11956 25540 12012 25542
rect 12036 25540 12092 25542
rect 12116 25540 12172 25542
rect 12196 25540 12252 25542
rect 11956 24506 12012 24508
rect 12036 24506 12092 24508
rect 12116 24506 12172 24508
rect 12196 24506 12252 24508
rect 11956 24454 12002 24506
rect 12002 24454 12012 24506
rect 12036 24454 12066 24506
rect 12066 24454 12078 24506
rect 12078 24454 12092 24506
rect 12116 24454 12130 24506
rect 12130 24454 12142 24506
rect 12142 24454 12172 24506
rect 12196 24454 12206 24506
rect 12206 24454 12252 24506
rect 11956 24452 12012 24454
rect 12036 24452 12092 24454
rect 12116 24452 12172 24454
rect 12196 24452 12252 24454
rect 11956 23418 12012 23420
rect 12036 23418 12092 23420
rect 12116 23418 12172 23420
rect 12196 23418 12252 23420
rect 11956 23366 12002 23418
rect 12002 23366 12012 23418
rect 12036 23366 12066 23418
rect 12066 23366 12078 23418
rect 12078 23366 12092 23418
rect 12116 23366 12130 23418
rect 12130 23366 12142 23418
rect 12142 23366 12172 23418
rect 12196 23366 12206 23418
rect 12206 23366 12252 23418
rect 11956 23364 12012 23366
rect 12036 23364 12092 23366
rect 12116 23364 12172 23366
rect 12196 23364 12252 23366
rect 11956 22330 12012 22332
rect 12036 22330 12092 22332
rect 12116 22330 12172 22332
rect 12196 22330 12252 22332
rect 11956 22278 12002 22330
rect 12002 22278 12012 22330
rect 12036 22278 12066 22330
rect 12066 22278 12078 22330
rect 12078 22278 12092 22330
rect 12116 22278 12130 22330
rect 12130 22278 12142 22330
rect 12142 22278 12172 22330
rect 12196 22278 12206 22330
rect 12206 22278 12252 22330
rect 11956 22276 12012 22278
rect 12036 22276 12092 22278
rect 12116 22276 12172 22278
rect 12196 22276 12252 22278
rect 11058 21956 11114 21992
rect 11058 21936 11060 21956
rect 11060 21936 11112 21956
rect 11112 21936 11114 21956
rect 11956 21242 12012 21244
rect 12036 21242 12092 21244
rect 12116 21242 12172 21244
rect 12196 21242 12252 21244
rect 11956 21190 12002 21242
rect 12002 21190 12012 21242
rect 12036 21190 12066 21242
rect 12066 21190 12078 21242
rect 12078 21190 12092 21242
rect 12116 21190 12130 21242
rect 12130 21190 12142 21242
rect 12142 21190 12172 21242
rect 12196 21190 12206 21242
rect 12206 21190 12252 21242
rect 11956 21188 12012 21190
rect 12036 21188 12092 21190
rect 12116 21188 12172 21190
rect 12196 21188 12252 21190
rect 11956 20154 12012 20156
rect 12036 20154 12092 20156
rect 12116 20154 12172 20156
rect 12196 20154 12252 20156
rect 11956 20102 12002 20154
rect 12002 20102 12012 20154
rect 12036 20102 12066 20154
rect 12066 20102 12078 20154
rect 12078 20102 12092 20154
rect 12116 20102 12130 20154
rect 12130 20102 12142 20154
rect 12142 20102 12172 20154
rect 12196 20102 12206 20154
rect 12206 20102 12252 20154
rect 11956 20100 12012 20102
rect 12036 20100 12092 20102
rect 12116 20100 12172 20102
rect 12196 20100 12252 20102
rect 11956 19066 12012 19068
rect 12036 19066 12092 19068
rect 12116 19066 12172 19068
rect 12196 19066 12252 19068
rect 11956 19014 12002 19066
rect 12002 19014 12012 19066
rect 12036 19014 12066 19066
rect 12066 19014 12078 19066
rect 12078 19014 12092 19066
rect 12116 19014 12130 19066
rect 12130 19014 12142 19066
rect 12142 19014 12172 19066
rect 12196 19014 12206 19066
rect 12206 19014 12252 19066
rect 11956 19012 12012 19014
rect 12036 19012 12092 19014
rect 12116 19012 12172 19014
rect 12196 19012 12252 19014
rect 11956 17978 12012 17980
rect 12036 17978 12092 17980
rect 12116 17978 12172 17980
rect 12196 17978 12252 17980
rect 11956 17926 12002 17978
rect 12002 17926 12012 17978
rect 12036 17926 12066 17978
rect 12066 17926 12078 17978
rect 12078 17926 12092 17978
rect 12116 17926 12130 17978
rect 12130 17926 12142 17978
rect 12142 17926 12172 17978
rect 12196 17926 12206 17978
rect 12206 17926 12252 17978
rect 11956 17924 12012 17926
rect 12036 17924 12092 17926
rect 12116 17924 12172 17926
rect 12196 17924 12252 17926
rect 11956 16890 12012 16892
rect 12036 16890 12092 16892
rect 12116 16890 12172 16892
rect 12196 16890 12252 16892
rect 11956 16838 12002 16890
rect 12002 16838 12012 16890
rect 12036 16838 12066 16890
rect 12066 16838 12078 16890
rect 12078 16838 12092 16890
rect 12116 16838 12130 16890
rect 12130 16838 12142 16890
rect 12142 16838 12172 16890
rect 12196 16838 12206 16890
rect 12206 16838 12252 16890
rect 11956 16836 12012 16838
rect 12036 16836 12092 16838
rect 12116 16836 12172 16838
rect 12196 16836 12252 16838
rect 11956 15802 12012 15804
rect 12036 15802 12092 15804
rect 12116 15802 12172 15804
rect 12196 15802 12252 15804
rect 11956 15750 12002 15802
rect 12002 15750 12012 15802
rect 12036 15750 12066 15802
rect 12066 15750 12078 15802
rect 12078 15750 12092 15802
rect 12116 15750 12130 15802
rect 12130 15750 12142 15802
rect 12142 15750 12172 15802
rect 12196 15750 12206 15802
rect 12206 15750 12252 15802
rect 11956 15748 12012 15750
rect 12036 15748 12092 15750
rect 12116 15748 12172 15750
rect 12196 15748 12252 15750
rect 11956 14714 12012 14716
rect 12036 14714 12092 14716
rect 12116 14714 12172 14716
rect 12196 14714 12252 14716
rect 11956 14662 12002 14714
rect 12002 14662 12012 14714
rect 12036 14662 12066 14714
rect 12066 14662 12078 14714
rect 12078 14662 12092 14714
rect 12116 14662 12130 14714
rect 12130 14662 12142 14714
rect 12142 14662 12172 14714
rect 12196 14662 12206 14714
rect 12206 14662 12252 14714
rect 11956 14660 12012 14662
rect 12036 14660 12092 14662
rect 12116 14660 12172 14662
rect 12196 14660 12252 14662
rect 11956 13626 12012 13628
rect 12036 13626 12092 13628
rect 12116 13626 12172 13628
rect 12196 13626 12252 13628
rect 11956 13574 12002 13626
rect 12002 13574 12012 13626
rect 12036 13574 12066 13626
rect 12066 13574 12078 13626
rect 12078 13574 12092 13626
rect 12116 13574 12130 13626
rect 12130 13574 12142 13626
rect 12142 13574 12172 13626
rect 12196 13574 12206 13626
rect 12206 13574 12252 13626
rect 11956 13572 12012 13574
rect 12036 13572 12092 13574
rect 12116 13572 12172 13574
rect 12196 13572 12252 13574
rect 11956 12538 12012 12540
rect 12036 12538 12092 12540
rect 12116 12538 12172 12540
rect 12196 12538 12252 12540
rect 11956 12486 12002 12538
rect 12002 12486 12012 12538
rect 12036 12486 12066 12538
rect 12066 12486 12078 12538
rect 12078 12486 12092 12538
rect 12116 12486 12130 12538
rect 12130 12486 12142 12538
rect 12142 12486 12172 12538
rect 12196 12486 12206 12538
rect 12206 12486 12252 12538
rect 11956 12484 12012 12486
rect 12036 12484 12092 12486
rect 12116 12484 12172 12486
rect 12196 12484 12252 12486
rect 11956 11450 12012 11452
rect 12036 11450 12092 11452
rect 12116 11450 12172 11452
rect 12196 11450 12252 11452
rect 11956 11398 12002 11450
rect 12002 11398 12012 11450
rect 12036 11398 12066 11450
rect 12066 11398 12078 11450
rect 12078 11398 12092 11450
rect 12116 11398 12130 11450
rect 12130 11398 12142 11450
rect 12142 11398 12172 11450
rect 12196 11398 12206 11450
rect 12206 11398 12252 11450
rect 11956 11396 12012 11398
rect 12036 11396 12092 11398
rect 12116 11396 12172 11398
rect 12196 11396 12252 11398
rect 11956 10362 12012 10364
rect 12036 10362 12092 10364
rect 12116 10362 12172 10364
rect 12196 10362 12252 10364
rect 11956 10310 12002 10362
rect 12002 10310 12012 10362
rect 12036 10310 12066 10362
rect 12066 10310 12078 10362
rect 12078 10310 12092 10362
rect 12116 10310 12130 10362
rect 12130 10310 12142 10362
rect 12142 10310 12172 10362
rect 12196 10310 12206 10362
rect 12206 10310 12252 10362
rect 11956 10308 12012 10310
rect 12036 10308 12092 10310
rect 12116 10308 12172 10310
rect 12196 10308 12252 10310
rect 11956 9274 12012 9276
rect 12036 9274 12092 9276
rect 12116 9274 12172 9276
rect 12196 9274 12252 9276
rect 11956 9222 12002 9274
rect 12002 9222 12012 9274
rect 12036 9222 12066 9274
rect 12066 9222 12078 9274
rect 12078 9222 12092 9274
rect 12116 9222 12130 9274
rect 12130 9222 12142 9274
rect 12142 9222 12172 9274
rect 12196 9222 12206 9274
rect 12206 9222 12252 9274
rect 11956 9220 12012 9222
rect 12036 9220 12092 9222
rect 12116 9220 12172 9222
rect 12196 9220 12252 9222
rect 11956 8186 12012 8188
rect 12036 8186 12092 8188
rect 12116 8186 12172 8188
rect 12196 8186 12252 8188
rect 11956 8134 12002 8186
rect 12002 8134 12012 8186
rect 12036 8134 12066 8186
rect 12066 8134 12078 8186
rect 12078 8134 12092 8186
rect 12116 8134 12130 8186
rect 12130 8134 12142 8186
rect 12142 8134 12172 8186
rect 12196 8134 12206 8186
rect 12206 8134 12252 8186
rect 11956 8132 12012 8134
rect 12036 8132 12092 8134
rect 12116 8132 12172 8134
rect 12196 8132 12252 8134
rect 11956 7098 12012 7100
rect 12036 7098 12092 7100
rect 12116 7098 12172 7100
rect 12196 7098 12252 7100
rect 11956 7046 12002 7098
rect 12002 7046 12012 7098
rect 12036 7046 12066 7098
rect 12066 7046 12078 7098
rect 12078 7046 12092 7098
rect 12116 7046 12130 7098
rect 12130 7046 12142 7098
rect 12142 7046 12172 7098
rect 12196 7046 12206 7098
rect 12206 7046 12252 7098
rect 11956 7044 12012 7046
rect 12036 7044 12092 7046
rect 12116 7044 12172 7046
rect 12196 7044 12252 7046
rect 11956 6010 12012 6012
rect 12036 6010 12092 6012
rect 12116 6010 12172 6012
rect 12196 6010 12252 6012
rect 11956 5958 12002 6010
rect 12002 5958 12012 6010
rect 12036 5958 12066 6010
rect 12066 5958 12078 6010
rect 12078 5958 12092 6010
rect 12116 5958 12130 6010
rect 12130 5958 12142 6010
rect 12142 5958 12172 6010
rect 12196 5958 12206 6010
rect 12206 5958 12252 6010
rect 11956 5956 12012 5958
rect 12036 5956 12092 5958
rect 12116 5956 12172 5958
rect 12196 5956 12252 5958
rect 11956 4922 12012 4924
rect 12036 4922 12092 4924
rect 12116 4922 12172 4924
rect 12196 4922 12252 4924
rect 11956 4870 12002 4922
rect 12002 4870 12012 4922
rect 12036 4870 12066 4922
rect 12066 4870 12078 4922
rect 12078 4870 12092 4922
rect 12116 4870 12130 4922
rect 12130 4870 12142 4922
rect 12142 4870 12172 4922
rect 12196 4870 12206 4922
rect 12206 4870 12252 4922
rect 11956 4868 12012 4870
rect 12036 4868 12092 4870
rect 12116 4868 12172 4870
rect 12196 4868 12252 4870
rect 12616 27226 12672 27228
rect 12696 27226 12752 27228
rect 12776 27226 12832 27228
rect 12856 27226 12912 27228
rect 12616 27174 12662 27226
rect 12662 27174 12672 27226
rect 12696 27174 12726 27226
rect 12726 27174 12738 27226
rect 12738 27174 12752 27226
rect 12776 27174 12790 27226
rect 12790 27174 12802 27226
rect 12802 27174 12832 27226
rect 12856 27174 12866 27226
rect 12866 27174 12912 27226
rect 12616 27172 12672 27174
rect 12696 27172 12752 27174
rect 12776 27172 12832 27174
rect 12856 27172 12912 27174
rect 12616 26138 12672 26140
rect 12696 26138 12752 26140
rect 12776 26138 12832 26140
rect 12856 26138 12912 26140
rect 12616 26086 12662 26138
rect 12662 26086 12672 26138
rect 12696 26086 12726 26138
rect 12726 26086 12738 26138
rect 12738 26086 12752 26138
rect 12776 26086 12790 26138
rect 12790 26086 12802 26138
rect 12802 26086 12832 26138
rect 12856 26086 12866 26138
rect 12866 26086 12912 26138
rect 12616 26084 12672 26086
rect 12696 26084 12752 26086
rect 12776 26084 12832 26086
rect 12856 26084 12912 26086
rect 12616 25050 12672 25052
rect 12696 25050 12752 25052
rect 12776 25050 12832 25052
rect 12856 25050 12912 25052
rect 12616 24998 12662 25050
rect 12662 24998 12672 25050
rect 12696 24998 12726 25050
rect 12726 24998 12738 25050
rect 12738 24998 12752 25050
rect 12776 24998 12790 25050
rect 12790 24998 12802 25050
rect 12802 24998 12832 25050
rect 12856 24998 12866 25050
rect 12866 24998 12912 25050
rect 12616 24996 12672 24998
rect 12696 24996 12752 24998
rect 12776 24996 12832 24998
rect 12856 24996 12912 24998
rect 12616 23962 12672 23964
rect 12696 23962 12752 23964
rect 12776 23962 12832 23964
rect 12856 23962 12912 23964
rect 12616 23910 12662 23962
rect 12662 23910 12672 23962
rect 12696 23910 12726 23962
rect 12726 23910 12738 23962
rect 12738 23910 12752 23962
rect 12776 23910 12790 23962
rect 12790 23910 12802 23962
rect 12802 23910 12832 23962
rect 12856 23910 12866 23962
rect 12866 23910 12912 23962
rect 12616 23908 12672 23910
rect 12696 23908 12752 23910
rect 12776 23908 12832 23910
rect 12856 23908 12912 23910
rect 12616 22874 12672 22876
rect 12696 22874 12752 22876
rect 12776 22874 12832 22876
rect 12856 22874 12912 22876
rect 12616 22822 12662 22874
rect 12662 22822 12672 22874
rect 12696 22822 12726 22874
rect 12726 22822 12738 22874
rect 12738 22822 12752 22874
rect 12776 22822 12790 22874
rect 12790 22822 12802 22874
rect 12802 22822 12832 22874
rect 12856 22822 12866 22874
rect 12866 22822 12912 22874
rect 12616 22820 12672 22822
rect 12696 22820 12752 22822
rect 12776 22820 12832 22822
rect 12856 22820 12912 22822
rect 12616 21786 12672 21788
rect 12696 21786 12752 21788
rect 12776 21786 12832 21788
rect 12856 21786 12912 21788
rect 12616 21734 12662 21786
rect 12662 21734 12672 21786
rect 12696 21734 12726 21786
rect 12726 21734 12738 21786
rect 12738 21734 12752 21786
rect 12776 21734 12790 21786
rect 12790 21734 12802 21786
rect 12802 21734 12832 21786
rect 12856 21734 12866 21786
rect 12866 21734 12912 21786
rect 12616 21732 12672 21734
rect 12696 21732 12752 21734
rect 12776 21732 12832 21734
rect 12856 21732 12912 21734
rect 12616 20698 12672 20700
rect 12696 20698 12752 20700
rect 12776 20698 12832 20700
rect 12856 20698 12912 20700
rect 12616 20646 12662 20698
rect 12662 20646 12672 20698
rect 12696 20646 12726 20698
rect 12726 20646 12738 20698
rect 12738 20646 12752 20698
rect 12776 20646 12790 20698
rect 12790 20646 12802 20698
rect 12802 20646 12832 20698
rect 12856 20646 12866 20698
rect 12866 20646 12912 20698
rect 12616 20644 12672 20646
rect 12696 20644 12752 20646
rect 12776 20644 12832 20646
rect 12856 20644 12912 20646
rect 12616 19610 12672 19612
rect 12696 19610 12752 19612
rect 12776 19610 12832 19612
rect 12856 19610 12912 19612
rect 12616 19558 12662 19610
rect 12662 19558 12672 19610
rect 12696 19558 12726 19610
rect 12726 19558 12738 19610
rect 12738 19558 12752 19610
rect 12776 19558 12790 19610
rect 12790 19558 12802 19610
rect 12802 19558 12832 19610
rect 12856 19558 12866 19610
rect 12866 19558 12912 19610
rect 12616 19556 12672 19558
rect 12696 19556 12752 19558
rect 12776 19556 12832 19558
rect 12856 19556 12912 19558
rect 12616 18522 12672 18524
rect 12696 18522 12752 18524
rect 12776 18522 12832 18524
rect 12856 18522 12912 18524
rect 12616 18470 12662 18522
rect 12662 18470 12672 18522
rect 12696 18470 12726 18522
rect 12726 18470 12738 18522
rect 12738 18470 12752 18522
rect 12776 18470 12790 18522
rect 12790 18470 12802 18522
rect 12802 18470 12832 18522
rect 12856 18470 12866 18522
rect 12866 18470 12912 18522
rect 12616 18468 12672 18470
rect 12696 18468 12752 18470
rect 12776 18468 12832 18470
rect 12856 18468 12912 18470
rect 12616 17434 12672 17436
rect 12696 17434 12752 17436
rect 12776 17434 12832 17436
rect 12856 17434 12912 17436
rect 12616 17382 12662 17434
rect 12662 17382 12672 17434
rect 12696 17382 12726 17434
rect 12726 17382 12738 17434
rect 12738 17382 12752 17434
rect 12776 17382 12790 17434
rect 12790 17382 12802 17434
rect 12802 17382 12832 17434
rect 12856 17382 12866 17434
rect 12866 17382 12912 17434
rect 12616 17380 12672 17382
rect 12696 17380 12752 17382
rect 12776 17380 12832 17382
rect 12856 17380 12912 17382
rect 12616 16346 12672 16348
rect 12696 16346 12752 16348
rect 12776 16346 12832 16348
rect 12856 16346 12912 16348
rect 12616 16294 12662 16346
rect 12662 16294 12672 16346
rect 12696 16294 12726 16346
rect 12726 16294 12738 16346
rect 12738 16294 12752 16346
rect 12776 16294 12790 16346
rect 12790 16294 12802 16346
rect 12802 16294 12832 16346
rect 12856 16294 12866 16346
rect 12866 16294 12912 16346
rect 12616 16292 12672 16294
rect 12696 16292 12752 16294
rect 12776 16292 12832 16294
rect 12856 16292 12912 16294
rect 12616 15258 12672 15260
rect 12696 15258 12752 15260
rect 12776 15258 12832 15260
rect 12856 15258 12912 15260
rect 12616 15206 12662 15258
rect 12662 15206 12672 15258
rect 12696 15206 12726 15258
rect 12726 15206 12738 15258
rect 12738 15206 12752 15258
rect 12776 15206 12790 15258
rect 12790 15206 12802 15258
rect 12802 15206 12832 15258
rect 12856 15206 12866 15258
rect 12866 15206 12912 15258
rect 12616 15204 12672 15206
rect 12696 15204 12752 15206
rect 12776 15204 12832 15206
rect 12856 15204 12912 15206
rect 12616 14170 12672 14172
rect 12696 14170 12752 14172
rect 12776 14170 12832 14172
rect 12856 14170 12912 14172
rect 12616 14118 12662 14170
rect 12662 14118 12672 14170
rect 12696 14118 12726 14170
rect 12726 14118 12738 14170
rect 12738 14118 12752 14170
rect 12776 14118 12790 14170
rect 12790 14118 12802 14170
rect 12802 14118 12832 14170
rect 12856 14118 12866 14170
rect 12866 14118 12912 14170
rect 12616 14116 12672 14118
rect 12696 14116 12752 14118
rect 12776 14116 12832 14118
rect 12856 14116 12912 14118
rect 12616 13082 12672 13084
rect 12696 13082 12752 13084
rect 12776 13082 12832 13084
rect 12856 13082 12912 13084
rect 12616 13030 12662 13082
rect 12662 13030 12672 13082
rect 12696 13030 12726 13082
rect 12726 13030 12738 13082
rect 12738 13030 12752 13082
rect 12776 13030 12790 13082
rect 12790 13030 12802 13082
rect 12802 13030 12832 13082
rect 12856 13030 12866 13082
rect 12866 13030 12912 13082
rect 12616 13028 12672 13030
rect 12696 13028 12752 13030
rect 12776 13028 12832 13030
rect 12856 13028 12912 13030
rect 12616 11994 12672 11996
rect 12696 11994 12752 11996
rect 12776 11994 12832 11996
rect 12856 11994 12912 11996
rect 12616 11942 12662 11994
rect 12662 11942 12672 11994
rect 12696 11942 12726 11994
rect 12726 11942 12738 11994
rect 12738 11942 12752 11994
rect 12776 11942 12790 11994
rect 12790 11942 12802 11994
rect 12802 11942 12832 11994
rect 12856 11942 12866 11994
rect 12866 11942 12912 11994
rect 12616 11940 12672 11942
rect 12696 11940 12752 11942
rect 12776 11940 12832 11942
rect 12856 11940 12912 11942
rect 12616 10906 12672 10908
rect 12696 10906 12752 10908
rect 12776 10906 12832 10908
rect 12856 10906 12912 10908
rect 12616 10854 12662 10906
rect 12662 10854 12672 10906
rect 12696 10854 12726 10906
rect 12726 10854 12738 10906
rect 12738 10854 12752 10906
rect 12776 10854 12790 10906
rect 12790 10854 12802 10906
rect 12802 10854 12832 10906
rect 12856 10854 12866 10906
rect 12866 10854 12912 10906
rect 12616 10852 12672 10854
rect 12696 10852 12752 10854
rect 12776 10852 12832 10854
rect 12856 10852 12912 10854
rect 12616 9818 12672 9820
rect 12696 9818 12752 9820
rect 12776 9818 12832 9820
rect 12856 9818 12912 9820
rect 12616 9766 12662 9818
rect 12662 9766 12672 9818
rect 12696 9766 12726 9818
rect 12726 9766 12738 9818
rect 12738 9766 12752 9818
rect 12776 9766 12790 9818
rect 12790 9766 12802 9818
rect 12802 9766 12832 9818
rect 12856 9766 12866 9818
rect 12866 9766 12912 9818
rect 12616 9764 12672 9766
rect 12696 9764 12752 9766
rect 12776 9764 12832 9766
rect 12856 9764 12912 9766
rect 12616 8730 12672 8732
rect 12696 8730 12752 8732
rect 12776 8730 12832 8732
rect 12856 8730 12912 8732
rect 12616 8678 12662 8730
rect 12662 8678 12672 8730
rect 12696 8678 12726 8730
rect 12726 8678 12738 8730
rect 12738 8678 12752 8730
rect 12776 8678 12790 8730
rect 12790 8678 12802 8730
rect 12802 8678 12832 8730
rect 12856 8678 12866 8730
rect 12866 8678 12912 8730
rect 12616 8676 12672 8678
rect 12696 8676 12752 8678
rect 12776 8676 12832 8678
rect 12856 8676 12912 8678
rect 12616 7642 12672 7644
rect 12696 7642 12752 7644
rect 12776 7642 12832 7644
rect 12856 7642 12912 7644
rect 12616 7590 12662 7642
rect 12662 7590 12672 7642
rect 12696 7590 12726 7642
rect 12726 7590 12738 7642
rect 12738 7590 12752 7642
rect 12776 7590 12790 7642
rect 12790 7590 12802 7642
rect 12802 7590 12832 7642
rect 12856 7590 12866 7642
rect 12866 7590 12912 7642
rect 12616 7588 12672 7590
rect 12696 7588 12752 7590
rect 12776 7588 12832 7590
rect 12856 7588 12912 7590
rect 12616 6554 12672 6556
rect 12696 6554 12752 6556
rect 12776 6554 12832 6556
rect 12856 6554 12912 6556
rect 12616 6502 12662 6554
rect 12662 6502 12672 6554
rect 12696 6502 12726 6554
rect 12726 6502 12738 6554
rect 12738 6502 12752 6554
rect 12776 6502 12790 6554
rect 12790 6502 12802 6554
rect 12802 6502 12832 6554
rect 12856 6502 12866 6554
rect 12866 6502 12912 6554
rect 12616 6500 12672 6502
rect 12696 6500 12752 6502
rect 12776 6500 12832 6502
rect 12856 6500 12912 6502
rect 12616 5466 12672 5468
rect 12696 5466 12752 5468
rect 12776 5466 12832 5468
rect 12856 5466 12912 5468
rect 12616 5414 12662 5466
rect 12662 5414 12672 5466
rect 12696 5414 12726 5466
rect 12726 5414 12738 5466
rect 12738 5414 12752 5466
rect 12776 5414 12790 5466
rect 12790 5414 12802 5466
rect 12802 5414 12832 5466
rect 12856 5414 12866 5466
rect 12866 5414 12912 5466
rect 12616 5412 12672 5414
rect 12696 5412 12752 5414
rect 12776 5412 12832 5414
rect 12856 5412 12912 5414
rect 12616 4378 12672 4380
rect 12696 4378 12752 4380
rect 12776 4378 12832 4380
rect 12856 4378 12912 4380
rect 12616 4326 12662 4378
rect 12662 4326 12672 4378
rect 12696 4326 12726 4378
rect 12726 4326 12738 4378
rect 12738 4326 12752 4378
rect 12776 4326 12790 4378
rect 12790 4326 12802 4378
rect 12802 4326 12832 4378
rect 12856 4326 12866 4378
rect 12866 4326 12912 4378
rect 12616 4324 12672 4326
rect 12696 4324 12752 4326
rect 12776 4324 12832 4326
rect 12856 4324 12912 4326
rect 11956 3834 12012 3836
rect 12036 3834 12092 3836
rect 12116 3834 12172 3836
rect 12196 3834 12252 3836
rect 11956 3782 12002 3834
rect 12002 3782 12012 3834
rect 12036 3782 12066 3834
rect 12066 3782 12078 3834
rect 12078 3782 12092 3834
rect 12116 3782 12130 3834
rect 12130 3782 12142 3834
rect 12142 3782 12172 3834
rect 12196 3782 12206 3834
rect 12206 3782 12252 3834
rect 11956 3780 12012 3782
rect 12036 3780 12092 3782
rect 12116 3780 12172 3782
rect 12196 3780 12252 3782
rect 14554 45892 14610 45928
rect 14554 45872 14556 45892
rect 14556 45872 14608 45892
rect 14608 45872 14610 45892
rect 12616 3290 12672 3292
rect 12696 3290 12752 3292
rect 12776 3290 12832 3292
rect 12856 3290 12912 3292
rect 12616 3238 12662 3290
rect 12662 3238 12672 3290
rect 12696 3238 12726 3290
rect 12726 3238 12738 3290
rect 12738 3238 12752 3290
rect 12776 3238 12790 3290
rect 12790 3238 12802 3290
rect 12802 3238 12832 3290
rect 12856 3238 12866 3290
rect 12866 3238 12912 3290
rect 12616 3236 12672 3238
rect 12696 3236 12752 3238
rect 12776 3236 12832 3238
rect 12856 3236 12912 3238
rect 11956 2746 12012 2748
rect 12036 2746 12092 2748
rect 12116 2746 12172 2748
rect 12196 2746 12252 2748
rect 11956 2694 12002 2746
rect 12002 2694 12012 2746
rect 12036 2694 12066 2746
rect 12066 2694 12078 2746
rect 12078 2694 12092 2746
rect 12116 2694 12130 2746
rect 12130 2694 12142 2746
rect 12142 2694 12172 2746
rect 12196 2694 12206 2746
rect 12206 2694 12252 2746
rect 11956 2692 12012 2694
rect 12036 2692 12092 2694
rect 12116 2692 12172 2694
rect 12196 2692 12252 2694
rect 16956 69114 17012 69116
rect 17036 69114 17092 69116
rect 17116 69114 17172 69116
rect 17196 69114 17252 69116
rect 16956 69062 17002 69114
rect 17002 69062 17012 69114
rect 17036 69062 17066 69114
rect 17066 69062 17078 69114
rect 17078 69062 17092 69114
rect 17116 69062 17130 69114
rect 17130 69062 17142 69114
rect 17142 69062 17172 69114
rect 17196 69062 17206 69114
rect 17206 69062 17252 69114
rect 16956 69060 17012 69062
rect 17036 69060 17092 69062
rect 17116 69060 17172 69062
rect 17196 69060 17252 69062
rect 17616 68570 17672 68572
rect 17696 68570 17752 68572
rect 17776 68570 17832 68572
rect 17856 68570 17912 68572
rect 17616 68518 17662 68570
rect 17662 68518 17672 68570
rect 17696 68518 17726 68570
rect 17726 68518 17738 68570
rect 17738 68518 17752 68570
rect 17776 68518 17790 68570
rect 17790 68518 17802 68570
rect 17802 68518 17832 68570
rect 17856 68518 17866 68570
rect 17866 68518 17912 68570
rect 17616 68516 17672 68518
rect 17696 68516 17752 68518
rect 17776 68516 17832 68518
rect 17856 68516 17912 68518
rect 16956 68026 17012 68028
rect 17036 68026 17092 68028
rect 17116 68026 17172 68028
rect 17196 68026 17252 68028
rect 16956 67974 17002 68026
rect 17002 67974 17012 68026
rect 17036 67974 17066 68026
rect 17066 67974 17078 68026
rect 17078 67974 17092 68026
rect 17116 67974 17130 68026
rect 17130 67974 17142 68026
rect 17142 67974 17172 68026
rect 17196 67974 17206 68026
rect 17206 67974 17252 68026
rect 16956 67972 17012 67974
rect 17036 67972 17092 67974
rect 17116 67972 17172 67974
rect 17196 67972 17252 67974
rect 17616 67482 17672 67484
rect 17696 67482 17752 67484
rect 17776 67482 17832 67484
rect 17856 67482 17912 67484
rect 17616 67430 17662 67482
rect 17662 67430 17672 67482
rect 17696 67430 17726 67482
rect 17726 67430 17738 67482
rect 17738 67430 17752 67482
rect 17776 67430 17790 67482
rect 17790 67430 17802 67482
rect 17802 67430 17832 67482
rect 17856 67430 17866 67482
rect 17866 67430 17912 67482
rect 17616 67428 17672 67430
rect 17696 67428 17752 67430
rect 17776 67428 17832 67430
rect 17856 67428 17912 67430
rect 16956 66938 17012 66940
rect 17036 66938 17092 66940
rect 17116 66938 17172 66940
rect 17196 66938 17252 66940
rect 16956 66886 17002 66938
rect 17002 66886 17012 66938
rect 17036 66886 17066 66938
rect 17066 66886 17078 66938
rect 17078 66886 17092 66938
rect 17116 66886 17130 66938
rect 17130 66886 17142 66938
rect 17142 66886 17172 66938
rect 17196 66886 17206 66938
rect 17206 66886 17252 66938
rect 16956 66884 17012 66886
rect 17036 66884 17092 66886
rect 17116 66884 17172 66886
rect 17196 66884 17252 66886
rect 16956 65850 17012 65852
rect 17036 65850 17092 65852
rect 17116 65850 17172 65852
rect 17196 65850 17252 65852
rect 16956 65798 17002 65850
rect 17002 65798 17012 65850
rect 17036 65798 17066 65850
rect 17066 65798 17078 65850
rect 17078 65798 17092 65850
rect 17116 65798 17130 65850
rect 17130 65798 17142 65850
rect 17142 65798 17172 65850
rect 17196 65798 17206 65850
rect 17206 65798 17252 65850
rect 16956 65796 17012 65798
rect 17036 65796 17092 65798
rect 17116 65796 17172 65798
rect 17196 65796 17252 65798
rect 16956 64762 17012 64764
rect 17036 64762 17092 64764
rect 17116 64762 17172 64764
rect 17196 64762 17252 64764
rect 16956 64710 17002 64762
rect 17002 64710 17012 64762
rect 17036 64710 17066 64762
rect 17066 64710 17078 64762
rect 17078 64710 17092 64762
rect 17116 64710 17130 64762
rect 17130 64710 17142 64762
rect 17142 64710 17172 64762
rect 17196 64710 17206 64762
rect 17206 64710 17252 64762
rect 16956 64708 17012 64710
rect 17036 64708 17092 64710
rect 17116 64708 17172 64710
rect 17196 64708 17252 64710
rect 16956 63674 17012 63676
rect 17036 63674 17092 63676
rect 17116 63674 17172 63676
rect 17196 63674 17252 63676
rect 16956 63622 17002 63674
rect 17002 63622 17012 63674
rect 17036 63622 17066 63674
rect 17066 63622 17078 63674
rect 17078 63622 17092 63674
rect 17116 63622 17130 63674
rect 17130 63622 17142 63674
rect 17142 63622 17172 63674
rect 17196 63622 17206 63674
rect 17206 63622 17252 63674
rect 16956 63620 17012 63622
rect 17036 63620 17092 63622
rect 17116 63620 17172 63622
rect 17196 63620 17252 63622
rect 16956 62586 17012 62588
rect 17036 62586 17092 62588
rect 17116 62586 17172 62588
rect 17196 62586 17252 62588
rect 16956 62534 17002 62586
rect 17002 62534 17012 62586
rect 17036 62534 17066 62586
rect 17066 62534 17078 62586
rect 17078 62534 17092 62586
rect 17116 62534 17130 62586
rect 17130 62534 17142 62586
rect 17142 62534 17172 62586
rect 17196 62534 17206 62586
rect 17206 62534 17252 62586
rect 16956 62532 17012 62534
rect 17036 62532 17092 62534
rect 17116 62532 17172 62534
rect 17196 62532 17252 62534
rect 16956 61498 17012 61500
rect 17036 61498 17092 61500
rect 17116 61498 17172 61500
rect 17196 61498 17252 61500
rect 16956 61446 17002 61498
rect 17002 61446 17012 61498
rect 17036 61446 17066 61498
rect 17066 61446 17078 61498
rect 17078 61446 17092 61498
rect 17116 61446 17130 61498
rect 17130 61446 17142 61498
rect 17142 61446 17172 61498
rect 17196 61446 17206 61498
rect 17206 61446 17252 61498
rect 16956 61444 17012 61446
rect 17036 61444 17092 61446
rect 17116 61444 17172 61446
rect 17196 61444 17252 61446
rect 16956 60410 17012 60412
rect 17036 60410 17092 60412
rect 17116 60410 17172 60412
rect 17196 60410 17252 60412
rect 16956 60358 17002 60410
rect 17002 60358 17012 60410
rect 17036 60358 17066 60410
rect 17066 60358 17078 60410
rect 17078 60358 17092 60410
rect 17116 60358 17130 60410
rect 17130 60358 17142 60410
rect 17142 60358 17172 60410
rect 17196 60358 17206 60410
rect 17206 60358 17252 60410
rect 16956 60356 17012 60358
rect 17036 60356 17092 60358
rect 17116 60356 17172 60358
rect 17196 60356 17252 60358
rect 16956 59322 17012 59324
rect 17036 59322 17092 59324
rect 17116 59322 17172 59324
rect 17196 59322 17252 59324
rect 16956 59270 17002 59322
rect 17002 59270 17012 59322
rect 17036 59270 17066 59322
rect 17066 59270 17078 59322
rect 17078 59270 17092 59322
rect 17116 59270 17130 59322
rect 17130 59270 17142 59322
rect 17142 59270 17172 59322
rect 17196 59270 17206 59322
rect 17206 59270 17252 59322
rect 16956 59268 17012 59270
rect 17036 59268 17092 59270
rect 17116 59268 17172 59270
rect 17196 59268 17252 59270
rect 16956 58234 17012 58236
rect 17036 58234 17092 58236
rect 17116 58234 17172 58236
rect 17196 58234 17252 58236
rect 16956 58182 17002 58234
rect 17002 58182 17012 58234
rect 17036 58182 17066 58234
rect 17066 58182 17078 58234
rect 17078 58182 17092 58234
rect 17116 58182 17130 58234
rect 17130 58182 17142 58234
rect 17142 58182 17172 58234
rect 17196 58182 17206 58234
rect 17206 58182 17252 58234
rect 16956 58180 17012 58182
rect 17036 58180 17092 58182
rect 17116 58180 17172 58182
rect 17196 58180 17252 58182
rect 16956 57146 17012 57148
rect 17036 57146 17092 57148
rect 17116 57146 17172 57148
rect 17196 57146 17252 57148
rect 16956 57094 17002 57146
rect 17002 57094 17012 57146
rect 17036 57094 17066 57146
rect 17066 57094 17078 57146
rect 17078 57094 17092 57146
rect 17116 57094 17130 57146
rect 17130 57094 17142 57146
rect 17142 57094 17172 57146
rect 17196 57094 17206 57146
rect 17206 57094 17252 57146
rect 16956 57092 17012 57094
rect 17036 57092 17092 57094
rect 17116 57092 17172 57094
rect 17196 57092 17252 57094
rect 16956 56058 17012 56060
rect 17036 56058 17092 56060
rect 17116 56058 17172 56060
rect 17196 56058 17252 56060
rect 16956 56006 17002 56058
rect 17002 56006 17012 56058
rect 17036 56006 17066 56058
rect 17066 56006 17078 56058
rect 17078 56006 17092 56058
rect 17116 56006 17130 56058
rect 17130 56006 17142 56058
rect 17142 56006 17172 56058
rect 17196 56006 17206 56058
rect 17206 56006 17252 56058
rect 16956 56004 17012 56006
rect 17036 56004 17092 56006
rect 17116 56004 17172 56006
rect 17196 56004 17252 56006
rect 16956 54970 17012 54972
rect 17036 54970 17092 54972
rect 17116 54970 17172 54972
rect 17196 54970 17252 54972
rect 16956 54918 17002 54970
rect 17002 54918 17012 54970
rect 17036 54918 17066 54970
rect 17066 54918 17078 54970
rect 17078 54918 17092 54970
rect 17116 54918 17130 54970
rect 17130 54918 17142 54970
rect 17142 54918 17172 54970
rect 17196 54918 17206 54970
rect 17206 54918 17252 54970
rect 16956 54916 17012 54918
rect 17036 54916 17092 54918
rect 17116 54916 17172 54918
rect 17196 54916 17252 54918
rect 16956 53882 17012 53884
rect 17036 53882 17092 53884
rect 17116 53882 17172 53884
rect 17196 53882 17252 53884
rect 16956 53830 17002 53882
rect 17002 53830 17012 53882
rect 17036 53830 17066 53882
rect 17066 53830 17078 53882
rect 17078 53830 17092 53882
rect 17116 53830 17130 53882
rect 17130 53830 17142 53882
rect 17142 53830 17172 53882
rect 17196 53830 17206 53882
rect 17206 53830 17252 53882
rect 16956 53828 17012 53830
rect 17036 53828 17092 53830
rect 17116 53828 17172 53830
rect 17196 53828 17252 53830
rect 17616 66394 17672 66396
rect 17696 66394 17752 66396
rect 17776 66394 17832 66396
rect 17856 66394 17912 66396
rect 17616 66342 17662 66394
rect 17662 66342 17672 66394
rect 17696 66342 17726 66394
rect 17726 66342 17738 66394
rect 17738 66342 17752 66394
rect 17776 66342 17790 66394
rect 17790 66342 17802 66394
rect 17802 66342 17832 66394
rect 17856 66342 17866 66394
rect 17866 66342 17912 66394
rect 17616 66340 17672 66342
rect 17696 66340 17752 66342
rect 17776 66340 17832 66342
rect 17856 66340 17912 66342
rect 17616 65306 17672 65308
rect 17696 65306 17752 65308
rect 17776 65306 17832 65308
rect 17856 65306 17912 65308
rect 17616 65254 17662 65306
rect 17662 65254 17672 65306
rect 17696 65254 17726 65306
rect 17726 65254 17738 65306
rect 17738 65254 17752 65306
rect 17776 65254 17790 65306
rect 17790 65254 17802 65306
rect 17802 65254 17832 65306
rect 17856 65254 17866 65306
rect 17866 65254 17912 65306
rect 17616 65252 17672 65254
rect 17696 65252 17752 65254
rect 17776 65252 17832 65254
rect 17856 65252 17912 65254
rect 16956 52794 17012 52796
rect 17036 52794 17092 52796
rect 17116 52794 17172 52796
rect 17196 52794 17252 52796
rect 16956 52742 17002 52794
rect 17002 52742 17012 52794
rect 17036 52742 17066 52794
rect 17066 52742 17078 52794
rect 17078 52742 17092 52794
rect 17116 52742 17130 52794
rect 17130 52742 17142 52794
rect 17142 52742 17172 52794
rect 17196 52742 17206 52794
rect 17206 52742 17252 52794
rect 16956 52740 17012 52742
rect 17036 52740 17092 52742
rect 17116 52740 17172 52742
rect 17196 52740 17252 52742
rect 16956 51706 17012 51708
rect 17036 51706 17092 51708
rect 17116 51706 17172 51708
rect 17196 51706 17252 51708
rect 16956 51654 17002 51706
rect 17002 51654 17012 51706
rect 17036 51654 17066 51706
rect 17066 51654 17078 51706
rect 17078 51654 17092 51706
rect 17116 51654 17130 51706
rect 17130 51654 17142 51706
rect 17142 51654 17172 51706
rect 17196 51654 17206 51706
rect 17206 51654 17252 51706
rect 16956 51652 17012 51654
rect 17036 51652 17092 51654
rect 17116 51652 17172 51654
rect 17196 51652 17252 51654
rect 16956 50618 17012 50620
rect 17036 50618 17092 50620
rect 17116 50618 17172 50620
rect 17196 50618 17252 50620
rect 16956 50566 17002 50618
rect 17002 50566 17012 50618
rect 17036 50566 17066 50618
rect 17066 50566 17078 50618
rect 17078 50566 17092 50618
rect 17116 50566 17130 50618
rect 17130 50566 17142 50618
rect 17142 50566 17172 50618
rect 17196 50566 17206 50618
rect 17206 50566 17252 50618
rect 16956 50564 17012 50566
rect 17036 50564 17092 50566
rect 17116 50564 17172 50566
rect 17196 50564 17252 50566
rect 16956 49530 17012 49532
rect 17036 49530 17092 49532
rect 17116 49530 17172 49532
rect 17196 49530 17252 49532
rect 16956 49478 17002 49530
rect 17002 49478 17012 49530
rect 17036 49478 17066 49530
rect 17066 49478 17078 49530
rect 17078 49478 17092 49530
rect 17116 49478 17130 49530
rect 17130 49478 17142 49530
rect 17142 49478 17172 49530
rect 17196 49478 17206 49530
rect 17206 49478 17252 49530
rect 16956 49476 17012 49478
rect 17036 49476 17092 49478
rect 17116 49476 17172 49478
rect 17196 49476 17252 49478
rect 16956 48442 17012 48444
rect 17036 48442 17092 48444
rect 17116 48442 17172 48444
rect 17196 48442 17252 48444
rect 16956 48390 17002 48442
rect 17002 48390 17012 48442
rect 17036 48390 17066 48442
rect 17066 48390 17078 48442
rect 17078 48390 17092 48442
rect 17116 48390 17130 48442
rect 17130 48390 17142 48442
rect 17142 48390 17172 48442
rect 17196 48390 17206 48442
rect 17206 48390 17252 48442
rect 16956 48388 17012 48390
rect 17036 48388 17092 48390
rect 17116 48388 17172 48390
rect 17196 48388 17252 48390
rect 16956 47354 17012 47356
rect 17036 47354 17092 47356
rect 17116 47354 17172 47356
rect 17196 47354 17252 47356
rect 16956 47302 17002 47354
rect 17002 47302 17012 47354
rect 17036 47302 17066 47354
rect 17066 47302 17078 47354
rect 17078 47302 17092 47354
rect 17116 47302 17130 47354
rect 17130 47302 17142 47354
rect 17142 47302 17172 47354
rect 17196 47302 17206 47354
rect 17206 47302 17252 47354
rect 16956 47300 17012 47302
rect 17036 47300 17092 47302
rect 17116 47300 17172 47302
rect 17196 47300 17252 47302
rect 16956 46266 17012 46268
rect 17036 46266 17092 46268
rect 17116 46266 17172 46268
rect 17196 46266 17252 46268
rect 16956 46214 17002 46266
rect 17002 46214 17012 46266
rect 17036 46214 17066 46266
rect 17066 46214 17078 46266
rect 17078 46214 17092 46266
rect 17116 46214 17130 46266
rect 17130 46214 17142 46266
rect 17142 46214 17172 46266
rect 17196 46214 17206 46266
rect 17206 46214 17252 46266
rect 16956 46212 17012 46214
rect 17036 46212 17092 46214
rect 17116 46212 17172 46214
rect 17196 46212 17252 46214
rect 16956 45178 17012 45180
rect 17036 45178 17092 45180
rect 17116 45178 17172 45180
rect 17196 45178 17252 45180
rect 16956 45126 17002 45178
rect 17002 45126 17012 45178
rect 17036 45126 17066 45178
rect 17066 45126 17078 45178
rect 17078 45126 17092 45178
rect 17116 45126 17130 45178
rect 17130 45126 17142 45178
rect 17142 45126 17172 45178
rect 17196 45126 17206 45178
rect 17206 45126 17252 45178
rect 16956 45124 17012 45126
rect 17036 45124 17092 45126
rect 17116 45124 17172 45126
rect 17196 45124 17252 45126
rect 16956 44090 17012 44092
rect 17036 44090 17092 44092
rect 17116 44090 17172 44092
rect 17196 44090 17252 44092
rect 16956 44038 17002 44090
rect 17002 44038 17012 44090
rect 17036 44038 17066 44090
rect 17066 44038 17078 44090
rect 17078 44038 17092 44090
rect 17116 44038 17130 44090
rect 17130 44038 17142 44090
rect 17142 44038 17172 44090
rect 17196 44038 17206 44090
rect 17206 44038 17252 44090
rect 16956 44036 17012 44038
rect 17036 44036 17092 44038
rect 17116 44036 17172 44038
rect 17196 44036 17252 44038
rect 16956 43002 17012 43004
rect 17036 43002 17092 43004
rect 17116 43002 17172 43004
rect 17196 43002 17252 43004
rect 16956 42950 17002 43002
rect 17002 42950 17012 43002
rect 17036 42950 17066 43002
rect 17066 42950 17078 43002
rect 17078 42950 17092 43002
rect 17116 42950 17130 43002
rect 17130 42950 17142 43002
rect 17142 42950 17172 43002
rect 17196 42950 17206 43002
rect 17206 42950 17252 43002
rect 16956 42948 17012 42950
rect 17036 42948 17092 42950
rect 17116 42948 17172 42950
rect 17196 42948 17252 42950
rect 16956 41914 17012 41916
rect 17036 41914 17092 41916
rect 17116 41914 17172 41916
rect 17196 41914 17252 41916
rect 16956 41862 17002 41914
rect 17002 41862 17012 41914
rect 17036 41862 17066 41914
rect 17066 41862 17078 41914
rect 17078 41862 17092 41914
rect 17116 41862 17130 41914
rect 17130 41862 17142 41914
rect 17142 41862 17172 41914
rect 17196 41862 17206 41914
rect 17206 41862 17252 41914
rect 16956 41860 17012 41862
rect 17036 41860 17092 41862
rect 17116 41860 17172 41862
rect 17196 41860 17252 41862
rect 16956 40826 17012 40828
rect 17036 40826 17092 40828
rect 17116 40826 17172 40828
rect 17196 40826 17252 40828
rect 16956 40774 17002 40826
rect 17002 40774 17012 40826
rect 17036 40774 17066 40826
rect 17066 40774 17078 40826
rect 17078 40774 17092 40826
rect 17116 40774 17130 40826
rect 17130 40774 17142 40826
rect 17142 40774 17172 40826
rect 17196 40774 17206 40826
rect 17206 40774 17252 40826
rect 16956 40772 17012 40774
rect 17036 40772 17092 40774
rect 17116 40772 17172 40774
rect 17196 40772 17252 40774
rect 16956 39738 17012 39740
rect 17036 39738 17092 39740
rect 17116 39738 17172 39740
rect 17196 39738 17252 39740
rect 16956 39686 17002 39738
rect 17002 39686 17012 39738
rect 17036 39686 17066 39738
rect 17066 39686 17078 39738
rect 17078 39686 17092 39738
rect 17116 39686 17130 39738
rect 17130 39686 17142 39738
rect 17142 39686 17172 39738
rect 17196 39686 17206 39738
rect 17206 39686 17252 39738
rect 16956 39684 17012 39686
rect 17036 39684 17092 39686
rect 17116 39684 17172 39686
rect 17196 39684 17252 39686
rect 16956 38650 17012 38652
rect 17036 38650 17092 38652
rect 17116 38650 17172 38652
rect 17196 38650 17252 38652
rect 16956 38598 17002 38650
rect 17002 38598 17012 38650
rect 17036 38598 17066 38650
rect 17066 38598 17078 38650
rect 17078 38598 17092 38650
rect 17116 38598 17130 38650
rect 17130 38598 17142 38650
rect 17142 38598 17172 38650
rect 17196 38598 17206 38650
rect 17206 38598 17252 38650
rect 16956 38596 17012 38598
rect 17036 38596 17092 38598
rect 17116 38596 17172 38598
rect 17196 38596 17252 38598
rect 16956 37562 17012 37564
rect 17036 37562 17092 37564
rect 17116 37562 17172 37564
rect 17196 37562 17252 37564
rect 16956 37510 17002 37562
rect 17002 37510 17012 37562
rect 17036 37510 17066 37562
rect 17066 37510 17078 37562
rect 17078 37510 17092 37562
rect 17116 37510 17130 37562
rect 17130 37510 17142 37562
rect 17142 37510 17172 37562
rect 17196 37510 17206 37562
rect 17206 37510 17252 37562
rect 16956 37508 17012 37510
rect 17036 37508 17092 37510
rect 17116 37508 17172 37510
rect 17196 37508 17252 37510
rect 16956 36474 17012 36476
rect 17036 36474 17092 36476
rect 17116 36474 17172 36476
rect 17196 36474 17252 36476
rect 16956 36422 17002 36474
rect 17002 36422 17012 36474
rect 17036 36422 17066 36474
rect 17066 36422 17078 36474
rect 17078 36422 17092 36474
rect 17116 36422 17130 36474
rect 17130 36422 17142 36474
rect 17142 36422 17172 36474
rect 17196 36422 17206 36474
rect 17206 36422 17252 36474
rect 16956 36420 17012 36422
rect 17036 36420 17092 36422
rect 17116 36420 17172 36422
rect 17196 36420 17252 36422
rect 16956 35386 17012 35388
rect 17036 35386 17092 35388
rect 17116 35386 17172 35388
rect 17196 35386 17252 35388
rect 16956 35334 17002 35386
rect 17002 35334 17012 35386
rect 17036 35334 17066 35386
rect 17066 35334 17078 35386
rect 17078 35334 17092 35386
rect 17116 35334 17130 35386
rect 17130 35334 17142 35386
rect 17142 35334 17172 35386
rect 17196 35334 17206 35386
rect 17206 35334 17252 35386
rect 16956 35332 17012 35334
rect 17036 35332 17092 35334
rect 17116 35332 17172 35334
rect 17196 35332 17252 35334
rect 16956 34298 17012 34300
rect 17036 34298 17092 34300
rect 17116 34298 17172 34300
rect 17196 34298 17252 34300
rect 16956 34246 17002 34298
rect 17002 34246 17012 34298
rect 17036 34246 17066 34298
rect 17066 34246 17078 34298
rect 17078 34246 17092 34298
rect 17116 34246 17130 34298
rect 17130 34246 17142 34298
rect 17142 34246 17172 34298
rect 17196 34246 17206 34298
rect 17206 34246 17252 34298
rect 16956 34244 17012 34246
rect 17036 34244 17092 34246
rect 17116 34244 17172 34246
rect 17196 34244 17252 34246
rect 16956 33210 17012 33212
rect 17036 33210 17092 33212
rect 17116 33210 17172 33212
rect 17196 33210 17252 33212
rect 16956 33158 17002 33210
rect 17002 33158 17012 33210
rect 17036 33158 17066 33210
rect 17066 33158 17078 33210
rect 17078 33158 17092 33210
rect 17116 33158 17130 33210
rect 17130 33158 17142 33210
rect 17142 33158 17172 33210
rect 17196 33158 17206 33210
rect 17206 33158 17252 33210
rect 16956 33156 17012 33158
rect 17036 33156 17092 33158
rect 17116 33156 17172 33158
rect 17196 33156 17252 33158
rect 16956 32122 17012 32124
rect 17036 32122 17092 32124
rect 17116 32122 17172 32124
rect 17196 32122 17252 32124
rect 16956 32070 17002 32122
rect 17002 32070 17012 32122
rect 17036 32070 17066 32122
rect 17066 32070 17078 32122
rect 17078 32070 17092 32122
rect 17116 32070 17130 32122
rect 17130 32070 17142 32122
rect 17142 32070 17172 32122
rect 17196 32070 17206 32122
rect 17206 32070 17252 32122
rect 16956 32068 17012 32070
rect 17036 32068 17092 32070
rect 17116 32068 17172 32070
rect 17196 32068 17252 32070
rect 16956 31034 17012 31036
rect 17036 31034 17092 31036
rect 17116 31034 17172 31036
rect 17196 31034 17252 31036
rect 16956 30982 17002 31034
rect 17002 30982 17012 31034
rect 17036 30982 17066 31034
rect 17066 30982 17078 31034
rect 17078 30982 17092 31034
rect 17116 30982 17130 31034
rect 17130 30982 17142 31034
rect 17142 30982 17172 31034
rect 17196 30982 17206 31034
rect 17206 30982 17252 31034
rect 16956 30980 17012 30982
rect 17036 30980 17092 30982
rect 17116 30980 17172 30982
rect 17196 30980 17252 30982
rect 16956 29946 17012 29948
rect 17036 29946 17092 29948
rect 17116 29946 17172 29948
rect 17196 29946 17252 29948
rect 16956 29894 17002 29946
rect 17002 29894 17012 29946
rect 17036 29894 17066 29946
rect 17066 29894 17078 29946
rect 17078 29894 17092 29946
rect 17116 29894 17130 29946
rect 17130 29894 17142 29946
rect 17142 29894 17172 29946
rect 17196 29894 17206 29946
rect 17206 29894 17252 29946
rect 16956 29892 17012 29894
rect 17036 29892 17092 29894
rect 17116 29892 17172 29894
rect 17196 29892 17252 29894
rect 16956 28858 17012 28860
rect 17036 28858 17092 28860
rect 17116 28858 17172 28860
rect 17196 28858 17252 28860
rect 16956 28806 17002 28858
rect 17002 28806 17012 28858
rect 17036 28806 17066 28858
rect 17066 28806 17078 28858
rect 17078 28806 17092 28858
rect 17116 28806 17130 28858
rect 17130 28806 17142 28858
rect 17142 28806 17172 28858
rect 17196 28806 17206 28858
rect 17206 28806 17252 28858
rect 16956 28804 17012 28806
rect 17036 28804 17092 28806
rect 17116 28804 17172 28806
rect 17196 28804 17252 28806
rect 16956 27770 17012 27772
rect 17036 27770 17092 27772
rect 17116 27770 17172 27772
rect 17196 27770 17252 27772
rect 16956 27718 17002 27770
rect 17002 27718 17012 27770
rect 17036 27718 17066 27770
rect 17066 27718 17078 27770
rect 17078 27718 17092 27770
rect 17116 27718 17130 27770
rect 17130 27718 17142 27770
rect 17142 27718 17172 27770
rect 17196 27718 17206 27770
rect 17206 27718 17252 27770
rect 16956 27716 17012 27718
rect 17036 27716 17092 27718
rect 17116 27716 17172 27718
rect 17196 27716 17252 27718
rect 16956 26682 17012 26684
rect 17036 26682 17092 26684
rect 17116 26682 17172 26684
rect 17196 26682 17252 26684
rect 16956 26630 17002 26682
rect 17002 26630 17012 26682
rect 17036 26630 17066 26682
rect 17066 26630 17078 26682
rect 17078 26630 17092 26682
rect 17116 26630 17130 26682
rect 17130 26630 17142 26682
rect 17142 26630 17172 26682
rect 17196 26630 17206 26682
rect 17206 26630 17252 26682
rect 16956 26628 17012 26630
rect 17036 26628 17092 26630
rect 17116 26628 17172 26630
rect 17196 26628 17252 26630
rect 16956 25594 17012 25596
rect 17036 25594 17092 25596
rect 17116 25594 17172 25596
rect 17196 25594 17252 25596
rect 16956 25542 17002 25594
rect 17002 25542 17012 25594
rect 17036 25542 17066 25594
rect 17066 25542 17078 25594
rect 17078 25542 17092 25594
rect 17116 25542 17130 25594
rect 17130 25542 17142 25594
rect 17142 25542 17172 25594
rect 17196 25542 17206 25594
rect 17206 25542 17252 25594
rect 16956 25540 17012 25542
rect 17036 25540 17092 25542
rect 17116 25540 17172 25542
rect 17196 25540 17252 25542
rect 16956 24506 17012 24508
rect 17036 24506 17092 24508
rect 17116 24506 17172 24508
rect 17196 24506 17252 24508
rect 16956 24454 17002 24506
rect 17002 24454 17012 24506
rect 17036 24454 17066 24506
rect 17066 24454 17078 24506
rect 17078 24454 17092 24506
rect 17116 24454 17130 24506
rect 17130 24454 17142 24506
rect 17142 24454 17172 24506
rect 17196 24454 17206 24506
rect 17206 24454 17252 24506
rect 16956 24452 17012 24454
rect 17036 24452 17092 24454
rect 17116 24452 17172 24454
rect 17196 24452 17252 24454
rect 16956 23418 17012 23420
rect 17036 23418 17092 23420
rect 17116 23418 17172 23420
rect 17196 23418 17252 23420
rect 16956 23366 17002 23418
rect 17002 23366 17012 23418
rect 17036 23366 17066 23418
rect 17066 23366 17078 23418
rect 17078 23366 17092 23418
rect 17116 23366 17130 23418
rect 17130 23366 17142 23418
rect 17142 23366 17172 23418
rect 17196 23366 17206 23418
rect 17206 23366 17252 23418
rect 16956 23364 17012 23366
rect 17036 23364 17092 23366
rect 17116 23364 17172 23366
rect 17196 23364 17252 23366
rect 16956 22330 17012 22332
rect 17036 22330 17092 22332
rect 17116 22330 17172 22332
rect 17196 22330 17252 22332
rect 16956 22278 17002 22330
rect 17002 22278 17012 22330
rect 17036 22278 17066 22330
rect 17066 22278 17078 22330
rect 17078 22278 17092 22330
rect 17116 22278 17130 22330
rect 17130 22278 17142 22330
rect 17142 22278 17172 22330
rect 17196 22278 17206 22330
rect 17206 22278 17252 22330
rect 16956 22276 17012 22278
rect 17036 22276 17092 22278
rect 17116 22276 17172 22278
rect 17196 22276 17252 22278
rect 16956 21242 17012 21244
rect 17036 21242 17092 21244
rect 17116 21242 17172 21244
rect 17196 21242 17252 21244
rect 16956 21190 17002 21242
rect 17002 21190 17012 21242
rect 17036 21190 17066 21242
rect 17066 21190 17078 21242
rect 17078 21190 17092 21242
rect 17116 21190 17130 21242
rect 17130 21190 17142 21242
rect 17142 21190 17172 21242
rect 17196 21190 17206 21242
rect 17206 21190 17252 21242
rect 16956 21188 17012 21190
rect 17036 21188 17092 21190
rect 17116 21188 17172 21190
rect 17196 21188 17252 21190
rect 16956 20154 17012 20156
rect 17036 20154 17092 20156
rect 17116 20154 17172 20156
rect 17196 20154 17252 20156
rect 16956 20102 17002 20154
rect 17002 20102 17012 20154
rect 17036 20102 17066 20154
rect 17066 20102 17078 20154
rect 17078 20102 17092 20154
rect 17116 20102 17130 20154
rect 17130 20102 17142 20154
rect 17142 20102 17172 20154
rect 17196 20102 17206 20154
rect 17206 20102 17252 20154
rect 16956 20100 17012 20102
rect 17036 20100 17092 20102
rect 17116 20100 17172 20102
rect 17196 20100 17252 20102
rect 16956 19066 17012 19068
rect 17036 19066 17092 19068
rect 17116 19066 17172 19068
rect 17196 19066 17252 19068
rect 16956 19014 17002 19066
rect 17002 19014 17012 19066
rect 17036 19014 17066 19066
rect 17066 19014 17078 19066
rect 17078 19014 17092 19066
rect 17116 19014 17130 19066
rect 17130 19014 17142 19066
rect 17142 19014 17172 19066
rect 17196 19014 17206 19066
rect 17206 19014 17252 19066
rect 16956 19012 17012 19014
rect 17036 19012 17092 19014
rect 17116 19012 17172 19014
rect 17196 19012 17252 19014
rect 17616 64218 17672 64220
rect 17696 64218 17752 64220
rect 17776 64218 17832 64220
rect 17856 64218 17912 64220
rect 17616 64166 17662 64218
rect 17662 64166 17672 64218
rect 17696 64166 17726 64218
rect 17726 64166 17738 64218
rect 17738 64166 17752 64218
rect 17776 64166 17790 64218
rect 17790 64166 17802 64218
rect 17802 64166 17832 64218
rect 17856 64166 17866 64218
rect 17866 64166 17912 64218
rect 17616 64164 17672 64166
rect 17696 64164 17752 64166
rect 17776 64164 17832 64166
rect 17856 64164 17912 64166
rect 17616 63130 17672 63132
rect 17696 63130 17752 63132
rect 17776 63130 17832 63132
rect 17856 63130 17912 63132
rect 17616 63078 17662 63130
rect 17662 63078 17672 63130
rect 17696 63078 17726 63130
rect 17726 63078 17738 63130
rect 17738 63078 17752 63130
rect 17776 63078 17790 63130
rect 17790 63078 17802 63130
rect 17802 63078 17832 63130
rect 17856 63078 17866 63130
rect 17866 63078 17912 63130
rect 17616 63076 17672 63078
rect 17696 63076 17752 63078
rect 17776 63076 17832 63078
rect 17856 63076 17912 63078
rect 17616 62042 17672 62044
rect 17696 62042 17752 62044
rect 17776 62042 17832 62044
rect 17856 62042 17912 62044
rect 17616 61990 17662 62042
rect 17662 61990 17672 62042
rect 17696 61990 17726 62042
rect 17726 61990 17738 62042
rect 17738 61990 17752 62042
rect 17776 61990 17790 62042
rect 17790 61990 17802 62042
rect 17802 61990 17832 62042
rect 17856 61990 17866 62042
rect 17866 61990 17912 62042
rect 17616 61988 17672 61990
rect 17696 61988 17752 61990
rect 17776 61988 17832 61990
rect 17856 61988 17912 61990
rect 17616 60954 17672 60956
rect 17696 60954 17752 60956
rect 17776 60954 17832 60956
rect 17856 60954 17912 60956
rect 17616 60902 17662 60954
rect 17662 60902 17672 60954
rect 17696 60902 17726 60954
rect 17726 60902 17738 60954
rect 17738 60902 17752 60954
rect 17776 60902 17790 60954
rect 17790 60902 17802 60954
rect 17802 60902 17832 60954
rect 17856 60902 17866 60954
rect 17866 60902 17912 60954
rect 17616 60900 17672 60902
rect 17696 60900 17752 60902
rect 17776 60900 17832 60902
rect 17856 60900 17912 60902
rect 17616 59866 17672 59868
rect 17696 59866 17752 59868
rect 17776 59866 17832 59868
rect 17856 59866 17912 59868
rect 17616 59814 17662 59866
rect 17662 59814 17672 59866
rect 17696 59814 17726 59866
rect 17726 59814 17738 59866
rect 17738 59814 17752 59866
rect 17776 59814 17790 59866
rect 17790 59814 17802 59866
rect 17802 59814 17832 59866
rect 17856 59814 17866 59866
rect 17866 59814 17912 59866
rect 17616 59812 17672 59814
rect 17696 59812 17752 59814
rect 17776 59812 17832 59814
rect 17856 59812 17912 59814
rect 17616 58778 17672 58780
rect 17696 58778 17752 58780
rect 17776 58778 17832 58780
rect 17856 58778 17912 58780
rect 17616 58726 17662 58778
rect 17662 58726 17672 58778
rect 17696 58726 17726 58778
rect 17726 58726 17738 58778
rect 17738 58726 17752 58778
rect 17776 58726 17790 58778
rect 17790 58726 17802 58778
rect 17802 58726 17832 58778
rect 17856 58726 17866 58778
rect 17866 58726 17912 58778
rect 17616 58724 17672 58726
rect 17696 58724 17752 58726
rect 17776 58724 17832 58726
rect 17856 58724 17912 58726
rect 17616 57690 17672 57692
rect 17696 57690 17752 57692
rect 17776 57690 17832 57692
rect 17856 57690 17912 57692
rect 17616 57638 17662 57690
rect 17662 57638 17672 57690
rect 17696 57638 17726 57690
rect 17726 57638 17738 57690
rect 17738 57638 17752 57690
rect 17776 57638 17790 57690
rect 17790 57638 17802 57690
rect 17802 57638 17832 57690
rect 17856 57638 17866 57690
rect 17866 57638 17912 57690
rect 17616 57636 17672 57638
rect 17696 57636 17752 57638
rect 17776 57636 17832 57638
rect 17856 57636 17912 57638
rect 17616 56602 17672 56604
rect 17696 56602 17752 56604
rect 17776 56602 17832 56604
rect 17856 56602 17912 56604
rect 17616 56550 17662 56602
rect 17662 56550 17672 56602
rect 17696 56550 17726 56602
rect 17726 56550 17738 56602
rect 17738 56550 17752 56602
rect 17776 56550 17790 56602
rect 17790 56550 17802 56602
rect 17802 56550 17832 56602
rect 17856 56550 17866 56602
rect 17866 56550 17912 56602
rect 17616 56548 17672 56550
rect 17696 56548 17752 56550
rect 17776 56548 17832 56550
rect 17856 56548 17912 56550
rect 17616 55514 17672 55516
rect 17696 55514 17752 55516
rect 17776 55514 17832 55516
rect 17856 55514 17912 55516
rect 17616 55462 17662 55514
rect 17662 55462 17672 55514
rect 17696 55462 17726 55514
rect 17726 55462 17738 55514
rect 17738 55462 17752 55514
rect 17776 55462 17790 55514
rect 17790 55462 17802 55514
rect 17802 55462 17832 55514
rect 17856 55462 17866 55514
rect 17866 55462 17912 55514
rect 17616 55460 17672 55462
rect 17696 55460 17752 55462
rect 17776 55460 17832 55462
rect 17856 55460 17912 55462
rect 17616 54426 17672 54428
rect 17696 54426 17752 54428
rect 17776 54426 17832 54428
rect 17856 54426 17912 54428
rect 17616 54374 17662 54426
rect 17662 54374 17672 54426
rect 17696 54374 17726 54426
rect 17726 54374 17738 54426
rect 17738 54374 17752 54426
rect 17776 54374 17790 54426
rect 17790 54374 17802 54426
rect 17802 54374 17832 54426
rect 17856 54374 17866 54426
rect 17866 54374 17912 54426
rect 17616 54372 17672 54374
rect 17696 54372 17752 54374
rect 17776 54372 17832 54374
rect 17856 54372 17912 54374
rect 17616 53338 17672 53340
rect 17696 53338 17752 53340
rect 17776 53338 17832 53340
rect 17856 53338 17912 53340
rect 17616 53286 17662 53338
rect 17662 53286 17672 53338
rect 17696 53286 17726 53338
rect 17726 53286 17738 53338
rect 17738 53286 17752 53338
rect 17776 53286 17790 53338
rect 17790 53286 17802 53338
rect 17802 53286 17832 53338
rect 17856 53286 17866 53338
rect 17866 53286 17912 53338
rect 17616 53284 17672 53286
rect 17696 53284 17752 53286
rect 17776 53284 17832 53286
rect 17856 53284 17912 53286
rect 17616 52250 17672 52252
rect 17696 52250 17752 52252
rect 17776 52250 17832 52252
rect 17856 52250 17912 52252
rect 17616 52198 17662 52250
rect 17662 52198 17672 52250
rect 17696 52198 17726 52250
rect 17726 52198 17738 52250
rect 17738 52198 17752 52250
rect 17776 52198 17790 52250
rect 17790 52198 17802 52250
rect 17802 52198 17832 52250
rect 17856 52198 17866 52250
rect 17866 52198 17912 52250
rect 17616 52196 17672 52198
rect 17696 52196 17752 52198
rect 17776 52196 17832 52198
rect 17856 52196 17912 52198
rect 17616 51162 17672 51164
rect 17696 51162 17752 51164
rect 17776 51162 17832 51164
rect 17856 51162 17912 51164
rect 17616 51110 17662 51162
rect 17662 51110 17672 51162
rect 17696 51110 17726 51162
rect 17726 51110 17738 51162
rect 17738 51110 17752 51162
rect 17776 51110 17790 51162
rect 17790 51110 17802 51162
rect 17802 51110 17832 51162
rect 17856 51110 17866 51162
rect 17866 51110 17912 51162
rect 17616 51108 17672 51110
rect 17696 51108 17752 51110
rect 17776 51108 17832 51110
rect 17856 51108 17912 51110
rect 17616 50074 17672 50076
rect 17696 50074 17752 50076
rect 17776 50074 17832 50076
rect 17856 50074 17912 50076
rect 17616 50022 17662 50074
rect 17662 50022 17672 50074
rect 17696 50022 17726 50074
rect 17726 50022 17738 50074
rect 17738 50022 17752 50074
rect 17776 50022 17790 50074
rect 17790 50022 17802 50074
rect 17802 50022 17832 50074
rect 17856 50022 17866 50074
rect 17866 50022 17912 50074
rect 17616 50020 17672 50022
rect 17696 50020 17752 50022
rect 17776 50020 17832 50022
rect 17856 50020 17912 50022
rect 17616 48986 17672 48988
rect 17696 48986 17752 48988
rect 17776 48986 17832 48988
rect 17856 48986 17912 48988
rect 17616 48934 17662 48986
rect 17662 48934 17672 48986
rect 17696 48934 17726 48986
rect 17726 48934 17738 48986
rect 17738 48934 17752 48986
rect 17776 48934 17790 48986
rect 17790 48934 17802 48986
rect 17802 48934 17832 48986
rect 17856 48934 17866 48986
rect 17866 48934 17912 48986
rect 17616 48932 17672 48934
rect 17696 48932 17752 48934
rect 17776 48932 17832 48934
rect 17856 48932 17912 48934
rect 17616 47898 17672 47900
rect 17696 47898 17752 47900
rect 17776 47898 17832 47900
rect 17856 47898 17912 47900
rect 17616 47846 17662 47898
rect 17662 47846 17672 47898
rect 17696 47846 17726 47898
rect 17726 47846 17738 47898
rect 17738 47846 17752 47898
rect 17776 47846 17790 47898
rect 17790 47846 17802 47898
rect 17802 47846 17832 47898
rect 17856 47846 17866 47898
rect 17866 47846 17912 47898
rect 17616 47844 17672 47846
rect 17696 47844 17752 47846
rect 17776 47844 17832 47846
rect 17856 47844 17912 47846
rect 17616 46810 17672 46812
rect 17696 46810 17752 46812
rect 17776 46810 17832 46812
rect 17856 46810 17912 46812
rect 17616 46758 17662 46810
rect 17662 46758 17672 46810
rect 17696 46758 17726 46810
rect 17726 46758 17738 46810
rect 17738 46758 17752 46810
rect 17776 46758 17790 46810
rect 17790 46758 17802 46810
rect 17802 46758 17832 46810
rect 17856 46758 17866 46810
rect 17866 46758 17912 46810
rect 17616 46756 17672 46758
rect 17696 46756 17752 46758
rect 17776 46756 17832 46758
rect 17856 46756 17912 46758
rect 17616 45722 17672 45724
rect 17696 45722 17752 45724
rect 17776 45722 17832 45724
rect 17856 45722 17912 45724
rect 17616 45670 17662 45722
rect 17662 45670 17672 45722
rect 17696 45670 17726 45722
rect 17726 45670 17738 45722
rect 17738 45670 17752 45722
rect 17776 45670 17790 45722
rect 17790 45670 17802 45722
rect 17802 45670 17832 45722
rect 17856 45670 17866 45722
rect 17866 45670 17912 45722
rect 17616 45668 17672 45670
rect 17696 45668 17752 45670
rect 17776 45668 17832 45670
rect 17856 45668 17912 45670
rect 17616 44634 17672 44636
rect 17696 44634 17752 44636
rect 17776 44634 17832 44636
rect 17856 44634 17912 44636
rect 17616 44582 17662 44634
rect 17662 44582 17672 44634
rect 17696 44582 17726 44634
rect 17726 44582 17738 44634
rect 17738 44582 17752 44634
rect 17776 44582 17790 44634
rect 17790 44582 17802 44634
rect 17802 44582 17832 44634
rect 17856 44582 17866 44634
rect 17866 44582 17912 44634
rect 17616 44580 17672 44582
rect 17696 44580 17752 44582
rect 17776 44580 17832 44582
rect 17856 44580 17912 44582
rect 17616 43546 17672 43548
rect 17696 43546 17752 43548
rect 17776 43546 17832 43548
rect 17856 43546 17912 43548
rect 17616 43494 17662 43546
rect 17662 43494 17672 43546
rect 17696 43494 17726 43546
rect 17726 43494 17738 43546
rect 17738 43494 17752 43546
rect 17776 43494 17790 43546
rect 17790 43494 17802 43546
rect 17802 43494 17832 43546
rect 17856 43494 17866 43546
rect 17866 43494 17912 43546
rect 17616 43492 17672 43494
rect 17696 43492 17752 43494
rect 17776 43492 17832 43494
rect 17856 43492 17912 43494
rect 17616 42458 17672 42460
rect 17696 42458 17752 42460
rect 17776 42458 17832 42460
rect 17856 42458 17912 42460
rect 17616 42406 17662 42458
rect 17662 42406 17672 42458
rect 17696 42406 17726 42458
rect 17726 42406 17738 42458
rect 17738 42406 17752 42458
rect 17776 42406 17790 42458
rect 17790 42406 17802 42458
rect 17802 42406 17832 42458
rect 17856 42406 17866 42458
rect 17866 42406 17912 42458
rect 17616 42404 17672 42406
rect 17696 42404 17752 42406
rect 17776 42404 17832 42406
rect 17856 42404 17912 42406
rect 17616 41370 17672 41372
rect 17696 41370 17752 41372
rect 17776 41370 17832 41372
rect 17856 41370 17912 41372
rect 17616 41318 17662 41370
rect 17662 41318 17672 41370
rect 17696 41318 17726 41370
rect 17726 41318 17738 41370
rect 17738 41318 17752 41370
rect 17776 41318 17790 41370
rect 17790 41318 17802 41370
rect 17802 41318 17832 41370
rect 17856 41318 17866 41370
rect 17866 41318 17912 41370
rect 17616 41316 17672 41318
rect 17696 41316 17752 41318
rect 17776 41316 17832 41318
rect 17856 41316 17912 41318
rect 17616 40282 17672 40284
rect 17696 40282 17752 40284
rect 17776 40282 17832 40284
rect 17856 40282 17912 40284
rect 17616 40230 17662 40282
rect 17662 40230 17672 40282
rect 17696 40230 17726 40282
rect 17726 40230 17738 40282
rect 17738 40230 17752 40282
rect 17776 40230 17790 40282
rect 17790 40230 17802 40282
rect 17802 40230 17832 40282
rect 17856 40230 17866 40282
rect 17866 40230 17912 40282
rect 17616 40228 17672 40230
rect 17696 40228 17752 40230
rect 17776 40228 17832 40230
rect 17856 40228 17912 40230
rect 17616 39194 17672 39196
rect 17696 39194 17752 39196
rect 17776 39194 17832 39196
rect 17856 39194 17912 39196
rect 17616 39142 17662 39194
rect 17662 39142 17672 39194
rect 17696 39142 17726 39194
rect 17726 39142 17738 39194
rect 17738 39142 17752 39194
rect 17776 39142 17790 39194
rect 17790 39142 17802 39194
rect 17802 39142 17832 39194
rect 17856 39142 17866 39194
rect 17866 39142 17912 39194
rect 17616 39140 17672 39142
rect 17696 39140 17752 39142
rect 17776 39140 17832 39142
rect 17856 39140 17912 39142
rect 17616 38106 17672 38108
rect 17696 38106 17752 38108
rect 17776 38106 17832 38108
rect 17856 38106 17912 38108
rect 17616 38054 17662 38106
rect 17662 38054 17672 38106
rect 17696 38054 17726 38106
rect 17726 38054 17738 38106
rect 17738 38054 17752 38106
rect 17776 38054 17790 38106
rect 17790 38054 17802 38106
rect 17802 38054 17832 38106
rect 17856 38054 17866 38106
rect 17866 38054 17912 38106
rect 17616 38052 17672 38054
rect 17696 38052 17752 38054
rect 17776 38052 17832 38054
rect 17856 38052 17912 38054
rect 17616 37018 17672 37020
rect 17696 37018 17752 37020
rect 17776 37018 17832 37020
rect 17856 37018 17912 37020
rect 17616 36966 17662 37018
rect 17662 36966 17672 37018
rect 17696 36966 17726 37018
rect 17726 36966 17738 37018
rect 17738 36966 17752 37018
rect 17776 36966 17790 37018
rect 17790 36966 17802 37018
rect 17802 36966 17832 37018
rect 17856 36966 17866 37018
rect 17866 36966 17912 37018
rect 17616 36964 17672 36966
rect 17696 36964 17752 36966
rect 17776 36964 17832 36966
rect 17856 36964 17912 36966
rect 17616 35930 17672 35932
rect 17696 35930 17752 35932
rect 17776 35930 17832 35932
rect 17856 35930 17912 35932
rect 17616 35878 17662 35930
rect 17662 35878 17672 35930
rect 17696 35878 17726 35930
rect 17726 35878 17738 35930
rect 17738 35878 17752 35930
rect 17776 35878 17790 35930
rect 17790 35878 17802 35930
rect 17802 35878 17832 35930
rect 17856 35878 17866 35930
rect 17866 35878 17912 35930
rect 17616 35876 17672 35878
rect 17696 35876 17752 35878
rect 17776 35876 17832 35878
rect 17856 35876 17912 35878
rect 17616 34842 17672 34844
rect 17696 34842 17752 34844
rect 17776 34842 17832 34844
rect 17856 34842 17912 34844
rect 17616 34790 17662 34842
rect 17662 34790 17672 34842
rect 17696 34790 17726 34842
rect 17726 34790 17738 34842
rect 17738 34790 17752 34842
rect 17776 34790 17790 34842
rect 17790 34790 17802 34842
rect 17802 34790 17832 34842
rect 17856 34790 17866 34842
rect 17866 34790 17912 34842
rect 17616 34788 17672 34790
rect 17696 34788 17752 34790
rect 17776 34788 17832 34790
rect 17856 34788 17912 34790
rect 17616 33754 17672 33756
rect 17696 33754 17752 33756
rect 17776 33754 17832 33756
rect 17856 33754 17912 33756
rect 17616 33702 17662 33754
rect 17662 33702 17672 33754
rect 17696 33702 17726 33754
rect 17726 33702 17738 33754
rect 17738 33702 17752 33754
rect 17776 33702 17790 33754
rect 17790 33702 17802 33754
rect 17802 33702 17832 33754
rect 17856 33702 17866 33754
rect 17866 33702 17912 33754
rect 17616 33700 17672 33702
rect 17696 33700 17752 33702
rect 17776 33700 17832 33702
rect 17856 33700 17912 33702
rect 17616 32666 17672 32668
rect 17696 32666 17752 32668
rect 17776 32666 17832 32668
rect 17856 32666 17912 32668
rect 17616 32614 17662 32666
rect 17662 32614 17672 32666
rect 17696 32614 17726 32666
rect 17726 32614 17738 32666
rect 17738 32614 17752 32666
rect 17776 32614 17790 32666
rect 17790 32614 17802 32666
rect 17802 32614 17832 32666
rect 17856 32614 17866 32666
rect 17866 32614 17912 32666
rect 17616 32612 17672 32614
rect 17696 32612 17752 32614
rect 17776 32612 17832 32614
rect 17856 32612 17912 32614
rect 17616 31578 17672 31580
rect 17696 31578 17752 31580
rect 17776 31578 17832 31580
rect 17856 31578 17912 31580
rect 17616 31526 17662 31578
rect 17662 31526 17672 31578
rect 17696 31526 17726 31578
rect 17726 31526 17738 31578
rect 17738 31526 17752 31578
rect 17776 31526 17790 31578
rect 17790 31526 17802 31578
rect 17802 31526 17832 31578
rect 17856 31526 17866 31578
rect 17866 31526 17912 31578
rect 17616 31524 17672 31526
rect 17696 31524 17752 31526
rect 17776 31524 17832 31526
rect 17856 31524 17912 31526
rect 17616 30490 17672 30492
rect 17696 30490 17752 30492
rect 17776 30490 17832 30492
rect 17856 30490 17912 30492
rect 17616 30438 17662 30490
rect 17662 30438 17672 30490
rect 17696 30438 17726 30490
rect 17726 30438 17738 30490
rect 17738 30438 17752 30490
rect 17776 30438 17790 30490
rect 17790 30438 17802 30490
rect 17802 30438 17832 30490
rect 17856 30438 17866 30490
rect 17866 30438 17912 30490
rect 17616 30436 17672 30438
rect 17696 30436 17752 30438
rect 17776 30436 17832 30438
rect 17856 30436 17912 30438
rect 17616 29402 17672 29404
rect 17696 29402 17752 29404
rect 17776 29402 17832 29404
rect 17856 29402 17912 29404
rect 17616 29350 17662 29402
rect 17662 29350 17672 29402
rect 17696 29350 17726 29402
rect 17726 29350 17738 29402
rect 17738 29350 17752 29402
rect 17776 29350 17790 29402
rect 17790 29350 17802 29402
rect 17802 29350 17832 29402
rect 17856 29350 17866 29402
rect 17866 29350 17912 29402
rect 17616 29348 17672 29350
rect 17696 29348 17752 29350
rect 17776 29348 17832 29350
rect 17856 29348 17912 29350
rect 17616 28314 17672 28316
rect 17696 28314 17752 28316
rect 17776 28314 17832 28316
rect 17856 28314 17912 28316
rect 17616 28262 17662 28314
rect 17662 28262 17672 28314
rect 17696 28262 17726 28314
rect 17726 28262 17738 28314
rect 17738 28262 17752 28314
rect 17776 28262 17790 28314
rect 17790 28262 17802 28314
rect 17802 28262 17832 28314
rect 17856 28262 17866 28314
rect 17866 28262 17912 28314
rect 17616 28260 17672 28262
rect 17696 28260 17752 28262
rect 17776 28260 17832 28262
rect 17856 28260 17912 28262
rect 17616 27226 17672 27228
rect 17696 27226 17752 27228
rect 17776 27226 17832 27228
rect 17856 27226 17912 27228
rect 17616 27174 17662 27226
rect 17662 27174 17672 27226
rect 17696 27174 17726 27226
rect 17726 27174 17738 27226
rect 17738 27174 17752 27226
rect 17776 27174 17790 27226
rect 17790 27174 17802 27226
rect 17802 27174 17832 27226
rect 17856 27174 17866 27226
rect 17866 27174 17912 27226
rect 17616 27172 17672 27174
rect 17696 27172 17752 27174
rect 17776 27172 17832 27174
rect 17856 27172 17912 27174
rect 17616 26138 17672 26140
rect 17696 26138 17752 26140
rect 17776 26138 17832 26140
rect 17856 26138 17912 26140
rect 17616 26086 17662 26138
rect 17662 26086 17672 26138
rect 17696 26086 17726 26138
rect 17726 26086 17738 26138
rect 17738 26086 17752 26138
rect 17776 26086 17790 26138
rect 17790 26086 17802 26138
rect 17802 26086 17832 26138
rect 17856 26086 17866 26138
rect 17866 26086 17912 26138
rect 17616 26084 17672 26086
rect 17696 26084 17752 26086
rect 17776 26084 17832 26086
rect 17856 26084 17912 26086
rect 17616 25050 17672 25052
rect 17696 25050 17752 25052
rect 17776 25050 17832 25052
rect 17856 25050 17912 25052
rect 17616 24998 17662 25050
rect 17662 24998 17672 25050
rect 17696 24998 17726 25050
rect 17726 24998 17738 25050
rect 17738 24998 17752 25050
rect 17776 24998 17790 25050
rect 17790 24998 17802 25050
rect 17802 24998 17832 25050
rect 17856 24998 17866 25050
rect 17866 24998 17912 25050
rect 17616 24996 17672 24998
rect 17696 24996 17752 24998
rect 17776 24996 17832 24998
rect 17856 24996 17912 24998
rect 17616 23962 17672 23964
rect 17696 23962 17752 23964
rect 17776 23962 17832 23964
rect 17856 23962 17912 23964
rect 17616 23910 17662 23962
rect 17662 23910 17672 23962
rect 17696 23910 17726 23962
rect 17726 23910 17738 23962
rect 17738 23910 17752 23962
rect 17776 23910 17790 23962
rect 17790 23910 17802 23962
rect 17802 23910 17832 23962
rect 17856 23910 17866 23962
rect 17866 23910 17912 23962
rect 17616 23908 17672 23910
rect 17696 23908 17752 23910
rect 17776 23908 17832 23910
rect 17856 23908 17912 23910
rect 17616 22874 17672 22876
rect 17696 22874 17752 22876
rect 17776 22874 17832 22876
rect 17856 22874 17912 22876
rect 17616 22822 17662 22874
rect 17662 22822 17672 22874
rect 17696 22822 17726 22874
rect 17726 22822 17738 22874
rect 17738 22822 17752 22874
rect 17776 22822 17790 22874
rect 17790 22822 17802 22874
rect 17802 22822 17832 22874
rect 17856 22822 17866 22874
rect 17866 22822 17912 22874
rect 17616 22820 17672 22822
rect 17696 22820 17752 22822
rect 17776 22820 17832 22822
rect 17856 22820 17912 22822
rect 17616 21786 17672 21788
rect 17696 21786 17752 21788
rect 17776 21786 17832 21788
rect 17856 21786 17912 21788
rect 17616 21734 17662 21786
rect 17662 21734 17672 21786
rect 17696 21734 17726 21786
rect 17726 21734 17738 21786
rect 17738 21734 17752 21786
rect 17776 21734 17790 21786
rect 17790 21734 17802 21786
rect 17802 21734 17832 21786
rect 17856 21734 17866 21786
rect 17866 21734 17912 21786
rect 17616 21732 17672 21734
rect 17696 21732 17752 21734
rect 17776 21732 17832 21734
rect 17856 21732 17912 21734
rect 17616 20698 17672 20700
rect 17696 20698 17752 20700
rect 17776 20698 17832 20700
rect 17856 20698 17912 20700
rect 17616 20646 17662 20698
rect 17662 20646 17672 20698
rect 17696 20646 17726 20698
rect 17726 20646 17738 20698
rect 17738 20646 17752 20698
rect 17776 20646 17790 20698
rect 17790 20646 17802 20698
rect 17802 20646 17832 20698
rect 17856 20646 17866 20698
rect 17866 20646 17912 20698
rect 17616 20644 17672 20646
rect 17696 20644 17752 20646
rect 17776 20644 17832 20646
rect 17856 20644 17912 20646
rect 17616 19610 17672 19612
rect 17696 19610 17752 19612
rect 17776 19610 17832 19612
rect 17856 19610 17912 19612
rect 17616 19558 17662 19610
rect 17662 19558 17672 19610
rect 17696 19558 17726 19610
rect 17726 19558 17738 19610
rect 17738 19558 17752 19610
rect 17776 19558 17790 19610
rect 17790 19558 17802 19610
rect 17802 19558 17832 19610
rect 17856 19558 17866 19610
rect 17866 19558 17912 19610
rect 17616 19556 17672 19558
rect 17696 19556 17752 19558
rect 17776 19556 17832 19558
rect 17856 19556 17912 19558
rect 17616 18522 17672 18524
rect 17696 18522 17752 18524
rect 17776 18522 17832 18524
rect 17856 18522 17912 18524
rect 17616 18470 17662 18522
rect 17662 18470 17672 18522
rect 17696 18470 17726 18522
rect 17726 18470 17738 18522
rect 17738 18470 17752 18522
rect 17776 18470 17790 18522
rect 17790 18470 17802 18522
rect 17802 18470 17832 18522
rect 17856 18470 17866 18522
rect 17866 18470 17912 18522
rect 17616 18468 17672 18470
rect 17696 18468 17752 18470
rect 17776 18468 17832 18470
rect 17856 18468 17912 18470
rect 16956 17978 17012 17980
rect 17036 17978 17092 17980
rect 17116 17978 17172 17980
rect 17196 17978 17252 17980
rect 16956 17926 17002 17978
rect 17002 17926 17012 17978
rect 17036 17926 17066 17978
rect 17066 17926 17078 17978
rect 17078 17926 17092 17978
rect 17116 17926 17130 17978
rect 17130 17926 17142 17978
rect 17142 17926 17172 17978
rect 17196 17926 17206 17978
rect 17206 17926 17252 17978
rect 16956 17924 17012 17926
rect 17036 17924 17092 17926
rect 17116 17924 17172 17926
rect 17196 17924 17252 17926
rect 17616 17434 17672 17436
rect 17696 17434 17752 17436
rect 17776 17434 17832 17436
rect 17856 17434 17912 17436
rect 17616 17382 17662 17434
rect 17662 17382 17672 17434
rect 17696 17382 17726 17434
rect 17726 17382 17738 17434
rect 17738 17382 17752 17434
rect 17776 17382 17790 17434
rect 17790 17382 17802 17434
rect 17802 17382 17832 17434
rect 17856 17382 17866 17434
rect 17866 17382 17912 17434
rect 17616 17380 17672 17382
rect 17696 17380 17752 17382
rect 17776 17380 17832 17382
rect 17856 17380 17912 17382
rect 16956 16890 17012 16892
rect 17036 16890 17092 16892
rect 17116 16890 17172 16892
rect 17196 16890 17252 16892
rect 16956 16838 17002 16890
rect 17002 16838 17012 16890
rect 17036 16838 17066 16890
rect 17066 16838 17078 16890
rect 17078 16838 17092 16890
rect 17116 16838 17130 16890
rect 17130 16838 17142 16890
rect 17142 16838 17172 16890
rect 17196 16838 17206 16890
rect 17206 16838 17252 16890
rect 16956 16836 17012 16838
rect 17036 16836 17092 16838
rect 17116 16836 17172 16838
rect 17196 16836 17252 16838
rect 16956 15802 17012 15804
rect 17036 15802 17092 15804
rect 17116 15802 17172 15804
rect 17196 15802 17252 15804
rect 16956 15750 17002 15802
rect 17002 15750 17012 15802
rect 17036 15750 17066 15802
rect 17066 15750 17078 15802
rect 17078 15750 17092 15802
rect 17116 15750 17130 15802
rect 17130 15750 17142 15802
rect 17142 15750 17172 15802
rect 17196 15750 17206 15802
rect 17206 15750 17252 15802
rect 16956 15748 17012 15750
rect 17036 15748 17092 15750
rect 17116 15748 17172 15750
rect 17196 15748 17252 15750
rect 16956 14714 17012 14716
rect 17036 14714 17092 14716
rect 17116 14714 17172 14716
rect 17196 14714 17252 14716
rect 16956 14662 17002 14714
rect 17002 14662 17012 14714
rect 17036 14662 17066 14714
rect 17066 14662 17078 14714
rect 17078 14662 17092 14714
rect 17116 14662 17130 14714
rect 17130 14662 17142 14714
rect 17142 14662 17172 14714
rect 17196 14662 17206 14714
rect 17206 14662 17252 14714
rect 16956 14660 17012 14662
rect 17036 14660 17092 14662
rect 17116 14660 17172 14662
rect 17196 14660 17252 14662
rect 16956 13626 17012 13628
rect 17036 13626 17092 13628
rect 17116 13626 17172 13628
rect 17196 13626 17252 13628
rect 16956 13574 17002 13626
rect 17002 13574 17012 13626
rect 17036 13574 17066 13626
rect 17066 13574 17078 13626
rect 17078 13574 17092 13626
rect 17116 13574 17130 13626
rect 17130 13574 17142 13626
rect 17142 13574 17172 13626
rect 17196 13574 17206 13626
rect 17206 13574 17252 13626
rect 16956 13572 17012 13574
rect 17036 13572 17092 13574
rect 17116 13572 17172 13574
rect 17196 13572 17252 13574
rect 16956 12538 17012 12540
rect 17036 12538 17092 12540
rect 17116 12538 17172 12540
rect 17196 12538 17252 12540
rect 16956 12486 17002 12538
rect 17002 12486 17012 12538
rect 17036 12486 17066 12538
rect 17066 12486 17078 12538
rect 17078 12486 17092 12538
rect 17116 12486 17130 12538
rect 17130 12486 17142 12538
rect 17142 12486 17172 12538
rect 17196 12486 17206 12538
rect 17206 12486 17252 12538
rect 16956 12484 17012 12486
rect 17036 12484 17092 12486
rect 17116 12484 17172 12486
rect 17196 12484 17252 12486
rect 16956 11450 17012 11452
rect 17036 11450 17092 11452
rect 17116 11450 17172 11452
rect 17196 11450 17252 11452
rect 16956 11398 17002 11450
rect 17002 11398 17012 11450
rect 17036 11398 17066 11450
rect 17066 11398 17078 11450
rect 17078 11398 17092 11450
rect 17116 11398 17130 11450
rect 17130 11398 17142 11450
rect 17142 11398 17172 11450
rect 17196 11398 17206 11450
rect 17206 11398 17252 11450
rect 16956 11396 17012 11398
rect 17036 11396 17092 11398
rect 17116 11396 17172 11398
rect 17196 11396 17252 11398
rect 16956 10362 17012 10364
rect 17036 10362 17092 10364
rect 17116 10362 17172 10364
rect 17196 10362 17252 10364
rect 16956 10310 17002 10362
rect 17002 10310 17012 10362
rect 17036 10310 17066 10362
rect 17066 10310 17078 10362
rect 17078 10310 17092 10362
rect 17116 10310 17130 10362
rect 17130 10310 17142 10362
rect 17142 10310 17172 10362
rect 17196 10310 17206 10362
rect 17206 10310 17252 10362
rect 16956 10308 17012 10310
rect 17036 10308 17092 10310
rect 17116 10308 17172 10310
rect 17196 10308 17252 10310
rect 17616 16346 17672 16348
rect 17696 16346 17752 16348
rect 17776 16346 17832 16348
rect 17856 16346 17912 16348
rect 17616 16294 17662 16346
rect 17662 16294 17672 16346
rect 17696 16294 17726 16346
rect 17726 16294 17738 16346
rect 17738 16294 17752 16346
rect 17776 16294 17790 16346
rect 17790 16294 17802 16346
rect 17802 16294 17832 16346
rect 17856 16294 17866 16346
rect 17866 16294 17912 16346
rect 17616 16292 17672 16294
rect 17696 16292 17752 16294
rect 17776 16292 17832 16294
rect 17856 16292 17912 16294
rect 17616 15258 17672 15260
rect 17696 15258 17752 15260
rect 17776 15258 17832 15260
rect 17856 15258 17912 15260
rect 17616 15206 17662 15258
rect 17662 15206 17672 15258
rect 17696 15206 17726 15258
rect 17726 15206 17738 15258
rect 17738 15206 17752 15258
rect 17776 15206 17790 15258
rect 17790 15206 17802 15258
rect 17802 15206 17832 15258
rect 17856 15206 17866 15258
rect 17866 15206 17912 15258
rect 17616 15204 17672 15206
rect 17696 15204 17752 15206
rect 17776 15204 17832 15206
rect 17856 15204 17912 15206
rect 17616 14170 17672 14172
rect 17696 14170 17752 14172
rect 17776 14170 17832 14172
rect 17856 14170 17912 14172
rect 17616 14118 17662 14170
rect 17662 14118 17672 14170
rect 17696 14118 17726 14170
rect 17726 14118 17738 14170
rect 17738 14118 17752 14170
rect 17776 14118 17790 14170
rect 17790 14118 17802 14170
rect 17802 14118 17832 14170
rect 17856 14118 17866 14170
rect 17866 14118 17912 14170
rect 17616 14116 17672 14118
rect 17696 14116 17752 14118
rect 17776 14116 17832 14118
rect 17856 14116 17912 14118
rect 17616 13082 17672 13084
rect 17696 13082 17752 13084
rect 17776 13082 17832 13084
rect 17856 13082 17912 13084
rect 17616 13030 17662 13082
rect 17662 13030 17672 13082
rect 17696 13030 17726 13082
rect 17726 13030 17738 13082
rect 17738 13030 17752 13082
rect 17776 13030 17790 13082
rect 17790 13030 17802 13082
rect 17802 13030 17832 13082
rect 17856 13030 17866 13082
rect 17866 13030 17912 13082
rect 17616 13028 17672 13030
rect 17696 13028 17752 13030
rect 17776 13028 17832 13030
rect 17856 13028 17912 13030
rect 19614 34448 19670 34504
rect 17616 11994 17672 11996
rect 17696 11994 17752 11996
rect 17776 11994 17832 11996
rect 17856 11994 17912 11996
rect 17616 11942 17662 11994
rect 17662 11942 17672 11994
rect 17696 11942 17726 11994
rect 17726 11942 17738 11994
rect 17738 11942 17752 11994
rect 17776 11942 17790 11994
rect 17790 11942 17802 11994
rect 17802 11942 17832 11994
rect 17856 11942 17866 11994
rect 17866 11942 17912 11994
rect 17616 11940 17672 11942
rect 17696 11940 17752 11942
rect 17776 11940 17832 11942
rect 17856 11940 17912 11942
rect 17616 10906 17672 10908
rect 17696 10906 17752 10908
rect 17776 10906 17832 10908
rect 17856 10906 17912 10908
rect 17616 10854 17662 10906
rect 17662 10854 17672 10906
rect 17696 10854 17726 10906
rect 17726 10854 17738 10906
rect 17738 10854 17752 10906
rect 17776 10854 17790 10906
rect 17790 10854 17802 10906
rect 17802 10854 17832 10906
rect 17856 10854 17866 10906
rect 17866 10854 17912 10906
rect 17616 10852 17672 10854
rect 17696 10852 17752 10854
rect 17776 10852 17832 10854
rect 17856 10852 17912 10854
rect 17616 9818 17672 9820
rect 17696 9818 17752 9820
rect 17776 9818 17832 9820
rect 17856 9818 17912 9820
rect 17616 9766 17662 9818
rect 17662 9766 17672 9818
rect 17696 9766 17726 9818
rect 17726 9766 17738 9818
rect 17738 9766 17752 9818
rect 17776 9766 17790 9818
rect 17790 9766 17802 9818
rect 17802 9766 17832 9818
rect 17856 9766 17866 9818
rect 17866 9766 17912 9818
rect 17616 9764 17672 9766
rect 17696 9764 17752 9766
rect 17776 9764 17832 9766
rect 17856 9764 17912 9766
rect 16956 9274 17012 9276
rect 17036 9274 17092 9276
rect 17116 9274 17172 9276
rect 17196 9274 17252 9276
rect 16956 9222 17002 9274
rect 17002 9222 17012 9274
rect 17036 9222 17066 9274
rect 17066 9222 17078 9274
rect 17078 9222 17092 9274
rect 17116 9222 17130 9274
rect 17130 9222 17142 9274
rect 17142 9222 17172 9274
rect 17196 9222 17206 9274
rect 17206 9222 17252 9274
rect 16956 9220 17012 9222
rect 17036 9220 17092 9222
rect 17116 9220 17172 9222
rect 17196 9220 17252 9222
rect 17616 8730 17672 8732
rect 17696 8730 17752 8732
rect 17776 8730 17832 8732
rect 17856 8730 17912 8732
rect 17616 8678 17662 8730
rect 17662 8678 17672 8730
rect 17696 8678 17726 8730
rect 17726 8678 17738 8730
rect 17738 8678 17752 8730
rect 17776 8678 17790 8730
rect 17790 8678 17802 8730
rect 17802 8678 17832 8730
rect 17856 8678 17866 8730
rect 17866 8678 17912 8730
rect 17616 8676 17672 8678
rect 17696 8676 17752 8678
rect 17776 8676 17832 8678
rect 17856 8676 17912 8678
rect 16956 8186 17012 8188
rect 17036 8186 17092 8188
rect 17116 8186 17172 8188
rect 17196 8186 17252 8188
rect 16956 8134 17002 8186
rect 17002 8134 17012 8186
rect 17036 8134 17066 8186
rect 17066 8134 17078 8186
rect 17078 8134 17092 8186
rect 17116 8134 17130 8186
rect 17130 8134 17142 8186
rect 17142 8134 17172 8186
rect 17196 8134 17206 8186
rect 17206 8134 17252 8186
rect 16956 8132 17012 8134
rect 17036 8132 17092 8134
rect 17116 8132 17172 8134
rect 17196 8132 17252 8134
rect 17616 7642 17672 7644
rect 17696 7642 17752 7644
rect 17776 7642 17832 7644
rect 17856 7642 17912 7644
rect 17616 7590 17662 7642
rect 17662 7590 17672 7642
rect 17696 7590 17726 7642
rect 17726 7590 17738 7642
rect 17738 7590 17752 7642
rect 17776 7590 17790 7642
rect 17790 7590 17802 7642
rect 17802 7590 17832 7642
rect 17856 7590 17866 7642
rect 17866 7590 17912 7642
rect 17616 7588 17672 7590
rect 17696 7588 17752 7590
rect 17776 7588 17832 7590
rect 17856 7588 17912 7590
rect 16956 7098 17012 7100
rect 17036 7098 17092 7100
rect 17116 7098 17172 7100
rect 17196 7098 17252 7100
rect 16956 7046 17002 7098
rect 17002 7046 17012 7098
rect 17036 7046 17066 7098
rect 17066 7046 17078 7098
rect 17078 7046 17092 7098
rect 17116 7046 17130 7098
rect 17130 7046 17142 7098
rect 17142 7046 17172 7098
rect 17196 7046 17206 7098
rect 17206 7046 17252 7098
rect 16956 7044 17012 7046
rect 17036 7044 17092 7046
rect 17116 7044 17172 7046
rect 17196 7044 17252 7046
rect 17616 6554 17672 6556
rect 17696 6554 17752 6556
rect 17776 6554 17832 6556
rect 17856 6554 17912 6556
rect 17616 6502 17662 6554
rect 17662 6502 17672 6554
rect 17696 6502 17726 6554
rect 17726 6502 17738 6554
rect 17738 6502 17752 6554
rect 17776 6502 17790 6554
rect 17790 6502 17802 6554
rect 17802 6502 17832 6554
rect 17856 6502 17866 6554
rect 17866 6502 17912 6554
rect 17616 6500 17672 6502
rect 17696 6500 17752 6502
rect 17776 6500 17832 6502
rect 17856 6500 17912 6502
rect 16956 6010 17012 6012
rect 17036 6010 17092 6012
rect 17116 6010 17172 6012
rect 17196 6010 17252 6012
rect 16956 5958 17002 6010
rect 17002 5958 17012 6010
rect 17036 5958 17066 6010
rect 17066 5958 17078 6010
rect 17078 5958 17092 6010
rect 17116 5958 17130 6010
rect 17130 5958 17142 6010
rect 17142 5958 17172 6010
rect 17196 5958 17206 6010
rect 17206 5958 17252 6010
rect 16956 5956 17012 5958
rect 17036 5956 17092 5958
rect 17116 5956 17172 5958
rect 17196 5956 17252 5958
rect 17616 5466 17672 5468
rect 17696 5466 17752 5468
rect 17776 5466 17832 5468
rect 17856 5466 17912 5468
rect 17616 5414 17662 5466
rect 17662 5414 17672 5466
rect 17696 5414 17726 5466
rect 17726 5414 17738 5466
rect 17738 5414 17752 5466
rect 17776 5414 17790 5466
rect 17790 5414 17802 5466
rect 17802 5414 17832 5466
rect 17856 5414 17866 5466
rect 17866 5414 17912 5466
rect 17616 5412 17672 5414
rect 17696 5412 17752 5414
rect 17776 5412 17832 5414
rect 17856 5412 17912 5414
rect 16956 4922 17012 4924
rect 17036 4922 17092 4924
rect 17116 4922 17172 4924
rect 17196 4922 17252 4924
rect 16956 4870 17002 4922
rect 17002 4870 17012 4922
rect 17036 4870 17066 4922
rect 17066 4870 17078 4922
rect 17078 4870 17092 4922
rect 17116 4870 17130 4922
rect 17130 4870 17142 4922
rect 17142 4870 17172 4922
rect 17196 4870 17206 4922
rect 17206 4870 17252 4922
rect 16956 4868 17012 4870
rect 17036 4868 17092 4870
rect 17116 4868 17172 4870
rect 17196 4868 17252 4870
rect 17616 4378 17672 4380
rect 17696 4378 17752 4380
rect 17776 4378 17832 4380
rect 17856 4378 17912 4380
rect 17616 4326 17662 4378
rect 17662 4326 17672 4378
rect 17696 4326 17726 4378
rect 17726 4326 17738 4378
rect 17738 4326 17752 4378
rect 17776 4326 17790 4378
rect 17790 4326 17802 4378
rect 17802 4326 17832 4378
rect 17856 4326 17866 4378
rect 17866 4326 17912 4378
rect 17616 4324 17672 4326
rect 17696 4324 17752 4326
rect 17776 4324 17832 4326
rect 17856 4324 17912 4326
rect 16956 3834 17012 3836
rect 17036 3834 17092 3836
rect 17116 3834 17172 3836
rect 17196 3834 17252 3836
rect 16956 3782 17002 3834
rect 17002 3782 17012 3834
rect 17036 3782 17066 3834
rect 17066 3782 17078 3834
rect 17078 3782 17092 3834
rect 17116 3782 17130 3834
rect 17130 3782 17142 3834
rect 17142 3782 17172 3834
rect 17196 3782 17206 3834
rect 17206 3782 17252 3834
rect 16956 3780 17012 3782
rect 17036 3780 17092 3782
rect 17116 3780 17172 3782
rect 17196 3780 17252 3782
rect 17616 3290 17672 3292
rect 17696 3290 17752 3292
rect 17776 3290 17832 3292
rect 17856 3290 17912 3292
rect 17616 3238 17662 3290
rect 17662 3238 17672 3290
rect 17696 3238 17726 3290
rect 17726 3238 17738 3290
rect 17738 3238 17752 3290
rect 17776 3238 17790 3290
rect 17790 3238 17802 3290
rect 17802 3238 17832 3290
rect 17856 3238 17866 3290
rect 17866 3238 17912 3290
rect 17616 3236 17672 3238
rect 17696 3236 17752 3238
rect 17776 3236 17832 3238
rect 17856 3236 17912 3238
rect 16956 2746 17012 2748
rect 17036 2746 17092 2748
rect 17116 2746 17172 2748
rect 17196 2746 17252 2748
rect 16956 2694 17002 2746
rect 17002 2694 17012 2746
rect 17036 2694 17066 2746
rect 17066 2694 17078 2746
rect 17078 2694 17092 2746
rect 17116 2694 17130 2746
rect 17130 2694 17142 2746
rect 17142 2694 17172 2746
rect 17196 2694 17206 2746
rect 17206 2694 17252 2746
rect 16956 2692 17012 2694
rect 17036 2692 17092 2694
rect 17116 2692 17172 2694
rect 17196 2692 17252 2694
rect 21086 33804 21088 33824
rect 21088 33804 21140 33824
rect 21140 33804 21142 33824
rect 21086 33768 21142 33804
rect 21956 69114 22012 69116
rect 22036 69114 22092 69116
rect 22116 69114 22172 69116
rect 22196 69114 22252 69116
rect 21956 69062 22002 69114
rect 22002 69062 22012 69114
rect 22036 69062 22066 69114
rect 22066 69062 22078 69114
rect 22078 69062 22092 69114
rect 22116 69062 22130 69114
rect 22130 69062 22142 69114
rect 22142 69062 22172 69114
rect 22196 69062 22206 69114
rect 22206 69062 22252 69114
rect 21956 69060 22012 69062
rect 22036 69060 22092 69062
rect 22116 69060 22172 69062
rect 22196 69060 22252 69062
rect 26956 69114 27012 69116
rect 27036 69114 27092 69116
rect 27116 69114 27172 69116
rect 27196 69114 27252 69116
rect 26956 69062 27002 69114
rect 27002 69062 27012 69114
rect 27036 69062 27066 69114
rect 27066 69062 27078 69114
rect 27078 69062 27092 69114
rect 27116 69062 27130 69114
rect 27130 69062 27142 69114
rect 27142 69062 27172 69114
rect 27196 69062 27206 69114
rect 27206 69062 27252 69114
rect 26956 69060 27012 69062
rect 27036 69060 27092 69062
rect 27116 69060 27172 69062
rect 27196 69060 27252 69062
rect 22616 68570 22672 68572
rect 22696 68570 22752 68572
rect 22776 68570 22832 68572
rect 22856 68570 22912 68572
rect 22616 68518 22662 68570
rect 22662 68518 22672 68570
rect 22696 68518 22726 68570
rect 22726 68518 22738 68570
rect 22738 68518 22752 68570
rect 22776 68518 22790 68570
rect 22790 68518 22802 68570
rect 22802 68518 22832 68570
rect 22856 68518 22866 68570
rect 22866 68518 22912 68570
rect 22616 68516 22672 68518
rect 22696 68516 22752 68518
rect 22776 68516 22832 68518
rect 22856 68516 22912 68518
rect 21956 68026 22012 68028
rect 22036 68026 22092 68028
rect 22116 68026 22172 68028
rect 22196 68026 22252 68028
rect 21956 67974 22002 68026
rect 22002 67974 22012 68026
rect 22036 67974 22066 68026
rect 22066 67974 22078 68026
rect 22078 67974 22092 68026
rect 22116 67974 22130 68026
rect 22130 67974 22142 68026
rect 22142 67974 22172 68026
rect 22196 67974 22206 68026
rect 22206 67974 22252 68026
rect 21956 67972 22012 67974
rect 22036 67972 22092 67974
rect 22116 67972 22172 67974
rect 22196 67972 22252 67974
rect 26956 68026 27012 68028
rect 27036 68026 27092 68028
rect 27116 68026 27172 68028
rect 27196 68026 27252 68028
rect 26956 67974 27002 68026
rect 27002 67974 27012 68026
rect 27036 67974 27066 68026
rect 27066 67974 27078 68026
rect 27078 67974 27092 68026
rect 27116 67974 27130 68026
rect 27130 67974 27142 68026
rect 27142 67974 27172 68026
rect 27196 67974 27206 68026
rect 27206 67974 27252 68026
rect 26956 67972 27012 67974
rect 27036 67972 27092 67974
rect 27116 67972 27172 67974
rect 27196 67972 27252 67974
rect 22616 67482 22672 67484
rect 22696 67482 22752 67484
rect 22776 67482 22832 67484
rect 22856 67482 22912 67484
rect 22616 67430 22662 67482
rect 22662 67430 22672 67482
rect 22696 67430 22726 67482
rect 22726 67430 22738 67482
rect 22738 67430 22752 67482
rect 22776 67430 22790 67482
rect 22790 67430 22802 67482
rect 22802 67430 22832 67482
rect 22856 67430 22866 67482
rect 22866 67430 22912 67482
rect 22616 67428 22672 67430
rect 22696 67428 22752 67430
rect 22776 67428 22832 67430
rect 22856 67428 22912 67430
rect 21956 66938 22012 66940
rect 22036 66938 22092 66940
rect 22116 66938 22172 66940
rect 22196 66938 22252 66940
rect 21956 66886 22002 66938
rect 22002 66886 22012 66938
rect 22036 66886 22066 66938
rect 22066 66886 22078 66938
rect 22078 66886 22092 66938
rect 22116 66886 22130 66938
rect 22130 66886 22142 66938
rect 22142 66886 22172 66938
rect 22196 66886 22206 66938
rect 22206 66886 22252 66938
rect 21956 66884 22012 66886
rect 22036 66884 22092 66886
rect 22116 66884 22172 66886
rect 22196 66884 22252 66886
rect 22616 66394 22672 66396
rect 22696 66394 22752 66396
rect 22776 66394 22832 66396
rect 22856 66394 22912 66396
rect 22616 66342 22662 66394
rect 22662 66342 22672 66394
rect 22696 66342 22726 66394
rect 22726 66342 22738 66394
rect 22738 66342 22752 66394
rect 22776 66342 22790 66394
rect 22790 66342 22802 66394
rect 22802 66342 22832 66394
rect 22856 66342 22866 66394
rect 22866 66342 22912 66394
rect 22616 66340 22672 66342
rect 22696 66340 22752 66342
rect 22776 66340 22832 66342
rect 22856 66340 22912 66342
rect 21956 65850 22012 65852
rect 22036 65850 22092 65852
rect 22116 65850 22172 65852
rect 22196 65850 22252 65852
rect 21956 65798 22002 65850
rect 22002 65798 22012 65850
rect 22036 65798 22066 65850
rect 22066 65798 22078 65850
rect 22078 65798 22092 65850
rect 22116 65798 22130 65850
rect 22130 65798 22142 65850
rect 22142 65798 22172 65850
rect 22196 65798 22206 65850
rect 22206 65798 22252 65850
rect 21956 65796 22012 65798
rect 22036 65796 22092 65798
rect 22116 65796 22172 65798
rect 22196 65796 22252 65798
rect 22616 65306 22672 65308
rect 22696 65306 22752 65308
rect 22776 65306 22832 65308
rect 22856 65306 22912 65308
rect 22616 65254 22662 65306
rect 22662 65254 22672 65306
rect 22696 65254 22726 65306
rect 22726 65254 22738 65306
rect 22738 65254 22752 65306
rect 22776 65254 22790 65306
rect 22790 65254 22802 65306
rect 22802 65254 22832 65306
rect 22856 65254 22866 65306
rect 22866 65254 22912 65306
rect 22616 65252 22672 65254
rect 22696 65252 22752 65254
rect 22776 65252 22832 65254
rect 22856 65252 22912 65254
rect 21956 64762 22012 64764
rect 22036 64762 22092 64764
rect 22116 64762 22172 64764
rect 22196 64762 22252 64764
rect 21956 64710 22002 64762
rect 22002 64710 22012 64762
rect 22036 64710 22066 64762
rect 22066 64710 22078 64762
rect 22078 64710 22092 64762
rect 22116 64710 22130 64762
rect 22130 64710 22142 64762
rect 22142 64710 22172 64762
rect 22196 64710 22206 64762
rect 22206 64710 22252 64762
rect 21956 64708 22012 64710
rect 22036 64708 22092 64710
rect 22116 64708 22172 64710
rect 22196 64708 22252 64710
rect 21956 63674 22012 63676
rect 22036 63674 22092 63676
rect 22116 63674 22172 63676
rect 22196 63674 22252 63676
rect 21956 63622 22002 63674
rect 22002 63622 22012 63674
rect 22036 63622 22066 63674
rect 22066 63622 22078 63674
rect 22078 63622 22092 63674
rect 22116 63622 22130 63674
rect 22130 63622 22142 63674
rect 22142 63622 22172 63674
rect 22196 63622 22206 63674
rect 22206 63622 22252 63674
rect 21956 63620 22012 63622
rect 22036 63620 22092 63622
rect 22116 63620 22172 63622
rect 22196 63620 22252 63622
rect 21956 62586 22012 62588
rect 22036 62586 22092 62588
rect 22116 62586 22172 62588
rect 22196 62586 22252 62588
rect 21956 62534 22002 62586
rect 22002 62534 22012 62586
rect 22036 62534 22066 62586
rect 22066 62534 22078 62586
rect 22078 62534 22092 62586
rect 22116 62534 22130 62586
rect 22130 62534 22142 62586
rect 22142 62534 22172 62586
rect 22196 62534 22206 62586
rect 22206 62534 22252 62586
rect 21956 62532 22012 62534
rect 22036 62532 22092 62534
rect 22116 62532 22172 62534
rect 22196 62532 22252 62534
rect 21956 61498 22012 61500
rect 22036 61498 22092 61500
rect 22116 61498 22172 61500
rect 22196 61498 22252 61500
rect 21956 61446 22002 61498
rect 22002 61446 22012 61498
rect 22036 61446 22066 61498
rect 22066 61446 22078 61498
rect 22078 61446 22092 61498
rect 22116 61446 22130 61498
rect 22130 61446 22142 61498
rect 22142 61446 22172 61498
rect 22196 61446 22206 61498
rect 22206 61446 22252 61498
rect 21956 61444 22012 61446
rect 22036 61444 22092 61446
rect 22116 61444 22172 61446
rect 22196 61444 22252 61446
rect 21956 60410 22012 60412
rect 22036 60410 22092 60412
rect 22116 60410 22172 60412
rect 22196 60410 22252 60412
rect 21956 60358 22002 60410
rect 22002 60358 22012 60410
rect 22036 60358 22066 60410
rect 22066 60358 22078 60410
rect 22078 60358 22092 60410
rect 22116 60358 22130 60410
rect 22130 60358 22142 60410
rect 22142 60358 22172 60410
rect 22196 60358 22206 60410
rect 22206 60358 22252 60410
rect 21956 60356 22012 60358
rect 22036 60356 22092 60358
rect 22116 60356 22172 60358
rect 22196 60356 22252 60358
rect 21956 59322 22012 59324
rect 22036 59322 22092 59324
rect 22116 59322 22172 59324
rect 22196 59322 22252 59324
rect 21956 59270 22002 59322
rect 22002 59270 22012 59322
rect 22036 59270 22066 59322
rect 22066 59270 22078 59322
rect 22078 59270 22092 59322
rect 22116 59270 22130 59322
rect 22130 59270 22142 59322
rect 22142 59270 22172 59322
rect 22196 59270 22206 59322
rect 22206 59270 22252 59322
rect 21956 59268 22012 59270
rect 22036 59268 22092 59270
rect 22116 59268 22172 59270
rect 22196 59268 22252 59270
rect 21956 58234 22012 58236
rect 22036 58234 22092 58236
rect 22116 58234 22172 58236
rect 22196 58234 22252 58236
rect 21956 58182 22002 58234
rect 22002 58182 22012 58234
rect 22036 58182 22066 58234
rect 22066 58182 22078 58234
rect 22078 58182 22092 58234
rect 22116 58182 22130 58234
rect 22130 58182 22142 58234
rect 22142 58182 22172 58234
rect 22196 58182 22206 58234
rect 22206 58182 22252 58234
rect 21956 58180 22012 58182
rect 22036 58180 22092 58182
rect 22116 58180 22172 58182
rect 22196 58180 22252 58182
rect 21956 57146 22012 57148
rect 22036 57146 22092 57148
rect 22116 57146 22172 57148
rect 22196 57146 22252 57148
rect 21956 57094 22002 57146
rect 22002 57094 22012 57146
rect 22036 57094 22066 57146
rect 22066 57094 22078 57146
rect 22078 57094 22092 57146
rect 22116 57094 22130 57146
rect 22130 57094 22142 57146
rect 22142 57094 22172 57146
rect 22196 57094 22206 57146
rect 22206 57094 22252 57146
rect 21956 57092 22012 57094
rect 22036 57092 22092 57094
rect 22116 57092 22172 57094
rect 22196 57092 22252 57094
rect 21956 56058 22012 56060
rect 22036 56058 22092 56060
rect 22116 56058 22172 56060
rect 22196 56058 22252 56060
rect 21956 56006 22002 56058
rect 22002 56006 22012 56058
rect 22036 56006 22066 56058
rect 22066 56006 22078 56058
rect 22078 56006 22092 56058
rect 22116 56006 22130 56058
rect 22130 56006 22142 56058
rect 22142 56006 22172 56058
rect 22196 56006 22206 56058
rect 22206 56006 22252 56058
rect 21956 56004 22012 56006
rect 22036 56004 22092 56006
rect 22116 56004 22172 56006
rect 22196 56004 22252 56006
rect 21956 54970 22012 54972
rect 22036 54970 22092 54972
rect 22116 54970 22172 54972
rect 22196 54970 22252 54972
rect 21956 54918 22002 54970
rect 22002 54918 22012 54970
rect 22036 54918 22066 54970
rect 22066 54918 22078 54970
rect 22078 54918 22092 54970
rect 22116 54918 22130 54970
rect 22130 54918 22142 54970
rect 22142 54918 22172 54970
rect 22196 54918 22206 54970
rect 22206 54918 22252 54970
rect 21956 54916 22012 54918
rect 22036 54916 22092 54918
rect 22116 54916 22172 54918
rect 22196 54916 22252 54918
rect 21956 53882 22012 53884
rect 22036 53882 22092 53884
rect 22116 53882 22172 53884
rect 22196 53882 22252 53884
rect 21956 53830 22002 53882
rect 22002 53830 22012 53882
rect 22036 53830 22066 53882
rect 22066 53830 22078 53882
rect 22078 53830 22092 53882
rect 22116 53830 22130 53882
rect 22130 53830 22142 53882
rect 22142 53830 22172 53882
rect 22196 53830 22206 53882
rect 22206 53830 22252 53882
rect 21956 53828 22012 53830
rect 22036 53828 22092 53830
rect 22116 53828 22172 53830
rect 22196 53828 22252 53830
rect 21956 52794 22012 52796
rect 22036 52794 22092 52796
rect 22116 52794 22172 52796
rect 22196 52794 22252 52796
rect 21956 52742 22002 52794
rect 22002 52742 22012 52794
rect 22036 52742 22066 52794
rect 22066 52742 22078 52794
rect 22078 52742 22092 52794
rect 22116 52742 22130 52794
rect 22130 52742 22142 52794
rect 22142 52742 22172 52794
rect 22196 52742 22206 52794
rect 22206 52742 22252 52794
rect 21956 52740 22012 52742
rect 22036 52740 22092 52742
rect 22116 52740 22172 52742
rect 22196 52740 22252 52742
rect 21956 51706 22012 51708
rect 22036 51706 22092 51708
rect 22116 51706 22172 51708
rect 22196 51706 22252 51708
rect 21956 51654 22002 51706
rect 22002 51654 22012 51706
rect 22036 51654 22066 51706
rect 22066 51654 22078 51706
rect 22078 51654 22092 51706
rect 22116 51654 22130 51706
rect 22130 51654 22142 51706
rect 22142 51654 22172 51706
rect 22196 51654 22206 51706
rect 22206 51654 22252 51706
rect 21956 51652 22012 51654
rect 22036 51652 22092 51654
rect 22116 51652 22172 51654
rect 22196 51652 22252 51654
rect 21956 50618 22012 50620
rect 22036 50618 22092 50620
rect 22116 50618 22172 50620
rect 22196 50618 22252 50620
rect 21956 50566 22002 50618
rect 22002 50566 22012 50618
rect 22036 50566 22066 50618
rect 22066 50566 22078 50618
rect 22078 50566 22092 50618
rect 22116 50566 22130 50618
rect 22130 50566 22142 50618
rect 22142 50566 22172 50618
rect 22196 50566 22206 50618
rect 22206 50566 22252 50618
rect 21956 50564 22012 50566
rect 22036 50564 22092 50566
rect 22116 50564 22172 50566
rect 22196 50564 22252 50566
rect 21956 49530 22012 49532
rect 22036 49530 22092 49532
rect 22116 49530 22172 49532
rect 22196 49530 22252 49532
rect 21956 49478 22002 49530
rect 22002 49478 22012 49530
rect 22036 49478 22066 49530
rect 22066 49478 22078 49530
rect 22078 49478 22092 49530
rect 22116 49478 22130 49530
rect 22130 49478 22142 49530
rect 22142 49478 22172 49530
rect 22196 49478 22206 49530
rect 22206 49478 22252 49530
rect 21956 49476 22012 49478
rect 22036 49476 22092 49478
rect 22116 49476 22172 49478
rect 22196 49476 22252 49478
rect 18878 7828 18880 7848
rect 18880 7828 18932 7848
rect 18932 7828 18934 7848
rect 18878 7792 18934 7828
rect 21956 48442 22012 48444
rect 22036 48442 22092 48444
rect 22116 48442 22172 48444
rect 22196 48442 22252 48444
rect 21956 48390 22002 48442
rect 22002 48390 22012 48442
rect 22036 48390 22066 48442
rect 22066 48390 22078 48442
rect 22078 48390 22092 48442
rect 22116 48390 22130 48442
rect 22130 48390 22142 48442
rect 22142 48390 22172 48442
rect 22196 48390 22206 48442
rect 22206 48390 22252 48442
rect 21956 48388 22012 48390
rect 22036 48388 22092 48390
rect 22116 48388 22172 48390
rect 22196 48388 22252 48390
rect 21956 47354 22012 47356
rect 22036 47354 22092 47356
rect 22116 47354 22172 47356
rect 22196 47354 22252 47356
rect 21956 47302 22002 47354
rect 22002 47302 22012 47354
rect 22036 47302 22066 47354
rect 22066 47302 22078 47354
rect 22078 47302 22092 47354
rect 22116 47302 22130 47354
rect 22130 47302 22142 47354
rect 22142 47302 22172 47354
rect 22196 47302 22206 47354
rect 22206 47302 22252 47354
rect 21956 47300 22012 47302
rect 22036 47300 22092 47302
rect 22116 47300 22172 47302
rect 22196 47300 22252 47302
rect 21956 46266 22012 46268
rect 22036 46266 22092 46268
rect 22116 46266 22172 46268
rect 22196 46266 22252 46268
rect 21956 46214 22002 46266
rect 22002 46214 22012 46266
rect 22036 46214 22066 46266
rect 22066 46214 22078 46266
rect 22078 46214 22092 46266
rect 22116 46214 22130 46266
rect 22130 46214 22142 46266
rect 22142 46214 22172 46266
rect 22196 46214 22206 46266
rect 22206 46214 22252 46266
rect 21956 46212 22012 46214
rect 22036 46212 22092 46214
rect 22116 46212 22172 46214
rect 22196 46212 22252 46214
rect 21956 45178 22012 45180
rect 22036 45178 22092 45180
rect 22116 45178 22172 45180
rect 22196 45178 22252 45180
rect 21956 45126 22002 45178
rect 22002 45126 22012 45178
rect 22036 45126 22066 45178
rect 22066 45126 22078 45178
rect 22078 45126 22092 45178
rect 22116 45126 22130 45178
rect 22130 45126 22142 45178
rect 22142 45126 22172 45178
rect 22196 45126 22206 45178
rect 22206 45126 22252 45178
rect 21956 45124 22012 45126
rect 22036 45124 22092 45126
rect 22116 45124 22172 45126
rect 22196 45124 22252 45126
rect 22616 64218 22672 64220
rect 22696 64218 22752 64220
rect 22776 64218 22832 64220
rect 22856 64218 22912 64220
rect 22616 64166 22662 64218
rect 22662 64166 22672 64218
rect 22696 64166 22726 64218
rect 22726 64166 22738 64218
rect 22738 64166 22752 64218
rect 22776 64166 22790 64218
rect 22790 64166 22802 64218
rect 22802 64166 22832 64218
rect 22856 64166 22866 64218
rect 22866 64166 22912 64218
rect 22616 64164 22672 64166
rect 22696 64164 22752 64166
rect 22776 64164 22832 64166
rect 22856 64164 22912 64166
rect 22616 63130 22672 63132
rect 22696 63130 22752 63132
rect 22776 63130 22832 63132
rect 22856 63130 22912 63132
rect 22616 63078 22662 63130
rect 22662 63078 22672 63130
rect 22696 63078 22726 63130
rect 22726 63078 22738 63130
rect 22738 63078 22752 63130
rect 22776 63078 22790 63130
rect 22790 63078 22802 63130
rect 22802 63078 22832 63130
rect 22856 63078 22866 63130
rect 22866 63078 22912 63130
rect 22616 63076 22672 63078
rect 22696 63076 22752 63078
rect 22776 63076 22832 63078
rect 22856 63076 22912 63078
rect 22616 62042 22672 62044
rect 22696 62042 22752 62044
rect 22776 62042 22832 62044
rect 22856 62042 22912 62044
rect 22616 61990 22662 62042
rect 22662 61990 22672 62042
rect 22696 61990 22726 62042
rect 22726 61990 22738 62042
rect 22738 61990 22752 62042
rect 22776 61990 22790 62042
rect 22790 61990 22802 62042
rect 22802 61990 22832 62042
rect 22856 61990 22866 62042
rect 22866 61990 22912 62042
rect 22616 61988 22672 61990
rect 22696 61988 22752 61990
rect 22776 61988 22832 61990
rect 22856 61988 22912 61990
rect 22616 60954 22672 60956
rect 22696 60954 22752 60956
rect 22776 60954 22832 60956
rect 22856 60954 22912 60956
rect 22616 60902 22662 60954
rect 22662 60902 22672 60954
rect 22696 60902 22726 60954
rect 22726 60902 22738 60954
rect 22738 60902 22752 60954
rect 22776 60902 22790 60954
rect 22790 60902 22802 60954
rect 22802 60902 22832 60954
rect 22856 60902 22866 60954
rect 22866 60902 22912 60954
rect 22616 60900 22672 60902
rect 22696 60900 22752 60902
rect 22776 60900 22832 60902
rect 22856 60900 22912 60902
rect 22616 59866 22672 59868
rect 22696 59866 22752 59868
rect 22776 59866 22832 59868
rect 22856 59866 22912 59868
rect 22616 59814 22662 59866
rect 22662 59814 22672 59866
rect 22696 59814 22726 59866
rect 22726 59814 22738 59866
rect 22738 59814 22752 59866
rect 22776 59814 22790 59866
rect 22790 59814 22802 59866
rect 22802 59814 22832 59866
rect 22856 59814 22866 59866
rect 22866 59814 22912 59866
rect 22616 59812 22672 59814
rect 22696 59812 22752 59814
rect 22776 59812 22832 59814
rect 22856 59812 22912 59814
rect 22616 58778 22672 58780
rect 22696 58778 22752 58780
rect 22776 58778 22832 58780
rect 22856 58778 22912 58780
rect 22616 58726 22662 58778
rect 22662 58726 22672 58778
rect 22696 58726 22726 58778
rect 22726 58726 22738 58778
rect 22738 58726 22752 58778
rect 22776 58726 22790 58778
rect 22790 58726 22802 58778
rect 22802 58726 22832 58778
rect 22856 58726 22866 58778
rect 22866 58726 22912 58778
rect 22616 58724 22672 58726
rect 22696 58724 22752 58726
rect 22776 58724 22832 58726
rect 22856 58724 22912 58726
rect 22616 57690 22672 57692
rect 22696 57690 22752 57692
rect 22776 57690 22832 57692
rect 22856 57690 22912 57692
rect 22616 57638 22662 57690
rect 22662 57638 22672 57690
rect 22696 57638 22726 57690
rect 22726 57638 22738 57690
rect 22738 57638 22752 57690
rect 22776 57638 22790 57690
rect 22790 57638 22802 57690
rect 22802 57638 22832 57690
rect 22856 57638 22866 57690
rect 22866 57638 22912 57690
rect 22616 57636 22672 57638
rect 22696 57636 22752 57638
rect 22776 57636 22832 57638
rect 22856 57636 22912 57638
rect 22616 56602 22672 56604
rect 22696 56602 22752 56604
rect 22776 56602 22832 56604
rect 22856 56602 22912 56604
rect 22616 56550 22662 56602
rect 22662 56550 22672 56602
rect 22696 56550 22726 56602
rect 22726 56550 22738 56602
rect 22738 56550 22752 56602
rect 22776 56550 22790 56602
rect 22790 56550 22802 56602
rect 22802 56550 22832 56602
rect 22856 56550 22866 56602
rect 22866 56550 22912 56602
rect 22616 56548 22672 56550
rect 22696 56548 22752 56550
rect 22776 56548 22832 56550
rect 22856 56548 22912 56550
rect 22616 55514 22672 55516
rect 22696 55514 22752 55516
rect 22776 55514 22832 55516
rect 22856 55514 22912 55516
rect 22616 55462 22662 55514
rect 22662 55462 22672 55514
rect 22696 55462 22726 55514
rect 22726 55462 22738 55514
rect 22738 55462 22752 55514
rect 22776 55462 22790 55514
rect 22790 55462 22802 55514
rect 22802 55462 22832 55514
rect 22856 55462 22866 55514
rect 22866 55462 22912 55514
rect 22616 55460 22672 55462
rect 22696 55460 22752 55462
rect 22776 55460 22832 55462
rect 22856 55460 22912 55462
rect 22616 54426 22672 54428
rect 22696 54426 22752 54428
rect 22776 54426 22832 54428
rect 22856 54426 22912 54428
rect 22616 54374 22662 54426
rect 22662 54374 22672 54426
rect 22696 54374 22726 54426
rect 22726 54374 22738 54426
rect 22738 54374 22752 54426
rect 22776 54374 22790 54426
rect 22790 54374 22802 54426
rect 22802 54374 22832 54426
rect 22856 54374 22866 54426
rect 22866 54374 22912 54426
rect 22616 54372 22672 54374
rect 22696 54372 22752 54374
rect 22776 54372 22832 54374
rect 22856 54372 22912 54374
rect 22616 53338 22672 53340
rect 22696 53338 22752 53340
rect 22776 53338 22832 53340
rect 22856 53338 22912 53340
rect 22616 53286 22662 53338
rect 22662 53286 22672 53338
rect 22696 53286 22726 53338
rect 22726 53286 22738 53338
rect 22738 53286 22752 53338
rect 22776 53286 22790 53338
rect 22790 53286 22802 53338
rect 22802 53286 22832 53338
rect 22856 53286 22866 53338
rect 22866 53286 22912 53338
rect 22616 53284 22672 53286
rect 22696 53284 22752 53286
rect 22776 53284 22832 53286
rect 22856 53284 22912 53286
rect 22616 52250 22672 52252
rect 22696 52250 22752 52252
rect 22776 52250 22832 52252
rect 22856 52250 22912 52252
rect 22616 52198 22662 52250
rect 22662 52198 22672 52250
rect 22696 52198 22726 52250
rect 22726 52198 22738 52250
rect 22738 52198 22752 52250
rect 22776 52198 22790 52250
rect 22790 52198 22802 52250
rect 22802 52198 22832 52250
rect 22856 52198 22866 52250
rect 22866 52198 22912 52250
rect 22616 52196 22672 52198
rect 22696 52196 22752 52198
rect 22776 52196 22832 52198
rect 22856 52196 22912 52198
rect 22616 51162 22672 51164
rect 22696 51162 22752 51164
rect 22776 51162 22832 51164
rect 22856 51162 22912 51164
rect 22616 51110 22662 51162
rect 22662 51110 22672 51162
rect 22696 51110 22726 51162
rect 22726 51110 22738 51162
rect 22738 51110 22752 51162
rect 22776 51110 22790 51162
rect 22790 51110 22802 51162
rect 22802 51110 22832 51162
rect 22856 51110 22866 51162
rect 22866 51110 22912 51162
rect 22616 51108 22672 51110
rect 22696 51108 22752 51110
rect 22776 51108 22832 51110
rect 22856 51108 22912 51110
rect 22616 50074 22672 50076
rect 22696 50074 22752 50076
rect 22776 50074 22832 50076
rect 22856 50074 22912 50076
rect 22616 50022 22662 50074
rect 22662 50022 22672 50074
rect 22696 50022 22726 50074
rect 22726 50022 22738 50074
rect 22738 50022 22752 50074
rect 22776 50022 22790 50074
rect 22790 50022 22802 50074
rect 22802 50022 22832 50074
rect 22856 50022 22866 50074
rect 22866 50022 22912 50074
rect 22616 50020 22672 50022
rect 22696 50020 22752 50022
rect 22776 50020 22832 50022
rect 22856 50020 22912 50022
rect 22616 48986 22672 48988
rect 22696 48986 22752 48988
rect 22776 48986 22832 48988
rect 22856 48986 22912 48988
rect 22616 48934 22662 48986
rect 22662 48934 22672 48986
rect 22696 48934 22726 48986
rect 22726 48934 22738 48986
rect 22738 48934 22752 48986
rect 22776 48934 22790 48986
rect 22790 48934 22802 48986
rect 22802 48934 22832 48986
rect 22856 48934 22866 48986
rect 22866 48934 22912 48986
rect 22616 48932 22672 48934
rect 22696 48932 22752 48934
rect 22776 48932 22832 48934
rect 22856 48932 22912 48934
rect 22616 47898 22672 47900
rect 22696 47898 22752 47900
rect 22776 47898 22832 47900
rect 22856 47898 22912 47900
rect 22616 47846 22662 47898
rect 22662 47846 22672 47898
rect 22696 47846 22726 47898
rect 22726 47846 22738 47898
rect 22738 47846 22752 47898
rect 22776 47846 22790 47898
rect 22790 47846 22802 47898
rect 22802 47846 22832 47898
rect 22856 47846 22866 47898
rect 22866 47846 22912 47898
rect 22616 47844 22672 47846
rect 22696 47844 22752 47846
rect 22776 47844 22832 47846
rect 22856 47844 22912 47846
rect 22616 46810 22672 46812
rect 22696 46810 22752 46812
rect 22776 46810 22832 46812
rect 22856 46810 22912 46812
rect 22616 46758 22662 46810
rect 22662 46758 22672 46810
rect 22696 46758 22726 46810
rect 22726 46758 22738 46810
rect 22738 46758 22752 46810
rect 22776 46758 22790 46810
rect 22790 46758 22802 46810
rect 22802 46758 22832 46810
rect 22856 46758 22866 46810
rect 22866 46758 22912 46810
rect 22616 46756 22672 46758
rect 22696 46756 22752 46758
rect 22776 46756 22832 46758
rect 22856 46756 22912 46758
rect 22616 45722 22672 45724
rect 22696 45722 22752 45724
rect 22776 45722 22832 45724
rect 22856 45722 22912 45724
rect 22616 45670 22662 45722
rect 22662 45670 22672 45722
rect 22696 45670 22726 45722
rect 22726 45670 22738 45722
rect 22738 45670 22752 45722
rect 22776 45670 22790 45722
rect 22790 45670 22802 45722
rect 22802 45670 22832 45722
rect 22856 45670 22866 45722
rect 22866 45670 22912 45722
rect 22616 45668 22672 45670
rect 22696 45668 22752 45670
rect 22776 45668 22832 45670
rect 22856 45668 22912 45670
rect 21956 44090 22012 44092
rect 22036 44090 22092 44092
rect 22116 44090 22172 44092
rect 22196 44090 22252 44092
rect 21956 44038 22002 44090
rect 22002 44038 22012 44090
rect 22036 44038 22066 44090
rect 22066 44038 22078 44090
rect 22078 44038 22092 44090
rect 22116 44038 22130 44090
rect 22130 44038 22142 44090
rect 22142 44038 22172 44090
rect 22196 44038 22206 44090
rect 22206 44038 22252 44090
rect 21956 44036 22012 44038
rect 22036 44036 22092 44038
rect 22116 44036 22172 44038
rect 22196 44036 22252 44038
rect 21956 43002 22012 43004
rect 22036 43002 22092 43004
rect 22116 43002 22172 43004
rect 22196 43002 22252 43004
rect 21956 42950 22002 43002
rect 22002 42950 22012 43002
rect 22036 42950 22066 43002
rect 22066 42950 22078 43002
rect 22078 42950 22092 43002
rect 22116 42950 22130 43002
rect 22130 42950 22142 43002
rect 22142 42950 22172 43002
rect 22196 42950 22206 43002
rect 22206 42950 22252 43002
rect 21956 42948 22012 42950
rect 22036 42948 22092 42950
rect 22116 42948 22172 42950
rect 22196 42948 22252 42950
rect 21956 41914 22012 41916
rect 22036 41914 22092 41916
rect 22116 41914 22172 41916
rect 22196 41914 22252 41916
rect 21956 41862 22002 41914
rect 22002 41862 22012 41914
rect 22036 41862 22066 41914
rect 22066 41862 22078 41914
rect 22078 41862 22092 41914
rect 22116 41862 22130 41914
rect 22130 41862 22142 41914
rect 22142 41862 22172 41914
rect 22196 41862 22206 41914
rect 22206 41862 22252 41914
rect 21956 41860 22012 41862
rect 22036 41860 22092 41862
rect 22116 41860 22172 41862
rect 22196 41860 22252 41862
rect 21956 40826 22012 40828
rect 22036 40826 22092 40828
rect 22116 40826 22172 40828
rect 22196 40826 22252 40828
rect 21956 40774 22002 40826
rect 22002 40774 22012 40826
rect 22036 40774 22066 40826
rect 22066 40774 22078 40826
rect 22078 40774 22092 40826
rect 22116 40774 22130 40826
rect 22130 40774 22142 40826
rect 22142 40774 22172 40826
rect 22196 40774 22206 40826
rect 22206 40774 22252 40826
rect 21956 40772 22012 40774
rect 22036 40772 22092 40774
rect 22116 40772 22172 40774
rect 22196 40772 22252 40774
rect 21956 39738 22012 39740
rect 22036 39738 22092 39740
rect 22116 39738 22172 39740
rect 22196 39738 22252 39740
rect 21956 39686 22002 39738
rect 22002 39686 22012 39738
rect 22036 39686 22066 39738
rect 22066 39686 22078 39738
rect 22078 39686 22092 39738
rect 22116 39686 22130 39738
rect 22130 39686 22142 39738
rect 22142 39686 22172 39738
rect 22196 39686 22206 39738
rect 22206 39686 22252 39738
rect 21956 39684 22012 39686
rect 22036 39684 22092 39686
rect 22116 39684 22172 39686
rect 22196 39684 22252 39686
rect 21956 38650 22012 38652
rect 22036 38650 22092 38652
rect 22116 38650 22172 38652
rect 22196 38650 22252 38652
rect 21956 38598 22002 38650
rect 22002 38598 22012 38650
rect 22036 38598 22066 38650
rect 22066 38598 22078 38650
rect 22078 38598 22092 38650
rect 22116 38598 22130 38650
rect 22130 38598 22142 38650
rect 22142 38598 22172 38650
rect 22196 38598 22206 38650
rect 22206 38598 22252 38650
rect 21956 38596 22012 38598
rect 22036 38596 22092 38598
rect 22116 38596 22172 38598
rect 22196 38596 22252 38598
rect 21956 37562 22012 37564
rect 22036 37562 22092 37564
rect 22116 37562 22172 37564
rect 22196 37562 22252 37564
rect 21956 37510 22002 37562
rect 22002 37510 22012 37562
rect 22036 37510 22066 37562
rect 22066 37510 22078 37562
rect 22078 37510 22092 37562
rect 22116 37510 22130 37562
rect 22130 37510 22142 37562
rect 22142 37510 22172 37562
rect 22196 37510 22206 37562
rect 22206 37510 22252 37562
rect 21956 37508 22012 37510
rect 22036 37508 22092 37510
rect 22116 37508 22172 37510
rect 22196 37508 22252 37510
rect 21956 36474 22012 36476
rect 22036 36474 22092 36476
rect 22116 36474 22172 36476
rect 22196 36474 22252 36476
rect 21956 36422 22002 36474
rect 22002 36422 22012 36474
rect 22036 36422 22066 36474
rect 22066 36422 22078 36474
rect 22078 36422 22092 36474
rect 22116 36422 22130 36474
rect 22130 36422 22142 36474
rect 22142 36422 22172 36474
rect 22196 36422 22206 36474
rect 22206 36422 22252 36474
rect 21956 36420 22012 36422
rect 22036 36420 22092 36422
rect 22116 36420 22172 36422
rect 22196 36420 22252 36422
rect 21956 35386 22012 35388
rect 22036 35386 22092 35388
rect 22116 35386 22172 35388
rect 22196 35386 22252 35388
rect 21956 35334 22002 35386
rect 22002 35334 22012 35386
rect 22036 35334 22066 35386
rect 22066 35334 22078 35386
rect 22078 35334 22092 35386
rect 22116 35334 22130 35386
rect 22130 35334 22142 35386
rect 22142 35334 22172 35386
rect 22196 35334 22206 35386
rect 22206 35334 22252 35386
rect 21956 35332 22012 35334
rect 22036 35332 22092 35334
rect 22116 35332 22172 35334
rect 22196 35332 22252 35334
rect 21956 34298 22012 34300
rect 22036 34298 22092 34300
rect 22116 34298 22172 34300
rect 22196 34298 22252 34300
rect 21956 34246 22002 34298
rect 22002 34246 22012 34298
rect 22036 34246 22066 34298
rect 22066 34246 22078 34298
rect 22078 34246 22092 34298
rect 22116 34246 22130 34298
rect 22130 34246 22142 34298
rect 22142 34246 22172 34298
rect 22196 34246 22206 34298
rect 22206 34246 22252 34298
rect 21956 34244 22012 34246
rect 22036 34244 22092 34246
rect 22116 34244 22172 34246
rect 22196 34244 22252 34246
rect 21956 33210 22012 33212
rect 22036 33210 22092 33212
rect 22116 33210 22172 33212
rect 22196 33210 22252 33212
rect 21956 33158 22002 33210
rect 22002 33158 22012 33210
rect 22036 33158 22066 33210
rect 22066 33158 22078 33210
rect 22078 33158 22092 33210
rect 22116 33158 22130 33210
rect 22130 33158 22142 33210
rect 22142 33158 22172 33210
rect 22196 33158 22206 33210
rect 22206 33158 22252 33210
rect 21956 33156 22012 33158
rect 22036 33156 22092 33158
rect 22116 33156 22172 33158
rect 22196 33156 22252 33158
rect 21956 32122 22012 32124
rect 22036 32122 22092 32124
rect 22116 32122 22172 32124
rect 22196 32122 22252 32124
rect 21956 32070 22002 32122
rect 22002 32070 22012 32122
rect 22036 32070 22066 32122
rect 22066 32070 22078 32122
rect 22078 32070 22092 32122
rect 22116 32070 22130 32122
rect 22130 32070 22142 32122
rect 22142 32070 22172 32122
rect 22196 32070 22206 32122
rect 22206 32070 22252 32122
rect 21956 32068 22012 32070
rect 22036 32068 22092 32070
rect 22116 32068 22172 32070
rect 22196 32068 22252 32070
rect 21956 31034 22012 31036
rect 22036 31034 22092 31036
rect 22116 31034 22172 31036
rect 22196 31034 22252 31036
rect 21956 30982 22002 31034
rect 22002 30982 22012 31034
rect 22036 30982 22066 31034
rect 22066 30982 22078 31034
rect 22078 30982 22092 31034
rect 22116 30982 22130 31034
rect 22130 30982 22142 31034
rect 22142 30982 22172 31034
rect 22196 30982 22206 31034
rect 22206 30982 22252 31034
rect 21956 30980 22012 30982
rect 22036 30980 22092 30982
rect 22116 30980 22172 30982
rect 22196 30980 22252 30982
rect 22616 44634 22672 44636
rect 22696 44634 22752 44636
rect 22776 44634 22832 44636
rect 22856 44634 22912 44636
rect 22616 44582 22662 44634
rect 22662 44582 22672 44634
rect 22696 44582 22726 44634
rect 22726 44582 22738 44634
rect 22738 44582 22752 44634
rect 22776 44582 22790 44634
rect 22790 44582 22802 44634
rect 22802 44582 22832 44634
rect 22856 44582 22866 44634
rect 22866 44582 22912 44634
rect 22616 44580 22672 44582
rect 22696 44580 22752 44582
rect 22776 44580 22832 44582
rect 22856 44580 22912 44582
rect 22616 43546 22672 43548
rect 22696 43546 22752 43548
rect 22776 43546 22832 43548
rect 22856 43546 22912 43548
rect 22616 43494 22662 43546
rect 22662 43494 22672 43546
rect 22696 43494 22726 43546
rect 22726 43494 22738 43546
rect 22738 43494 22752 43546
rect 22776 43494 22790 43546
rect 22790 43494 22802 43546
rect 22802 43494 22832 43546
rect 22856 43494 22866 43546
rect 22866 43494 22912 43546
rect 22616 43492 22672 43494
rect 22696 43492 22752 43494
rect 22776 43492 22832 43494
rect 22856 43492 22912 43494
rect 22616 42458 22672 42460
rect 22696 42458 22752 42460
rect 22776 42458 22832 42460
rect 22856 42458 22912 42460
rect 22616 42406 22662 42458
rect 22662 42406 22672 42458
rect 22696 42406 22726 42458
rect 22726 42406 22738 42458
rect 22738 42406 22752 42458
rect 22776 42406 22790 42458
rect 22790 42406 22802 42458
rect 22802 42406 22832 42458
rect 22856 42406 22866 42458
rect 22866 42406 22912 42458
rect 22616 42404 22672 42406
rect 22696 42404 22752 42406
rect 22776 42404 22832 42406
rect 22856 42404 22912 42406
rect 22616 41370 22672 41372
rect 22696 41370 22752 41372
rect 22776 41370 22832 41372
rect 22856 41370 22912 41372
rect 22616 41318 22662 41370
rect 22662 41318 22672 41370
rect 22696 41318 22726 41370
rect 22726 41318 22738 41370
rect 22738 41318 22752 41370
rect 22776 41318 22790 41370
rect 22790 41318 22802 41370
rect 22802 41318 22832 41370
rect 22856 41318 22866 41370
rect 22866 41318 22912 41370
rect 22616 41316 22672 41318
rect 22696 41316 22752 41318
rect 22776 41316 22832 41318
rect 22856 41316 22912 41318
rect 22616 40282 22672 40284
rect 22696 40282 22752 40284
rect 22776 40282 22832 40284
rect 22856 40282 22912 40284
rect 22616 40230 22662 40282
rect 22662 40230 22672 40282
rect 22696 40230 22726 40282
rect 22726 40230 22738 40282
rect 22738 40230 22752 40282
rect 22776 40230 22790 40282
rect 22790 40230 22802 40282
rect 22802 40230 22832 40282
rect 22856 40230 22866 40282
rect 22866 40230 22912 40282
rect 22616 40228 22672 40230
rect 22696 40228 22752 40230
rect 22776 40228 22832 40230
rect 22856 40228 22912 40230
rect 22616 39194 22672 39196
rect 22696 39194 22752 39196
rect 22776 39194 22832 39196
rect 22856 39194 22912 39196
rect 22616 39142 22662 39194
rect 22662 39142 22672 39194
rect 22696 39142 22726 39194
rect 22726 39142 22738 39194
rect 22738 39142 22752 39194
rect 22776 39142 22790 39194
rect 22790 39142 22802 39194
rect 22802 39142 22832 39194
rect 22856 39142 22866 39194
rect 22866 39142 22912 39194
rect 22616 39140 22672 39142
rect 22696 39140 22752 39142
rect 22776 39140 22832 39142
rect 22856 39140 22912 39142
rect 22616 38106 22672 38108
rect 22696 38106 22752 38108
rect 22776 38106 22832 38108
rect 22856 38106 22912 38108
rect 22616 38054 22662 38106
rect 22662 38054 22672 38106
rect 22696 38054 22726 38106
rect 22726 38054 22738 38106
rect 22738 38054 22752 38106
rect 22776 38054 22790 38106
rect 22790 38054 22802 38106
rect 22802 38054 22832 38106
rect 22856 38054 22866 38106
rect 22866 38054 22912 38106
rect 22616 38052 22672 38054
rect 22696 38052 22752 38054
rect 22776 38052 22832 38054
rect 22856 38052 22912 38054
rect 22616 37018 22672 37020
rect 22696 37018 22752 37020
rect 22776 37018 22832 37020
rect 22856 37018 22912 37020
rect 22616 36966 22662 37018
rect 22662 36966 22672 37018
rect 22696 36966 22726 37018
rect 22726 36966 22738 37018
rect 22738 36966 22752 37018
rect 22776 36966 22790 37018
rect 22790 36966 22802 37018
rect 22802 36966 22832 37018
rect 22856 36966 22866 37018
rect 22866 36966 22912 37018
rect 22616 36964 22672 36966
rect 22696 36964 22752 36966
rect 22776 36964 22832 36966
rect 22856 36964 22912 36966
rect 22616 35930 22672 35932
rect 22696 35930 22752 35932
rect 22776 35930 22832 35932
rect 22856 35930 22912 35932
rect 22616 35878 22662 35930
rect 22662 35878 22672 35930
rect 22696 35878 22726 35930
rect 22726 35878 22738 35930
rect 22738 35878 22752 35930
rect 22776 35878 22790 35930
rect 22790 35878 22802 35930
rect 22802 35878 22832 35930
rect 22856 35878 22866 35930
rect 22866 35878 22912 35930
rect 22616 35876 22672 35878
rect 22696 35876 22752 35878
rect 22776 35876 22832 35878
rect 22856 35876 22912 35878
rect 22616 34842 22672 34844
rect 22696 34842 22752 34844
rect 22776 34842 22832 34844
rect 22856 34842 22912 34844
rect 22616 34790 22662 34842
rect 22662 34790 22672 34842
rect 22696 34790 22726 34842
rect 22726 34790 22738 34842
rect 22738 34790 22752 34842
rect 22776 34790 22790 34842
rect 22790 34790 22802 34842
rect 22802 34790 22832 34842
rect 22856 34790 22866 34842
rect 22866 34790 22912 34842
rect 22616 34788 22672 34790
rect 22696 34788 22752 34790
rect 22776 34788 22832 34790
rect 22856 34788 22912 34790
rect 22616 33754 22672 33756
rect 22696 33754 22752 33756
rect 22776 33754 22832 33756
rect 22856 33754 22912 33756
rect 22616 33702 22662 33754
rect 22662 33702 22672 33754
rect 22696 33702 22726 33754
rect 22726 33702 22738 33754
rect 22738 33702 22752 33754
rect 22776 33702 22790 33754
rect 22790 33702 22802 33754
rect 22802 33702 22832 33754
rect 22856 33702 22866 33754
rect 22866 33702 22912 33754
rect 22616 33700 22672 33702
rect 22696 33700 22752 33702
rect 22776 33700 22832 33702
rect 22856 33700 22912 33702
rect 22616 32666 22672 32668
rect 22696 32666 22752 32668
rect 22776 32666 22832 32668
rect 22856 32666 22912 32668
rect 22616 32614 22662 32666
rect 22662 32614 22672 32666
rect 22696 32614 22726 32666
rect 22726 32614 22738 32666
rect 22738 32614 22752 32666
rect 22776 32614 22790 32666
rect 22790 32614 22802 32666
rect 22802 32614 22832 32666
rect 22856 32614 22866 32666
rect 22866 32614 22912 32666
rect 22616 32612 22672 32614
rect 22696 32612 22752 32614
rect 22776 32612 22832 32614
rect 22856 32612 22912 32614
rect 22616 31578 22672 31580
rect 22696 31578 22752 31580
rect 22776 31578 22832 31580
rect 22856 31578 22912 31580
rect 22616 31526 22662 31578
rect 22662 31526 22672 31578
rect 22696 31526 22726 31578
rect 22726 31526 22738 31578
rect 22738 31526 22752 31578
rect 22776 31526 22790 31578
rect 22790 31526 22802 31578
rect 22802 31526 22832 31578
rect 22856 31526 22866 31578
rect 22866 31526 22912 31578
rect 22616 31524 22672 31526
rect 22696 31524 22752 31526
rect 22776 31524 22832 31526
rect 22856 31524 22912 31526
rect 22616 30490 22672 30492
rect 22696 30490 22752 30492
rect 22776 30490 22832 30492
rect 22856 30490 22912 30492
rect 22616 30438 22662 30490
rect 22662 30438 22672 30490
rect 22696 30438 22726 30490
rect 22726 30438 22738 30490
rect 22738 30438 22752 30490
rect 22776 30438 22790 30490
rect 22790 30438 22802 30490
rect 22802 30438 22832 30490
rect 22856 30438 22866 30490
rect 22866 30438 22912 30490
rect 22616 30436 22672 30438
rect 22696 30436 22752 30438
rect 22776 30436 22832 30438
rect 22856 30436 22912 30438
rect 21956 29946 22012 29948
rect 22036 29946 22092 29948
rect 22116 29946 22172 29948
rect 22196 29946 22252 29948
rect 21956 29894 22002 29946
rect 22002 29894 22012 29946
rect 22036 29894 22066 29946
rect 22066 29894 22078 29946
rect 22078 29894 22092 29946
rect 22116 29894 22130 29946
rect 22130 29894 22142 29946
rect 22142 29894 22172 29946
rect 22196 29894 22206 29946
rect 22206 29894 22252 29946
rect 21956 29892 22012 29894
rect 22036 29892 22092 29894
rect 22116 29892 22172 29894
rect 22196 29892 22252 29894
rect 22616 29402 22672 29404
rect 22696 29402 22752 29404
rect 22776 29402 22832 29404
rect 22856 29402 22912 29404
rect 22616 29350 22662 29402
rect 22662 29350 22672 29402
rect 22696 29350 22726 29402
rect 22726 29350 22738 29402
rect 22738 29350 22752 29402
rect 22776 29350 22790 29402
rect 22790 29350 22802 29402
rect 22802 29350 22832 29402
rect 22856 29350 22866 29402
rect 22866 29350 22912 29402
rect 22616 29348 22672 29350
rect 22696 29348 22752 29350
rect 22776 29348 22832 29350
rect 22856 29348 22912 29350
rect 21956 28858 22012 28860
rect 22036 28858 22092 28860
rect 22116 28858 22172 28860
rect 22196 28858 22252 28860
rect 21956 28806 22002 28858
rect 22002 28806 22012 28858
rect 22036 28806 22066 28858
rect 22066 28806 22078 28858
rect 22078 28806 22092 28858
rect 22116 28806 22130 28858
rect 22130 28806 22142 28858
rect 22142 28806 22172 28858
rect 22196 28806 22206 28858
rect 22206 28806 22252 28858
rect 21956 28804 22012 28806
rect 22036 28804 22092 28806
rect 22116 28804 22172 28806
rect 22196 28804 22252 28806
rect 22616 28314 22672 28316
rect 22696 28314 22752 28316
rect 22776 28314 22832 28316
rect 22856 28314 22912 28316
rect 22616 28262 22662 28314
rect 22662 28262 22672 28314
rect 22696 28262 22726 28314
rect 22726 28262 22738 28314
rect 22738 28262 22752 28314
rect 22776 28262 22790 28314
rect 22790 28262 22802 28314
rect 22802 28262 22832 28314
rect 22856 28262 22866 28314
rect 22866 28262 22912 28314
rect 22616 28260 22672 28262
rect 22696 28260 22752 28262
rect 22776 28260 22832 28262
rect 22856 28260 22912 28262
rect 21956 27770 22012 27772
rect 22036 27770 22092 27772
rect 22116 27770 22172 27772
rect 22196 27770 22252 27772
rect 21956 27718 22002 27770
rect 22002 27718 22012 27770
rect 22036 27718 22066 27770
rect 22066 27718 22078 27770
rect 22078 27718 22092 27770
rect 22116 27718 22130 27770
rect 22130 27718 22142 27770
rect 22142 27718 22172 27770
rect 22196 27718 22206 27770
rect 22206 27718 22252 27770
rect 21956 27716 22012 27718
rect 22036 27716 22092 27718
rect 22116 27716 22172 27718
rect 22196 27716 22252 27718
rect 21956 26682 22012 26684
rect 22036 26682 22092 26684
rect 22116 26682 22172 26684
rect 22196 26682 22252 26684
rect 21956 26630 22002 26682
rect 22002 26630 22012 26682
rect 22036 26630 22066 26682
rect 22066 26630 22078 26682
rect 22078 26630 22092 26682
rect 22116 26630 22130 26682
rect 22130 26630 22142 26682
rect 22142 26630 22172 26682
rect 22196 26630 22206 26682
rect 22206 26630 22252 26682
rect 21956 26628 22012 26630
rect 22036 26628 22092 26630
rect 22116 26628 22172 26630
rect 22196 26628 22252 26630
rect 21956 25594 22012 25596
rect 22036 25594 22092 25596
rect 22116 25594 22172 25596
rect 22196 25594 22252 25596
rect 21956 25542 22002 25594
rect 22002 25542 22012 25594
rect 22036 25542 22066 25594
rect 22066 25542 22078 25594
rect 22078 25542 22092 25594
rect 22116 25542 22130 25594
rect 22130 25542 22142 25594
rect 22142 25542 22172 25594
rect 22196 25542 22206 25594
rect 22206 25542 22252 25594
rect 21956 25540 22012 25542
rect 22036 25540 22092 25542
rect 22116 25540 22172 25542
rect 22196 25540 22252 25542
rect 21956 24506 22012 24508
rect 22036 24506 22092 24508
rect 22116 24506 22172 24508
rect 22196 24506 22252 24508
rect 21956 24454 22002 24506
rect 22002 24454 22012 24506
rect 22036 24454 22066 24506
rect 22066 24454 22078 24506
rect 22078 24454 22092 24506
rect 22116 24454 22130 24506
rect 22130 24454 22142 24506
rect 22142 24454 22172 24506
rect 22196 24454 22206 24506
rect 22206 24454 22252 24506
rect 21956 24452 22012 24454
rect 22036 24452 22092 24454
rect 22116 24452 22172 24454
rect 22196 24452 22252 24454
rect 21956 23418 22012 23420
rect 22036 23418 22092 23420
rect 22116 23418 22172 23420
rect 22196 23418 22252 23420
rect 21956 23366 22002 23418
rect 22002 23366 22012 23418
rect 22036 23366 22066 23418
rect 22066 23366 22078 23418
rect 22078 23366 22092 23418
rect 22116 23366 22130 23418
rect 22130 23366 22142 23418
rect 22142 23366 22172 23418
rect 22196 23366 22206 23418
rect 22206 23366 22252 23418
rect 21956 23364 22012 23366
rect 22036 23364 22092 23366
rect 22116 23364 22172 23366
rect 22196 23364 22252 23366
rect 21956 22330 22012 22332
rect 22036 22330 22092 22332
rect 22116 22330 22172 22332
rect 22196 22330 22252 22332
rect 21956 22278 22002 22330
rect 22002 22278 22012 22330
rect 22036 22278 22066 22330
rect 22066 22278 22078 22330
rect 22078 22278 22092 22330
rect 22116 22278 22130 22330
rect 22130 22278 22142 22330
rect 22142 22278 22172 22330
rect 22196 22278 22206 22330
rect 22206 22278 22252 22330
rect 21956 22276 22012 22278
rect 22036 22276 22092 22278
rect 22116 22276 22172 22278
rect 22196 22276 22252 22278
rect 21956 21242 22012 21244
rect 22036 21242 22092 21244
rect 22116 21242 22172 21244
rect 22196 21242 22252 21244
rect 21956 21190 22002 21242
rect 22002 21190 22012 21242
rect 22036 21190 22066 21242
rect 22066 21190 22078 21242
rect 22078 21190 22092 21242
rect 22116 21190 22130 21242
rect 22130 21190 22142 21242
rect 22142 21190 22172 21242
rect 22196 21190 22206 21242
rect 22206 21190 22252 21242
rect 21956 21188 22012 21190
rect 22036 21188 22092 21190
rect 22116 21188 22172 21190
rect 22196 21188 22252 21190
rect 21956 20154 22012 20156
rect 22036 20154 22092 20156
rect 22116 20154 22172 20156
rect 22196 20154 22252 20156
rect 21956 20102 22002 20154
rect 22002 20102 22012 20154
rect 22036 20102 22066 20154
rect 22066 20102 22078 20154
rect 22078 20102 22092 20154
rect 22116 20102 22130 20154
rect 22130 20102 22142 20154
rect 22142 20102 22172 20154
rect 22196 20102 22206 20154
rect 22206 20102 22252 20154
rect 21956 20100 22012 20102
rect 22036 20100 22092 20102
rect 22116 20100 22172 20102
rect 22196 20100 22252 20102
rect 21956 19066 22012 19068
rect 22036 19066 22092 19068
rect 22116 19066 22172 19068
rect 22196 19066 22252 19068
rect 21956 19014 22002 19066
rect 22002 19014 22012 19066
rect 22036 19014 22066 19066
rect 22066 19014 22078 19066
rect 22078 19014 22092 19066
rect 22116 19014 22130 19066
rect 22130 19014 22142 19066
rect 22142 19014 22172 19066
rect 22196 19014 22206 19066
rect 22206 19014 22252 19066
rect 21956 19012 22012 19014
rect 22036 19012 22092 19014
rect 22116 19012 22172 19014
rect 22196 19012 22252 19014
rect 21956 17978 22012 17980
rect 22036 17978 22092 17980
rect 22116 17978 22172 17980
rect 22196 17978 22252 17980
rect 21956 17926 22002 17978
rect 22002 17926 22012 17978
rect 22036 17926 22066 17978
rect 22066 17926 22078 17978
rect 22078 17926 22092 17978
rect 22116 17926 22130 17978
rect 22130 17926 22142 17978
rect 22142 17926 22172 17978
rect 22196 17926 22206 17978
rect 22206 17926 22252 17978
rect 21956 17924 22012 17926
rect 22036 17924 22092 17926
rect 22116 17924 22172 17926
rect 22196 17924 22252 17926
rect 21956 16890 22012 16892
rect 22036 16890 22092 16892
rect 22116 16890 22172 16892
rect 22196 16890 22252 16892
rect 21956 16838 22002 16890
rect 22002 16838 22012 16890
rect 22036 16838 22066 16890
rect 22066 16838 22078 16890
rect 22078 16838 22092 16890
rect 22116 16838 22130 16890
rect 22130 16838 22142 16890
rect 22142 16838 22172 16890
rect 22196 16838 22206 16890
rect 22206 16838 22252 16890
rect 21956 16836 22012 16838
rect 22036 16836 22092 16838
rect 22116 16836 22172 16838
rect 22196 16836 22252 16838
rect 21956 15802 22012 15804
rect 22036 15802 22092 15804
rect 22116 15802 22172 15804
rect 22196 15802 22252 15804
rect 21956 15750 22002 15802
rect 22002 15750 22012 15802
rect 22036 15750 22066 15802
rect 22066 15750 22078 15802
rect 22078 15750 22092 15802
rect 22116 15750 22130 15802
rect 22130 15750 22142 15802
rect 22142 15750 22172 15802
rect 22196 15750 22206 15802
rect 22206 15750 22252 15802
rect 21956 15748 22012 15750
rect 22036 15748 22092 15750
rect 22116 15748 22172 15750
rect 22196 15748 22252 15750
rect 21956 14714 22012 14716
rect 22036 14714 22092 14716
rect 22116 14714 22172 14716
rect 22196 14714 22252 14716
rect 21956 14662 22002 14714
rect 22002 14662 22012 14714
rect 22036 14662 22066 14714
rect 22066 14662 22078 14714
rect 22078 14662 22092 14714
rect 22116 14662 22130 14714
rect 22130 14662 22142 14714
rect 22142 14662 22172 14714
rect 22196 14662 22206 14714
rect 22206 14662 22252 14714
rect 21956 14660 22012 14662
rect 22036 14660 22092 14662
rect 22116 14660 22172 14662
rect 22196 14660 22252 14662
rect 21956 13626 22012 13628
rect 22036 13626 22092 13628
rect 22116 13626 22172 13628
rect 22196 13626 22252 13628
rect 21956 13574 22002 13626
rect 22002 13574 22012 13626
rect 22036 13574 22066 13626
rect 22066 13574 22078 13626
rect 22078 13574 22092 13626
rect 22116 13574 22130 13626
rect 22130 13574 22142 13626
rect 22142 13574 22172 13626
rect 22196 13574 22206 13626
rect 22206 13574 22252 13626
rect 21956 13572 22012 13574
rect 22036 13572 22092 13574
rect 22116 13572 22172 13574
rect 22196 13572 22252 13574
rect 21956 12538 22012 12540
rect 22036 12538 22092 12540
rect 22116 12538 22172 12540
rect 22196 12538 22252 12540
rect 21956 12486 22002 12538
rect 22002 12486 22012 12538
rect 22036 12486 22066 12538
rect 22066 12486 22078 12538
rect 22078 12486 22092 12538
rect 22116 12486 22130 12538
rect 22130 12486 22142 12538
rect 22142 12486 22172 12538
rect 22196 12486 22206 12538
rect 22206 12486 22252 12538
rect 21956 12484 22012 12486
rect 22036 12484 22092 12486
rect 22116 12484 22172 12486
rect 22196 12484 22252 12486
rect 21956 11450 22012 11452
rect 22036 11450 22092 11452
rect 22116 11450 22172 11452
rect 22196 11450 22252 11452
rect 21956 11398 22002 11450
rect 22002 11398 22012 11450
rect 22036 11398 22066 11450
rect 22066 11398 22078 11450
rect 22078 11398 22092 11450
rect 22116 11398 22130 11450
rect 22130 11398 22142 11450
rect 22142 11398 22172 11450
rect 22196 11398 22206 11450
rect 22206 11398 22252 11450
rect 21956 11396 22012 11398
rect 22036 11396 22092 11398
rect 22116 11396 22172 11398
rect 22196 11396 22252 11398
rect 21956 10362 22012 10364
rect 22036 10362 22092 10364
rect 22116 10362 22172 10364
rect 22196 10362 22252 10364
rect 21956 10310 22002 10362
rect 22002 10310 22012 10362
rect 22036 10310 22066 10362
rect 22066 10310 22078 10362
rect 22078 10310 22092 10362
rect 22116 10310 22130 10362
rect 22130 10310 22142 10362
rect 22142 10310 22172 10362
rect 22196 10310 22206 10362
rect 22206 10310 22252 10362
rect 21956 10308 22012 10310
rect 22036 10308 22092 10310
rect 22116 10308 22172 10310
rect 22196 10308 22252 10310
rect 21956 9274 22012 9276
rect 22036 9274 22092 9276
rect 22116 9274 22172 9276
rect 22196 9274 22252 9276
rect 21956 9222 22002 9274
rect 22002 9222 22012 9274
rect 22036 9222 22066 9274
rect 22066 9222 22078 9274
rect 22078 9222 22092 9274
rect 22116 9222 22130 9274
rect 22130 9222 22142 9274
rect 22142 9222 22172 9274
rect 22196 9222 22206 9274
rect 22206 9222 22252 9274
rect 21956 9220 22012 9222
rect 22036 9220 22092 9222
rect 22116 9220 22172 9222
rect 22196 9220 22252 9222
rect 22616 27226 22672 27228
rect 22696 27226 22752 27228
rect 22776 27226 22832 27228
rect 22856 27226 22912 27228
rect 22616 27174 22662 27226
rect 22662 27174 22672 27226
rect 22696 27174 22726 27226
rect 22726 27174 22738 27226
rect 22738 27174 22752 27226
rect 22776 27174 22790 27226
rect 22790 27174 22802 27226
rect 22802 27174 22832 27226
rect 22856 27174 22866 27226
rect 22866 27174 22912 27226
rect 22616 27172 22672 27174
rect 22696 27172 22752 27174
rect 22776 27172 22832 27174
rect 22856 27172 22912 27174
rect 22616 26138 22672 26140
rect 22696 26138 22752 26140
rect 22776 26138 22832 26140
rect 22856 26138 22912 26140
rect 22616 26086 22662 26138
rect 22662 26086 22672 26138
rect 22696 26086 22726 26138
rect 22726 26086 22738 26138
rect 22738 26086 22752 26138
rect 22776 26086 22790 26138
rect 22790 26086 22802 26138
rect 22802 26086 22832 26138
rect 22856 26086 22866 26138
rect 22866 26086 22912 26138
rect 22616 26084 22672 26086
rect 22696 26084 22752 26086
rect 22776 26084 22832 26086
rect 22856 26084 22912 26086
rect 22616 25050 22672 25052
rect 22696 25050 22752 25052
rect 22776 25050 22832 25052
rect 22856 25050 22912 25052
rect 22616 24998 22662 25050
rect 22662 24998 22672 25050
rect 22696 24998 22726 25050
rect 22726 24998 22738 25050
rect 22738 24998 22752 25050
rect 22776 24998 22790 25050
rect 22790 24998 22802 25050
rect 22802 24998 22832 25050
rect 22856 24998 22866 25050
rect 22866 24998 22912 25050
rect 22616 24996 22672 24998
rect 22696 24996 22752 24998
rect 22776 24996 22832 24998
rect 22856 24996 22912 24998
rect 22616 23962 22672 23964
rect 22696 23962 22752 23964
rect 22776 23962 22832 23964
rect 22856 23962 22912 23964
rect 22616 23910 22662 23962
rect 22662 23910 22672 23962
rect 22696 23910 22726 23962
rect 22726 23910 22738 23962
rect 22738 23910 22752 23962
rect 22776 23910 22790 23962
rect 22790 23910 22802 23962
rect 22802 23910 22832 23962
rect 22856 23910 22866 23962
rect 22866 23910 22912 23962
rect 22616 23908 22672 23910
rect 22696 23908 22752 23910
rect 22776 23908 22832 23910
rect 22856 23908 22912 23910
rect 22616 22874 22672 22876
rect 22696 22874 22752 22876
rect 22776 22874 22832 22876
rect 22856 22874 22912 22876
rect 22616 22822 22662 22874
rect 22662 22822 22672 22874
rect 22696 22822 22726 22874
rect 22726 22822 22738 22874
rect 22738 22822 22752 22874
rect 22776 22822 22790 22874
rect 22790 22822 22802 22874
rect 22802 22822 22832 22874
rect 22856 22822 22866 22874
rect 22866 22822 22912 22874
rect 22616 22820 22672 22822
rect 22696 22820 22752 22822
rect 22776 22820 22832 22822
rect 22856 22820 22912 22822
rect 22616 21786 22672 21788
rect 22696 21786 22752 21788
rect 22776 21786 22832 21788
rect 22856 21786 22912 21788
rect 22616 21734 22662 21786
rect 22662 21734 22672 21786
rect 22696 21734 22726 21786
rect 22726 21734 22738 21786
rect 22738 21734 22752 21786
rect 22776 21734 22790 21786
rect 22790 21734 22802 21786
rect 22802 21734 22832 21786
rect 22856 21734 22866 21786
rect 22866 21734 22912 21786
rect 22616 21732 22672 21734
rect 22696 21732 22752 21734
rect 22776 21732 22832 21734
rect 22856 21732 22912 21734
rect 22616 20698 22672 20700
rect 22696 20698 22752 20700
rect 22776 20698 22832 20700
rect 22856 20698 22912 20700
rect 22616 20646 22662 20698
rect 22662 20646 22672 20698
rect 22696 20646 22726 20698
rect 22726 20646 22738 20698
rect 22738 20646 22752 20698
rect 22776 20646 22790 20698
rect 22790 20646 22802 20698
rect 22802 20646 22832 20698
rect 22856 20646 22866 20698
rect 22866 20646 22912 20698
rect 22616 20644 22672 20646
rect 22696 20644 22752 20646
rect 22776 20644 22832 20646
rect 22856 20644 22912 20646
rect 22616 19610 22672 19612
rect 22696 19610 22752 19612
rect 22776 19610 22832 19612
rect 22856 19610 22912 19612
rect 22616 19558 22662 19610
rect 22662 19558 22672 19610
rect 22696 19558 22726 19610
rect 22726 19558 22738 19610
rect 22738 19558 22752 19610
rect 22776 19558 22790 19610
rect 22790 19558 22802 19610
rect 22802 19558 22832 19610
rect 22856 19558 22866 19610
rect 22866 19558 22912 19610
rect 22616 19556 22672 19558
rect 22696 19556 22752 19558
rect 22776 19556 22832 19558
rect 22856 19556 22912 19558
rect 22616 18522 22672 18524
rect 22696 18522 22752 18524
rect 22776 18522 22832 18524
rect 22856 18522 22912 18524
rect 22616 18470 22662 18522
rect 22662 18470 22672 18522
rect 22696 18470 22726 18522
rect 22726 18470 22738 18522
rect 22738 18470 22752 18522
rect 22776 18470 22790 18522
rect 22790 18470 22802 18522
rect 22802 18470 22832 18522
rect 22856 18470 22866 18522
rect 22866 18470 22912 18522
rect 22616 18468 22672 18470
rect 22696 18468 22752 18470
rect 22776 18468 22832 18470
rect 22856 18468 22912 18470
rect 22616 17434 22672 17436
rect 22696 17434 22752 17436
rect 22776 17434 22832 17436
rect 22856 17434 22912 17436
rect 22616 17382 22662 17434
rect 22662 17382 22672 17434
rect 22696 17382 22726 17434
rect 22726 17382 22738 17434
rect 22738 17382 22752 17434
rect 22776 17382 22790 17434
rect 22790 17382 22802 17434
rect 22802 17382 22832 17434
rect 22856 17382 22866 17434
rect 22866 17382 22912 17434
rect 22616 17380 22672 17382
rect 22696 17380 22752 17382
rect 22776 17380 22832 17382
rect 22856 17380 22912 17382
rect 22616 16346 22672 16348
rect 22696 16346 22752 16348
rect 22776 16346 22832 16348
rect 22856 16346 22912 16348
rect 22616 16294 22662 16346
rect 22662 16294 22672 16346
rect 22696 16294 22726 16346
rect 22726 16294 22738 16346
rect 22738 16294 22752 16346
rect 22776 16294 22790 16346
rect 22790 16294 22802 16346
rect 22802 16294 22832 16346
rect 22856 16294 22866 16346
rect 22866 16294 22912 16346
rect 22616 16292 22672 16294
rect 22696 16292 22752 16294
rect 22776 16292 22832 16294
rect 22856 16292 22912 16294
rect 22616 15258 22672 15260
rect 22696 15258 22752 15260
rect 22776 15258 22832 15260
rect 22856 15258 22912 15260
rect 22616 15206 22662 15258
rect 22662 15206 22672 15258
rect 22696 15206 22726 15258
rect 22726 15206 22738 15258
rect 22738 15206 22752 15258
rect 22776 15206 22790 15258
rect 22790 15206 22802 15258
rect 22802 15206 22832 15258
rect 22856 15206 22866 15258
rect 22866 15206 22912 15258
rect 22616 15204 22672 15206
rect 22696 15204 22752 15206
rect 22776 15204 22832 15206
rect 22856 15204 22912 15206
rect 22616 14170 22672 14172
rect 22696 14170 22752 14172
rect 22776 14170 22832 14172
rect 22856 14170 22912 14172
rect 22616 14118 22662 14170
rect 22662 14118 22672 14170
rect 22696 14118 22726 14170
rect 22726 14118 22738 14170
rect 22738 14118 22752 14170
rect 22776 14118 22790 14170
rect 22790 14118 22802 14170
rect 22802 14118 22832 14170
rect 22856 14118 22866 14170
rect 22866 14118 22912 14170
rect 22616 14116 22672 14118
rect 22696 14116 22752 14118
rect 22776 14116 22832 14118
rect 22856 14116 22912 14118
rect 22616 13082 22672 13084
rect 22696 13082 22752 13084
rect 22776 13082 22832 13084
rect 22856 13082 22912 13084
rect 22616 13030 22662 13082
rect 22662 13030 22672 13082
rect 22696 13030 22726 13082
rect 22726 13030 22738 13082
rect 22738 13030 22752 13082
rect 22776 13030 22790 13082
rect 22790 13030 22802 13082
rect 22802 13030 22832 13082
rect 22856 13030 22866 13082
rect 22866 13030 22912 13082
rect 22616 13028 22672 13030
rect 22696 13028 22752 13030
rect 22776 13028 22832 13030
rect 22856 13028 22912 13030
rect 26956 66938 27012 66940
rect 27036 66938 27092 66940
rect 27116 66938 27172 66940
rect 27196 66938 27252 66940
rect 26956 66886 27002 66938
rect 27002 66886 27012 66938
rect 27036 66886 27066 66938
rect 27066 66886 27078 66938
rect 27078 66886 27092 66938
rect 27116 66886 27130 66938
rect 27130 66886 27142 66938
rect 27142 66886 27172 66938
rect 27196 66886 27206 66938
rect 27206 66886 27252 66938
rect 26956 66884 27012 66886
rect 27036 66884 27092 66886
rect 27116 66884 27172 66886
rect 27196 66884 27252 66886
rect 24582 22652 24584 22672
rect 24584 22652 24636 22672
rect 24636 22652 24638 22672
rect 24582 22616 24638 22652
rect 26956 65850 27012 65852
rect 27036 65850 27092 65852
rect 27116 65850 27172 65852
rect 27196 65850 27252 65852
rect 26956 65798 27002 65850
rect 27002 65798 27012 65850
rect 27036 65798 27066 65850
rect 27066 65798 27078 65850
rect 27078 65798 27092 65850
rect 27116 65798 27130 65850
rect 27130 65798 27142 65850
rect 27142 65798 27172 65850
rect 27196 65798 27206 65850
rect 27206 65798 27252 65850
rect 26956 65796 27012 65798
rect 27036 65796 27092 65798
rect 27116 65796 27172 65798
rect 27196 65796 27252 65798
rect 26956 64762 27012 64764
rect 27036 64762 27092 64764
rect 27116 64762 27172 64764
rect 27196 64762 27252 64764
rect 26956 64710 27002 64762
rect 27002 64710 27012 64762
rect 27036 64710 27066 64762
rect 27066 64710 27078 64762
rect 27078 64710 27092 64762
rect 27116 64710 27130 64762
rect 27130 64710 27142 64762
rect 27142 64710 27172 64762
rect 27196 64710 27206 64762
rect 27206 64710 27252 64762
rect 26956 64708 27012 64710
rect 27036 64708 27092 64710
rect 27116 64708 27172 64710
rect 27196 64708 27252 64710
rect 26956 63674 27012 63676
rect 27036 63674 27092 63676
rect 27116 63674 27172 63676
rect 27196 63674 27252 63676
rect 26956 63622 27002 63674
rect 27002 63622 27012 63674
rect 27036 63622 27066 63674
rect 27066 63622 27078 63674
rect 27078 63622 27092 63674
rect 27116 63622 27130 63674
rect 27130 63622 27142 63674
rect 27142 63622 27172 63674
rect 27196 63622 27206 63674
rect 27206 63622 27252 63674
rect 26956 63620 27012 63622
rect 27036 63620 27092 63622
rect 27116 63620 27172 63622
rect 27196 63620 27252 63622
rect 26956 62586 27012 62588
rect 27036 62586 27092 62588
rect 27116 62586 27172 62588
rect 27196 62586 27252 62588
rect 26956 62534 27002 62586
rect 27002 62534 27012 62586
rect 27036 62534 27066 62586
rect 27066 62534 27078 62586
rect 27078 62534 27092 62586
rect 27116 62534 27130 62586
rect 27130 62534 27142 62586
rect 27142 62534 27172 62586
rect 27196 62534 27206 62586
rect 27206 62534 27252 62586
rect 26956 62532 27012 62534
rect 27036 62532 27092 62534
rect 27116 62532 27172 62534
rect 27196 62532 27252 62534
rect 22616 11994 22672 11996
rect 22696 11994 22752 11996
rect 22776 11994 22832 11996
rect 22856 11994 22912 11996
rect 22616 11942 22662 11994
rect 22662 11942 22672 11994
rect 22696 11942 22726 11994
rect 22726 11942 22738 11994
rect 22738 11942 22752 11994
rect 22776 11942 22790 11994
rect 22790 11942 22802 11994
rect 22802 11942 22832 11994
rect 22856 11942 22866 11994
rect 22866 11942 22912 11994
rect 22616 11940 22672 11942
rect 22696 11940 22752 11942
rect 22776 11940 22832 11942
rect 22856 11940 22912 11942
rect 22616 10906 22672 10908
rect 22696 10906 22752 10908
rect 22776 10906 22832 10908
rect 22856 10906 22912 10908
rect 22616 10854 22662 10906
rect 22662 10854 22672 10906
rect 22696 10854 22726 10906
rect 22726 10854 22738 10906
rect 22738 10854 22752 10906
rect 22776 10854 22790 10906
rect 22790 10854 22802 10906
rect 22802 10854 22832 10906
rect 22856 10854 22866 10906
rect 22866 10854 22912 10906
rect 22616 10852 22672 10854
rect 22696 10852 22752 10854
rect 22776 10852 22832 10854
rect 22856 10852 22912 10854
rect 22616 9818 22672 9820
rect 22696 9818 22752 9820
rect 22776 9818 22832 9820
rect 22856 9818 22912 9820
rect 22616 9766 22662 9818
rect 22662 9766 22672 9818
rect 22696 9766 22726 9818
rect 22726 9766 22738 9818
rect 22738 9766 22752 9818
rect 22776 9766 22790 9818
rect 22790 9766 22802 9818
rect 22802 9766 22832 9818
rect 22856 9766 22866 9818
rect 22866 9766 22912 9818
rect 22616 9764 22672 9766
rect 22696 9764 22752 9766
rect 22776 9764 22832 9766
rect 22856 9764 22912 9766
rect 22616 8730 22672 8732
rect 22696 8730 22752 8732
rect 22776 8730 22832 8732
rect 22856 8730 22912 8732
rect 22616 8678 22662 8730
rect 22662 8678 22672 8730
rect 22696 8678 22726 8730
rect 22726 8678 22738 8730
rect 22738 8678 22752 8730
rect 22776 8678 22790 8730
rect 22790 8678 22802 8730
rect 22802 8678 22832 8730
rect 22856 8678 22866 8730
rect 22866 8678 22912 8730
rect 22616 8676 22672 8678
rect 22696 8676 22752 8678
rect 22776 8676 22832 8678
rect 22856 8676 22912 8678
rect 21956 8186 22012 8188
rect 22036 8186 22092 8188
rect 22116 8186 22172 8188
rect 22196 8186 22252 8188
rect 21956 8134 22002 8186
rect 22002 8134 22012 8186
rect 22036 8134 22066 8186
rect 22066 8134 22078 8186
rect 22078 8134 22092 8186
rect 22116 8134 22130 8186
rect 22130 8134 22142 8186
rect 22142 8134 22172 8186
rect 22196 8134 22206 8186
rect 22206 8134 22252 8186
rect 21956 8132 22012 8134
rect 22036 8132 22092 8134
rect 22116 8132 22172 8134
rect 22196 8132 22252 8134
rect 22616 7642 22672 7644
rect 22696 7642 22752 7644
rect 22776 7642 22832 7644
rect 22856 7642 22912 7644
rect 22616 7590 22662 7642
rect 22662 7590 22672 7642
rect 22696 7590 22726 7642
rect 22726 7590 22738 7642
rect 22738 7590 22752 7642
rect 22776 7590 22790 7642
rect 22790 7590 22802 7642
rect 22802 7590 22832 7642
rect 22856 7590 22866 7642
rect 22866 7590 22912 7642
rect 22616 7588 22672 7590
rect 22696 7588 22752 7590
rect 22776 7588 22832 7590
rect 22856 7588 22912 7590
rect 21956 7098 22012 7100
rect 22036 7098 22092 7100
rect 22116 7098 22172 7100
rect 22196 7098 22252 7100
rect 21956 7046 22002 7098
rect 22002 7046 22012 7098
rect 22036 7046 22066 7098
rect 22066 7046 22078 7098
rect 22078 7046 22092 7098
rect 22116 7046 22130 7098
rect 22130 7046 22142 7098
rect 22142 7046 22172 7098
rect 22196 7046 22206 7098
rect 22206 7046 22252 7098
rect 21956 7044 22012 7046
rect 22036 7044 22092 7046
rect 22116 7044 22172 7046
rect 22196 7044 22252 7046
rect 22616 6554 22672 6556
rect 22696 6554 22752 6556
rect 22776 6554 22832 6556
rect 22856 6554 22912 6556
rect 22616 6502 22662 6554
rect 22662 6502 22672 6554
rect 22696 6502 22726 6554
rect 22726 6502 22738 6554
rect 22738 6502 22752 6554
rect 22776 6502 22790 6554
rect 22790 6502 22802 6554
rect 22802 6502 22832 6554
rect 22856 6502 22866 6554
rect 22866 6502 22912 6554
rect 22616 6500 22672 6502
rect 22696 6500 22752 6502
rect 22776 6500 22832 6502
rect 22856 6500 22912 6502
rect 21956 6010 22012 6012
rect 22036 6010 22092 6012
rect 22116 6010 22172 6012
rect 22196 6010 22252 6012
rect 21956 5958 22002 6010
rect 22002 5958 22012 6010
rect 22036 5958 22066 6010
rect 22066 5958 22078 6010
rect 22078 5958 22092 6010
rect 22116 5958 22130 6010
rect 22130 5958 22142 6010
rect 22142 5958 22172 6010
rect 22196 5958 22206 6010
rect 22206 5958 22252 6010
rect 21956 5956 22012 5958
rect 22036 5956 22092 5958
rect 22116 5956 22172 5958
rect 22196 5956 22252 5958
rect 22616 5466 22672 5468
rect 22696 5466 22752 5468
rect 22776 5466 22832 5468
rect 22856 5466 22912 5468
rect 22616 5414 22662 5466
rect 22662 5414 22672 5466
rect 22696 5414 22726 5466
rect 22726 5414 22738 5466
rect 22738 5414 22752 5466
rect 22776 5414 22790 5466
rect 22790 5414 22802 5466
rect 22802 5414 22832 5466
rect 22856 5414 22866 5466
rect 22866 5414 22912 5466
rect 22616 5412 22672 5414
rect 22696 5412 22752 5414
rect 22776 5412 22832 5414
rect 22856 5412 22912 5414
rect 21956 4922 22012 4924
rect 22036 4922 22092 4924
rect 22116 4922 22172 4924
rect 22196 4922 22252 4924
rect 21956 4870 22002 4922
rect 22002 4870 22012 4922
rect 22036 4870 22066 4922
rect 22066 4870 22078 4922
rect 22078 4870 22092 4922
rect 22116 4870 22130 4922
rect 22130 4870 22142 4922
rect 22142 4870 22172 4922
rect 22196 4870 22206 4922
rect 22206 4870 22252 4922
rect 21956 4868 22012 4870
rect 22036 4868 22092 4870
rect 22116 4868 22172 4870
rect 22196 4868 22252 4870
rect 26956 61498 27012 61500
rect 27036 61498 27092 61500
rect 27116 61498 27172 61500
rect 27196 61498 27252 61500
rect 26956 61446 27002 61498
rect 27002 61446 27012 61498
rect 27036 61446 27066 61498
rect 27066 61446 27078 61498
rect 27078 61446 27092 61498
rect 27116 61446 27130 61498
rect 27130 61446 27142 61498
rect 27142 61446 27172 61498
rect 27196 61446 27206 61498
rect 27206 61446 27252 61498
rect 26956 61444 27012 61446
rect 27036 61444 27092 61446
rect 27116 61444 27172 61446
rect 27196 61444 27252 61446
rect 26956 60410 27012 60412
rect 27036 60410 27092 60412
rect 27116 60410 27172 60412
rect 27196 60410 27252 60412
rect 26956 60358 27002 60410
rect 27002 60358 27012 60410
rect 27036 60358 27066 60410
rect 27066 60358 27078 60410
rect 27078 60358 27092 60410
rect 27116 60358 27130 60410
rect 27130 60358 27142 60410
rect 27142 60358 27172 60410
rect 27196 60358 27206 60410
rect 27206 60358 27252 60410
rect 26956 60356 27012 60358
rect 27036 60356 27092 60358
rect 27116 60356 27172 60358
rect 27196 60356 27252 60358
rect 26956 59322 27012 59324
rect 27036 59322 27092 59324
rect 27116 59322 27172 59324
rect 27196 59322 27252 59324
rect 26956 59270 27002 59322
rect 27002 59270 27012 59322
rect 27036 59270 27066 59322
rect 27066 59270 27078 59322
rect 27078 59270 27092 59322
rect 27116 59270 27130 59322
rect 27130 59270 27142 59322
rect 27142 59270 27172 59322
rect 27196 59270 27206 59322
rect 27206 59270 27252 59322
rect 26956 59268 27012 59270
rect 27036 59268 27092 59270
rect 27116 59268 27172 59270
rect 27196 59268 27252 59270
rect 26956 58234 27012 58236
rect 27036 58234 27092 58236
rect 27116 58234 27172 58236
rect 27196 58234 27252 58236
rect 26956 58182 27002 58234
rect 27002 58182 27012 58234
rect 27036 58182 27066 58234
rect 27066 58182 27078 58234
rect 27078 58182 27092 58234
rect 27116 58182 27130 58234
rect 27130 58182 27142 58234
rect 27142 58182 27172 58234
rect 27196 58182 27206 58234
rect 27206 58182 27252 58234
rect 26956 58180 27012 58182
rect 27036 58180 27092 58182
rect 27116 58180 27172 58182
rect 27196 58180 27252 58182
rect 26956 57146 27012 57148
rect 27036 57146 27092 57148
rect 27116 57146 27172 57148
rect 27196 57146 27252 57148
rect 26956 57094 27002 57146
rect 27002 57094 27012 57146
rect 27036 57094 27066 57146
rect 27066 57094 27078 57146
rect 27078 57094 27092 57146
rect 27116 57094 27130 57146
rect 27130 57094 27142 57146
rect 27142 57094 27172 57146
rect 27196 57094 27206 57146
rect 27206 57094 27252 57146
rect 26956 57092 27012 57094
rect 27036 57092 27092 57094
rect 27116 57092 27172 57094
rect 27196 57092 27252 57094
rect 26956 56058 27012 56060
rect 27036 56058 27092 56060
rect 27116 56058 27172 56060
rect 27196 56058 27252 56060
rect 26956 56006 27002 56058
rect 27002 56006 27012 56058
rect 27036 56006 27066 56058
rect 27066 56006 27078 56058
rect 27078 56006 27092 56058
rect 27116 56006 27130 56058
rect 27130 56006 27142 56058
rect 27142 56006 27172 56058
rect 27196 56006 27206 56058
rect 27206 56006 27252 56058
rect 26956 56004 27012 56006
rect 27036 56004 27092 56006
rect 27116 56004 27172 56006
rect 27196 56004 27252 56006
rect 26956 54970 27012 54972
rect 27036 54970 27092 54972
rect 27116 54970 27172 54972
rect 27196 54970 27252 54972
rect 26956 54918 27002 54970
rect 27002 54918 27012 54970
rect 27036 54918 27066 54970
rect 27066 54918 27078 54970
rect 27078 54918 27092 54970
rect 27116 54918 27130 54970
rect 27130 54918 27142 54970
rect 27142 54918 27172 54970
rect 27196 54918 27206 54970
rect 27206 54918 27252 54970
rect 26956 54916 27012 54918
rect 27036 54916 27092 54918
rect 27116 54916 27172 54918
rect 27196 54916 27252 54918
rect 26956 53882 27012 53884
rect 27036 53882 27092 53884
rect 27116 53882 27172 53884
rect 27196 53882 27252 53884
rect 26956 53830 27002 53882
rect 27002 53830 27012 53882
rect 27036 53830 27066 53882
rect 27066 53830 27078 53882
rect 27078 53830 27092 53882
rect 27116 53830 27130 53882
rect 27130 53830 27142 53882
rect 27142 53830 27172 53882
rect 27196 53830 27206 53882
rect 27206 53830 27252 53882
rect 26956 53828 27012 53830
rect 27036 53828 27092 53830
rect 27116 53828 27172 53830
rect 27196 53828 27252 53830
rect 26956 52794 27012 52796
rect 27036 52794 27092 52796
rect 27116 52794 27172 52796
rect 27196 52794 27252 52796
rect 26956 52742 27002 52794
rect 27002 52742 27012 52794
rect 27036 52742 27066 52794
rect 27066 52742 27078 52794
rect 27078 52742 27092 52794
rect 27116 52742 27130 52794
rect 27130 52742 27142 52794
rect 27142 52742 27172 52794
rect 27196 52742 27206 52794
rect 27206 52742 27252 52794
rect 26956 52740 27012 52742
rect 27036 52740 27092 52742
rect 27116 52740 27172 52742
rect 27196 52740 27252 52742
rect 26956 51706 27012 51708
rect 27036 51706 27092 51708
rect 27116 51706 27172 51708
rect 27196 51706 27252 51708
rect 26956 51654 27002 51706
rect 27002 51654 27012 51706
rect 27036 51654 27066 51706
rect 27066 51654 27078 51706
rect 27078 51654 27092 51706
rect 27116 51654 27130 51706
rect 27130 51654 27142 51706
rect 27142 51654 27172 51706
rect 27196 51654 27206 51706
rect 27206 51654 27252 51706
rect 26956 51652 27012 51654
rect 27036 51652 27092 51654
rect 27116 51652 27172 51654
rect 27196 51652 27252 51654
rect 26956 50618 27012 50620
rect 27036 50618 27092 50620
rect 27116 50618 27172 50620
rect 27196 50618 27252 50620
rect 26956 50566 27002 50618
rect 27002 50566 27012 50618
rect 27036 50566 27066 50618
rect 27066 50566 27078 50618
rect 27078 50566 27092 50618
rect 27116 50566 27130 50618
rect 27130 50566 27142 50618
rect 27142 50566 27172 50618
rect 27196 50566 27206 50618
rect 27206 50566 27252 50618
rect 26956 50564 27012 50566
rect 27036 50564 27092 50566
rect 27116 50564 27172 50566
rect 27196 50564 27252 50566
rect 26956 49530 27012 49532
rect 27036 49530 27092 49532
rect 27116 49530 27172 49532
rect 27196 49530 27252 49532
rect 26956 49478 27002 49530
rect 27002 49478 27012 49530
rect 27036 49478 27066 49530
rect 27066 49478 27078 49530
rect 27078 49478 27092 49530
rect 27116 49478 27130 49530
rect 27130 49478 27142 49530
rect 27142 49478 27172 49530
rect 27196 49478 27206 49530
rect 27206 49478 27252 49530
rect 26956 49476 27012 49478
rect 27036 49476 27092 49478
rect 27116 49476 27172 49478
rect 27196 49476 27252 49478
rect 26956 48442 27012 48444
rect 27036 48442 27092 48444
rect 27116 48442 27172 48444
rect 27196 48442 27252 48444
rect 26956 48390 27002 48442
rect 27002 48390 27012 48442
rect 27036 48390 27066 48442
rect 27066 48390 27078 48442
rect 27078 48390 27092 48442
rect 27116 48390 27130 48442
rect 27130 48390 27142 48442
rect 27142 48390 27172 48442
rect 27196 48390 27206 48442
rect 27206 48390 27252 48442
rect 26956 48388 27012 48390
rect 27036 48388 27092 48390
rect 27116 48388 27172 48390
rect 27196 48388 27252 48390
rect 26956 47354 27012 47356
rect 27036 47354 27092 47356
rect 27116 47354 27172 47356
rect 27196 47354 27252 47356
rect 26956 47302 27002 47354
rect 27002 47302 27012 47354
rect 27036 47302 27066 47354
rect 27066 47302 27078 47354
rect 27078 47302 27092 47354
rect 27116 47302 27130 47354
rect 27130 47302 27142 47354
rect 27142 47302 27172 47354
rect 27196 47302 27206 47354
rect 27206 47302 27252 47354
rect 26956 47300 27012 47302
rect 27036 47300 27092 47302
rect 27116 47300 27172 47302
rect 27196 47300 27252 47302
rect 26956 46266 27012 46268
rect 27036 46266 27092 46268
rect 27116 46266 27172 46268
rect 27196 46266 27252 46268
rect 26956 46214 27002 46266
rect 27002 46214 27012 46266
rect 27036 46214 27066 46266
rect 27066 46214 27078 46266
rect 27078 46214 27092 46266
rect 27116 46214 27130 46266
rect 27130 46214 27142 46266
rect 27142 46214 27172 46266
rect 27196 46214 27206 46266
rect 27206 46214 27252 46266
rect 26956 46212 27012 46214
rect 27036 46212 27092 46214
rect 27116 46212 27172 46214
rect 27196 46212 27252 46214
rect 26956 45178 27012 45180
rect 27036 45178 27092 45180
rect 27116 45178 27172 45180
rect 27196 45178 27252 45180
rect 26956 45126 27002 45178
rect 27002 45126 27012 45178
rect 27036 45126 27066 45178
rect 27066 45126 27078 45178
rect 27078 45126 27092 45178
rect 27116 45126 27130 45178
rect 27130 45126 27142 45178
rect 27142 45126 27172 45178
rect 27196 45126 27206 45178
rect 27206 45126 27252 45178
rect 26956 45124 27012 45126
rect 27036 45124 27092 45126
rect 27116 45124 27172 45126
rect 27196 45124 27252 45126
rect 26956 44090 27012 44092
rect 27036 44090 27092 44092
rect 27116 44090 27172 44092
rect 27196 44090 27252 44092
rect 26956 44038 27002 44090
rect 27002 44038 27012 44090
rect 27036 44038 27066 44090
rect 27066 44038 27078 44090
rect 27078 44038 27092 44090
rect 27116 44038 27130 44090
rect 27130 44038 27142 44090
rect 27142 44038 27172 44090
rect 27196 44038 27206 44090
rect 27206 44038 27252 44090
rect 26956 44036 27012 44038
rect 27036 44036 27092 44038
rect 27116 44036 27172 44038
rect 27196 44036 27252 44038
rect 26956 43002 27012 43004
rect 27036 43002 27092 43004
rect 27116 43002 27172 43004
rect 27196 43002 27252 43004
rect 26956 42950 27002 43002
rect 27002 42950 27012 43002
rect 27036 42950 27066 43002
rect 27066 42950 27078 43002
rect 27078 42950 27092 43002
rect 27116 42950 27130 43002
rect 27130 42950 27142 43002
rect 27142 42950 27172 43002
rect 27196 42950 27206 43002
rect 27206 42950 27252 43002
rect 26956 42948 27012 42950
rect 27036 42948 27092 42950
rect 27116 42948 27172 42950
rect 27196 42948 27252 42950
rect 26956 41914 27012 41916
rect 27036 41914 27092 41916
rect 27116 41914 27172 41916
rect 27196 41914 27252 41916
rect 26956 41862 27002 41914
rect 27002 41862 27012 41914
rect 27036 41862 27066 41914
rect 27066 41862 27078 41914
rect 27078 41862 27092 41914
rect 27116 41862 27130 41914
rect 27130 41862 27142 41914
rect 27142 41862 27172 41914
rect 27196 41862 27206 41914
rect 27206 41862 27252 41914
rect 26956 41860 27012 41862
rect 27036 41860 27092 41862
rect 27116 41860 27172 41862
rect 27196 41860 27252 41862
rect 26956 40826 27012 40828
rect 27036 40826 27092 40828
rect 27116 40826 27172 40828
rect 27196 40826 27252 40828
rect 26956 40774 27002 40826
rect 27002 40774 27012 40826
rect 27036 40774 27066 40826
rect 27066 40774 27078 40826
rect 27078 40774 27092 40826
rect 27116 40774 27130 40826
rect 27130 40774 27142 40826
rect 27142 40774 27172 40826
rect 27196 40774 27206 40826
rect 27206 40774 27252 40826
rect 26956 40772 27012 40774
rect 27036 40772 27092 40774
rect 27116 40772 27172 40774
rect 27196 40772 27252 40774
rect 26956 39738 27012 39740
rect 27036 39738 27092 39740
rect 27116 39738 27172 39740
rect 27196 39738 27252 39740
rect 26956 39686 27002 39738
rect 27002 39686 27012 39738
rect 27036 39686 27066 39738
rect 27066 39686 27078 39738
rect 27078 39686 27092 39738
rect 27116 39686 27130 39738
rect 27130 39686 27142 39738
rect 27142 39686 27172 39738
rect 27196 39686 27206 39738
rect 27206 39686 27252 39738
rect 26956 39684 27012 39686
rect 27036 39684 27092 39686
rect 27116 39684 27172 39686
rect 27196 39684 27252 39686
rect 26956 38650 27012 38652
rect 27036 38650 27092 38652
rect 27116 38650 27172 38652
rect 27196 38650 27252 38652
rect 26956 38598 27002 38650
rect 27002 38598 27012 38650
rect 27036 38598 27066 38650
rect 27066 38598 27078 38650
rect 27078 38598 27092 38650
rect 27116 38598 27130 38650
rect 27130 38598 27142 38650
rect 27142 38598 27172 38650
rect 27196 38598 27206 38650
rect 27206 38598 27252 38650
rect 26956 38596 27012 38598
rect 27036 38596 27092 38598
rect 27116 38596 27172 38598
rect 27196 38596 27252 38598
rect 26956 37562 27012 37564
rect 27036 37562 27092 37564
rect 27116 37562 27172 37564
rect 27196 37562 27252 37564
rect 26956 37510 27002 37562
rect 27002 37510 27012 37562
rect 27036 37510 27066 37562
rect 27066 37510 27078 37562
rect 27078 37510 27092 37562
rect 27116 37510 27130 37562
rect 27130 37510 27142 37562
rect 27142 37510 27172 37562
rect 27196 37510 27206 37562
rect 27206 37510 27252 37562
rect 26956 37508 27012 37510
rect 27036 37508 27092 37510
rect 27116 37508 27172 37510
rect 27196 37508 27252 37510
rect 26956 36474 27012 36476
rect 27036 36474 27092 36476
rect 27116 36474 27172 36476
rect 27196 36474 27252 36476
rect 26956 36422 27002 36474
rect 27002 36422 27012 36474
rect 27036 36422 27066 36474
rect 27066 36422 27078 36474
rect 27078 36422 27092 36474
rect 27116 36422 27130 36474
rect 27130 36422 27142 36474
rect 27142 36422 27172 36474
rect 27196 36422 27206 36474
rect 27206 36422 27252 36474
rect 26956 36420 27012 36422
rect 27036 36420 27092 36422
rect 27116 36420 27172 36422
rect 27196 36420 27252 36422
rect 26956 35386 27012 35388
rect 27036 35386 27092 35388
rect 27116 35386 27172 35388
rect 27196 35386 27252 35388
rect 26956 35334 27002 35386
rect 27002 35334 27012 35386
rect 27036 35334 27066 35386
rect 27066 35334 27078 35386
rect 27078 35334 27092 35386
rect 27116 35334 27130 35386
rect 27130 35334 27142 35386
rect 27142 35334 27172 35386
rect 27196 35334 27206 35386
rect 27206 35334 27252 35386
rect 26956 35332 27012 35334
rect 27036 35332 27092 35334
rect 27116 35332 27172 35334
rect 27196 35332 27252 35334
rect 26956 34298 27012 34300
rect 27036 34298 27092 34300
rect 27116 34298 27172 34300
rect 27196 34298 27252 34300
rect 26956 34246 27002 34298
rect 27002 34246 27012 34298
rect 27036 34246 27066 34298
rect 27066 34246 27078 34298
rect 27078 34246 27092 34298
rect 27116 34246 27130 34298
rect 27130 34246 27142 34298
rect 27142 34246 27172 34298
rect 27196 34246 27206 34298
rect 27206 34246 27252 34298
rect 26956 34244 27012 34246
rect 27036 34244 27092 34246
rect 27116 34244 27172 34246
rect 27196 34244 27252 34246
rect 26956 33210 27012 33212
rect 27036 33210 27092 33212
rect 27116 33210 27172 33212
rect 27196 33210 27252 33212
rect 26956 33158 27002 33210
rect 27002 33158 27012 33210
rect 27036 33158 27066 33210
rect 27066 33158 27078 33210
rect 27078 33158 27092 33210
rect 27116 33158 27130 33210
rect 27130 33158 27142 33210
rect 27142 33158 27172 33210
rect 27196 33158 27206 33210
rect 27206 33158 27252 33210
rect 26956 33156 27012 33158
rect 27036 33156 27092 33158
rect 27116 33156 27172 33158
rect 27196 33156 27252 33158
rect 26956 32122 27012 32124
rect 27036 32122 27092 32124
rect 27116 32122 27172 32124
rect 27196 32122 27252 32124
rect 26956 32070 27002 32122
rect 27002 32070 27012 32122
rect 27036 32070 27066 32122
rect 27066 32070 27078 32122
rect 27078 32070 27092 32122
rect 27116 32070 27130 32122
rect 27130 32070 27142 32122
rect 27142 32070 27172 32122
rect 27196 32070 27206 32122
rect 27206 32070 27252 32122
rect 26956 32068 27012 32070
rect 27036 32068 27092 32070
rect 27116 32068 27172 32070
rect 27196 32068 27252 32070
rect 26956 31034 27012 31036
rect 27036 31034 27092 31036
rect 27116 31034 27172 31036
rect 27196 31034 27252 31036
rect 26956 30982 27002 31034
rect 27002 30982 27012 31034
rect 27036 30982 27066 31034
rect 27066 30982 27078 31034
rect 27078 30982 27092 31034
rect 27116 30982 27130 31034
rect 27130 30982 27142 31034
rect 27142 30982 27172 31034
rect 27196 30982 27206 31034
rect 27206 30982 27252 31034
rect 26956 30980 27012 30982
rect 27036 30980 27092 30982
rect 27116 30980 27172 30982
rect 27196 30980 27252 30982
rect 26956 29946 27012 29948
rect 27036 29946 27092 29948
rect 27116 29946 27172 29948
rect 27196 29946 27252 29948
rect 26956 29894 27002 29946
rect 27002 29894 27012 29946
rect 27036 29894 27066 29946
rect 27066 29894 27078 29946
rect 27078 29894 27092 29946
rect 27116 29894 27130 29946
rect 27130 29894 27142 29946
rect 27142 29894 27172 29946
rect 27196 29894 27206 29946
rect 27206 29894 27252 29946
rect 26956 29892 27012 29894
rect 27036 29892 27092 29894
rect 27116 29892 27172 29894
rect 27196 29892 27252 29894
rect 26956 28858 27012 28860
rect 27036 28858 27092 28860
rect 27116 28858 27172 28860
rect 27196 28858 27252 28860
rect 26956 28806 27002 28858
rect 27002 28806 27012 28858
rect 27036 28806 27066 28858
rect 27066 28806 27078 28858
rect 27078 28806 27092 28858
rect 27116 28806 27130 28858
rect 27130 28806 27142 28858
rect 27142 28806 27172 28858
rect 27196 28806 27206 28858
rect 27206 28806 27252 28858
rect 26956 28804 27012 28806
rect 27036 28804 27092 28806
rect 27116 28804 27172 28806
rect 27196 28804 27252 28806
rect 26956 27770 27012 27772
rect 27036 27770 27092 27772
rect 27116 27770 27172 27772
rect 27196 27770 27252 27772
rect 26956 27718 27002 27770
rect 27002 27718 27012 27770
rect 27036 27718 27066 27770
rect 27066 27718 27078 27770
rect 27078 27718 27092 27770
rect 27116 27718 27130 27770
rect 27130 27718 27142 27770
rect 27142 27718 27172 27770
rect 27196 27718 27206 27770
rect 27206 27718 27252 27770
rect 26956 27716 27012 27718
rect 27036 27716 27092 27718
rect 27116 27716 27172 27718
rect 27196 27716 27252 27718
rect 26956 26682 27012 26684
rect 27036 26682 27092 26684
rect 27116 26682 27172 26684
rect 27196 26682 27252 26684
rect 26956 26630 27002 26682
rect 27002 26630 27012 26682
rect 27036 26630 27066 26682
rect 27066 26630 27078 26682
rect 27078 26630 27092 26682
rect 27116 26630 27130 26682
rect 27130 26630 27142 26682
rect 27142 26630 27172 26682
rect 27196 26630 27206 26682
rect 27206 26630 27252 26682
rect 26956 26628 27012 26630
rect 27036 26628 27092 26630
rect 27116 26628 27172 26630
rect 27196 26628 27252 26630
rect 26956 25594 27012 25596
rect 27036 25594 27092 25596
rect 27116 25594 27172 25596
rect 27196 25594 27252 25596
rect 26956 25542 27002 25594
rect 27002 25542 27012 25594
rect 27036 25542 27066 25594
rect 27066 25542 27078 25594
rect 27078 25542 27092 25594
rect 27116 25542 27130 25594
rect 27130 25542 27142 25594
rect 27142 25542 27172 25594
rect 27196 25542 27206 25594
rect 27206 25542 27252 25594
rect 26956 25540 27012 25542
rect 27036 25540 27092 25542
rect 27116 25540 27172 25542
rect 27196 25540 27252 25542
rect 26956 24506 27012 24508
rect 27036 24506 27092 24508
rect 27116 24506 27172 24508
rect 27196 24506 27252 24508
rect 26956 24454 27002 24506
rect 27002 24454 27012 24506
rect 27036 24454 27066 24506
rect 27066 24454 27078 24506
rect 27078 24454 27092 24506
rect 27116 24454 27130 24506
rect 27130 24454 27142 24506
rect 27142 24454 27172 24506
rect 27196 24454 27206 24506
rect 27206 24454 27252 24506
rect 26956 24452 27012 24454
rect 27036 24452 27092 24454
rect 27116 24452 27172 24454
rect 27196 24452 27252 24454
rect 31956 69114 32012 69116
rect 32036 69114 32092 69116
rect 32116 69114 32172 69116
rect 32196 69114 32252 69116
rect 31956 69062 32002 69114
rect 32002 69062 32012 69114
rect 32036 69062 32066 69114
rect 32066 69062 32078 69114
rect 32078 69062 32092 69114
rect 32116 69062 32130 69114
rect 32130 69062 32142 69114
rect 32142 69062 32172 69114
rect 32196 69062 32206 69114
rect 32206 69062 32252 69114
rect 31956 69060 32012 69062
rect 32036 69060 32092 69062
rect 32116 69060 32172 69062
rect 32196 69060 32252 69062
rect 27616 68570 27672 68572
rect 27696 68570 27752 68572
rect 27776 68570 27832 68572
rect 27856 68570 27912 68572
rect 27616 68518 27662 68570
rect 27662 68518 27672 68570
rect 27696 68518 27726 68570
rect 27726 68518 27738 68570
rect 27738 68518 27752 68570
rect 27776 68518 27790 68570
rect 27790 68518 27802 68570
rect 27802 68518 27832 68570
rect 27856 68518 27866 68570
rect 27866 68518 27912 68570
rect 27616 68516 27672 68518
rect 27696 68516 27752 68518
rect 27776 68516 27832 68518
rect 27856 68516 27912 68518
rect 32616 68570 32672 68572
rect 32696 68570 32752 68572
rect 32776 68570 32832 68572
rect 32856 68570 32912 68572
rect 32616 68518 32662 68570
rect 32662 68518 32672 68570
rect 32696 68518 32726 68570
rect 32726 68518 32738 68570
rect 32738 68518 32752 68570
rect 32776 68518 32790 68570
rect 32790 68518 32802 68570
rect 32802 68518 32832 68570
rect 32856 68518 32866 68570
rect 32866 68518 32912 68570
rect 32616 68516 32672 68518
rect 32696 68516 32752 68518
rect 32776 68516 32832 68518
rect 32856 68516 32912 68518
rect 27616 67482 27672 67484
rect 27696 67482 27752 67484
rect 27776 67482 27832 67484
rect 27856 67482 27912 67484
rect 27616 67430 27662 67482
rect 27662 67430 27672 67482
rect 27696 67430 27726 67482
rect 27726 67430 27738 67482
rect 27738 67430 27752 67482
rect 27776 67430 27790 67482
rect 27790 67430 27802 67482
rect 27802 67430 27832 67482
rect 27856 67430 27866 67482
rect 27866 67430 27912 67482
rect 27616 67428 27672 67430
rect 27696 67428 27752 67430
rect 27776 67428 27832 67430
rect 27856 67428 27912 67430
rect 27616 66394 27672 66396
rect 27696 66394 27752 66396
rect 27776 66394 27832 66396
rect 27856 66394 27912 66396
rect 27616 66342 27662 66394
rect 27662 66342 27672 66394
rect 27696 66342 27726 66394
rect 27726 66342 27738 66394
rect 27738 66342 27752 66394
rect 27776 66342 27790 66394
rect 27790 66342 27802 66394
rect 27802 66342 27832 66394
rect 27856 66342 27866 66394
rect 27866 66342 27912 66394
rect 27616 66340 27672 66342
rect 27696 66340 27752 66342
rect 27776 66340 27832 66342
rect 27856 66340 27912 66342
rect 27616 65306 27672 65308
rect 27696 65306 27752 65308
rect 27776 65306 27832 65308
rect 27856 65306 27912 65308
rect 27616 65254 27662 65306
rect 27662 65254 27672 65306
rect 27696 65254 27726 65306
rect 27726 65254 27738 65306
rect 27738 65254 27752 65306
rect 27776 65254 27790 65306
rect 27790 65254 27802 65306
rect 27802 65254 27832 65306
rect 27856 65254 27866 65306
rect 27866 65254 27912 65306
rect 27616 65252 27672 65254
rect 27696 65252 27752 65254
rect 27776 65252 27832 65254
rect 27856 65252 27912 65254
rect 27616 64218 27672 64220
rect 27696 64218 27752 64220
rect 27776 64218 27832 64220
rect 27856 64218 27912 64220
rect 27616 64166 27662 64218
rect 27662 64166 27672 64218
rect 27696 64166 27726 64218
rect 27726 64166 27738 64218
rect 27738 64166 27752 64218
rect 27776 64166 27790 64218
rect 27790 64166 27802 64218
rect 27802 64166 27832 64218
rect 27856 64166 27866 64218
rect 27866 64166 27912 64218
rect 27616 64164 27672 64166
rect 27696 64164 27752 64166
rect 27776 64164 27832 64166
rect 27856 64164 27912 64166
rect 27616 63130 27672 63132
rect 27696 63130 27752 63132
rect 27776 63130 27832 63132
rect 27856 63130 27912 63132
rect 27616 63078 27662 63130
rect 27662 63078 27672 63130
rect 27696 63078 27726 63130
rect 27726 63078 27738 63130
rect 27738 63078 27752 63130
rect 27776 63078 27790 63130
rect 27790 63078 27802 63130
rect 27802 63078 27832 63130
rect 27856 63078 27866 63130
rect 27866 63078 27912 63130
rect 27616 63076 27672 63078
rect 27696 63076 27752 63078
rect 27776 63076 27832 63078
rect 27856 63076 27912 63078
rect 27616 62042 27672 62044
rect 27696 62042 27752 62044
rect 27776 62042 27832 62044
rect 27856 62042 27912 62044
rect 27616 61990 27662 62042
rect 27662 61990 27672 62042
rect 27696 61990 27726 62042
rect 27726 61990 27738 62042
rect 27738 61990 27752 62042
rect 27776 61990 27790 62042
rect 27790 61990 27802 62042
rect 27802 61990 27832 62042
rect 27856 61990 27866 62042
rect 27866 61990 27912 62042
rect 27616 61988 27672 61990
rect 27696 61988 27752 61990
rect 27776 61988 27832 61990
rect 27856 61988 27912 61990
rect 27616 60954 27672 60956
rect 27696 60954 27752 60956
rect 27776 60954 27832 60956
rect 27856 60954 27912 60956
rect 27616 60902 27662 60954
rect 27662 60902 27672 60954
rect 27696 60902 27726 60954
rect 27726 60902 27738 60954
rect 27738 60902 27752 60954
rect 27776 60902 27790 60954
rect 27790 60902 27802 60954
rect 27802 60902 27832 60954
rect 27856 60902 27866 60954
rect 27866 60902 27912 60954
rect 27616 60900 27672 60902
rect 27696 60900 27752 60902
rect 27776 60900 27832 60902
rect 27856 60900 27912 60902
rect 27616 59866 27672 59868
rect 27696 59866 27752 59868
rect 27776 59866 27832 59868
rect 27856 59866 27912 59868
rect 27616 59814 27662 59866
rect 27662 59814 27672 59866
rect 27696 59814 27726 59866
rect 27726 59814 27738 59866
rect 27738 59814 27752 59866
rect 27776 59814 27790 59866
rect 27790 59814 27802 59866
rect 27802 59814 27832 59866
rect 27856 59814 27866 59866
rect 27866 59814 27912 59866
rect 27616 59812 27672 59814
rect 27696 59812 27752 59814
rect 27776 59812 27832 59814
rect 27856 59812 27912 59814
rect 27616 58778 27672 58780
rect 27696 58778 27752 58780
rect 27776 58778 27832 58780
rect 27856 58778 27912 58780
rect 27616 58726 27662 58778
rect 27662 58726 27672 58778
rect 27696 58726 27726 58778
rect 27726 58726 27738 58778
rect 27738 58726 27752 58778
rect 27776 58726 27790 58778
rect 27790 58726 27802 58778
rect 27802 58726 27832 58778
rect 27856 58726 27866 58778
rect 27866 58726 27912 58778
rect 27616 58724 27672 58726
rect 27696 58724 27752 58726
rect 27776 58724 27832 58726
rect 27856 58724 27912 58726
rect 27616 57690 27672 57692
rect 27696 57690 27752 57692
rect 27776 57690 27832 57692
rect 27856 57690 27912 57692
rect 27616 57638 27662 57690
rect 27662 57638 27672 57690
rect 27696 57638 27726 57690
rect 27726 57638 27738 57690
rect 27738 57638 27752 57690
rect 27776 57638 27790 57690
rect 27790 57638 27802 57690
rect 27802 57638 27832 57690
rect 27856 57638 27866 57690
rect 27866 57638 27912 57690
rect 27616 57636 27672 57638
rect 27696 57636 27752 57638
rect 27776 57636 27832 57638
rect 27856 57636 27912 57638
rect 27616 56602 27672 56604
rect 27696 56602 27752 56604
rect 27776 56602 27832 56604
rect 27856 56602 27912 56604
rect 27616 56550 27662 56602
rect 27662 56550 27672 56602
rect 27696 56550 27726 56602
rect 27726 56550 27738 56602
rect 27738 56550 27752 56602
rect 27776 56550 27790 56602
rect 27790 56550 27802 56602
rect 27802 56550 27832 56602
rect 27856 56550 27866 56602
rect 27866 56550 27912 56602
rect 27616 56548 27672 56550
rect 27696 56548 27752 56550
rect 27776 56548 27832 56550
rect 27856 56548 27912 56550
rect 27616 55514 27672 55516
rect 27696 55514 27752 55516
rect 27776 55514 27832 55516
rect 27856 55514 27912 55516
rect 27616 55462 27662 55514
rect 27662 55462 27672 55514
rect 27696 55462 27726 55514
rect 27726 55462 27738 55514
rect 27738 55462 27752 55514
rect 27776 55462 27790 55514
rect 27790 55462 27802 55514
rect 27802 55462 27832 55514
rect 27856 55462 27866 55514
rect 27866 55462 27912 55514
rect 27616 55460 27672 55462
rect 27696 55460 27752 55462
rect 27776 55460 27832 55462
rect 27856 55460 27912 55462
rect 27616 54426 27672 54428
rect 27696 54426 27752 54428
rect 27776 54426 27832 54428
rect 27856 54426 27912 54428
rect 27616 54374 27662 54426
rect 27662 54374 27672 54426
rect 27696 54374 27726 54426
rect 27726 54374 27738 54426
rect 27738 54374 27752 54426
rect 27776 54374 27790 54426
rect 27790 54374 27802 54426
rect 27802 54374 27832 54426
rect 27856 54374 27866 54426
rect 27866 54374 27912 54426
rect 27616 54372 27672 54374
rect 27696 54372 27752 54374
rect 27776 54372 27832 54374
rect 27856 54372 27912 54374
rect 27616 53338 27672 53340
rect 27696 53338 27752 53340
rect 27776 53338 27832 53340
rect 27856 53338 27912 53340
rect 27616 53286 27662 53338
rect 27662 53286 27672 53338
rect 27696 53286 27726 53338
rect 27726 53286 27738 53338
rect 27738 53286 27752 53338
rect 27776 53286 27790 53338
rect 27790 53286 27802 53338
rect 27802 53286 27832 53338
rect 27856 53286 27866 53338
rect 27866 53286 27912 53338
rect 27616 53284 27672 53286
rect 27696 53284 27752 53286
rect 27776 53284 27832 53286
rect 27856 53284 27912 53286
rect 27616 52250 27672 52252
rect 27696 52250 27752 52252
rect 27776 52250 27832 52252
rect 27856 52250 27912 52252
rect 27616 52198 27662 52250
rect 27662 52198 27672 52250
rect 27696 52198 27726 52250
rect 27726 52198 27738 52250
rect 27738 52198 27752 52250
rect 27776 52198 27790 52250
rect 27790 52198 27802 52250
rect 27802 52198 27832 52250
rect 27856 52198 27866 52250
rect 27866 52198 27912 52250
rect 27616 52196 27672 52198
rect 27696 52196 27752 52198
rect 27776 52196 27832 52198
rect 27856 52196 27912 52198
rect 27616 51162 27672 51164
rect 27696 51162 27752 51164
rect 27776 51162 27832 51164
rect 27856 51162 27912 51164
rect 27616 51110 27662 51162
rect 27662 51110 27672 51162
rect 27696 51110 27726 51162
rect 27726 51110 27738 51162
rect 27738 51110 27752 51162
rect 27776 51110 27790 51162
rect 27790 51110 27802 51162
rect 27802 51110 27832 51162
rect 27856 51110 27866 51162
rect 27866 51110 27912 51162
rect 27616 51108 27672 51110
rect 27696 51108 27752 51110
rect 27776 51108 27832 51110
rect 27856 51108 27912 51110
rect 27616 50074 27672 50076
rect 27696 50074 27752 50076
rect 27776 50074 27832 50076
rect 27856 50074 27912 50076
rect 27616 50022 27662 50074
rect 27662 50022 27672 50074
rect 27696 50022 27726 50074
rect 27726 50022 27738 50074
rect 27738 50022 27752 50074
rect 27776 50022 27790 50074
rect 27790 50022 27802 50074
rect 27802 50022 27832 50074
rect 27856 50022 27866 50074
rect 27866 50022 27912 50074
rect 27616 50020 27672 50022
rect 27696 50020 27752 50022
rect 27776 50020 27832 50022
rect 27856 50020 27912 50022
rect 27616 48986 27672 48988
rect 27696 48986 27752 48988
rect 27776 48986 27832 48988
rect 27856 48986 27912 48988
rect 27616 48934 27662 48986
rect 27662 48934 27672 48986
rect 27696 48934 27726 48986
rect 27726 48934 27738 48986
rect 27738 48934 27752 48986
rect 27776 48934 27790 48986
rect 27790 48934 27802 48986
rect 27802 48934 27832 48986
rect 27856 48934 27866 48986
rect 27866 48934 27912 48986
rect 27616 48932 27672 48934
rect 27696 48932 27752 48934
rect 27776 48932 27832 48934
rect 27856 48932 27912 48934
rect 27616 47898 27672 47900
rect 27696 47898 27752 47900
rect 27776 47898 27832 47900
rect 27856 47898 27912 47900
rect 27616 47846 27662 47898
rect 27662 47846 27672 47898
rect 27696 47846 27726 47898
rect 27726 47846 27738 47898
rect 27738 47846 27752 47898
rect 27776 47846 27790 47898
rect 27790 47846 27802 47898
rect 27802 47846 27832 47898
rect 27856 47846 27866 47898
rect 27866 47846 27912 47898
rect 27616 47844 27672 47846
rect 27696 47844 27752 47846
rect 27776 47844 27832 47846
rect 27856 47844 27912 47846
rect 27616 46810 27672 46812
rect 27696 46810 27752 46812
rect 27776 46810 27832 46812
rect 27856 46810 27912 46812
rect 27616 46758 27662 46810
rect 27662 46758 27672 46810
rect 27696 46758 27726 46810
rect 27726 46758 27738 46810
rect 27738 46758 27752 46810
rect 27776 46758 27790 46810
rect 27790 46758 27802 46810
rect 27802 46758 27832 46810
rect 27856 46758 27866 46810
rect 27866 46758 27912 46810
rect 27616 46756 27672 46758
rect 27696 46756 27752 46758
rect 27776 46756 27832 46758
rect 27856 46756 27912 46758
rect 27616 45722 27672 45724
rect 27696 45722 27752 45724
rect 27776 45722 27832 45724
rect 27856 45722 27912 45724
rect 27616 45670 27662 45722
rect 27662 45670 27672 45722
rect 27696 45670 27726 45722
rect 27726 45670 27738 45722
rect 27738 45670 27752 45722
rect 27776 45670 27790 45722
rect 27790 45670 27802 45722
rect 27802 45670 27832 45722
rect 27856 45670 27866 45722
rect 27866 45670 27912 45722
rect 27616 45668 27672 45670
rect 27696 45668 27752 45670
rect 27776 45668 27832 45670
rect 27856 45668 27912 45670
rect 27616 44634 27672 44636
rect 27696 44634 27752 44636
rect 27776 44634 27832 44636
rect 27856 44634 27912 44636
rect 27616 44582 27662 44634
rect 27662 44582 27672 44634
rect 27696 44582 27726 44634
rect 27726 44582 27738 44634
rect 27738 44582 27752 44634
rect 27776 44582 27790 44634
rect 27790 44582 27802 44634
rect 27802 44582 27832 44634
rect 27856 44582 27866 44634
rect 27866 44582 27912 44634
rect 27616 44580 27672 44582
rect 27696 44580 27752 44582
rect 27776 44580 27832 44582
rect 27856 44580 27912 44582
rect 27616 43546 27672 43548
rect 27696 43546 27752 43548
rect 27776 43546 27832 43548
rect 27856 43546 27912 43548
rect 27616 43494 27662 43546
rect 27662 43494 27672 43546
rect 27696 43494 27726 43546
rect 27726 43494 27738 43546
rect 27738 43494 27752 43546
rect 27776 43494 27790 43546
rect 27790 43494 27802 43546
rect 27802 43494 27832 43546
rect 27856 43494 27866 43546
rect 27866 43494 27912 43546
rect 27616 43492 27672 43494
rect 27696 43492 27752 43494
rect 27776 43492 27832 43494
rect 27856 43492 27912 43494
rect 27616 42458 27672 42460
rect 27696 42458 27752 42460
rect 27776 42458 27832 42460
rect 27856 42458 27912 42460
rect 27616 42406 27662 42458
rect 27662 42406 27672 42458
rect 27696 42406 27726 42458
rect 27726 42406 27738 42458
rect 27738 42406 27752 42458
rect 27776 42406 27790 42458
rect 27790 42406 27802 42458
rect 27802 42406 27832 42458
rect 27856 42406 27866 42458
rect 27866 42406 27912 42458
rect 27616 42404 27672 42406
rect 27696 42404 27752 42406
rect 27776 42404 27832 42406
rect 27856 42404 27912 42406
rect 27616 41370 27672 41372
rect 27696 41370 27752 41372
rect 27776 41370 27832 41372
rect 27856 41370 27912 41372
rect 27616 41318 27662 41370
rect 27662 41318 27672 41370
rect 27696 41318 27726 41370
rect 27726 41318 27738 41370
rect 27738 41318 27752 41370
rect 27776 41318 27790 41370
rect 27790 41318 27802 41370
rect 27802 41318 27832 41370
rect 27856 41318 27866 41370
rect 27866 41318 27912 41370
rect 27616 41316 27672 41318
rect 27696 41316 27752 41318
rect 27776 41316 27832 41318
rect 27856 41316 27912 41318
rect 27616 40282 27672 40284
rect 27696 40282 27752 40284
rect 27776 40282 27832 40284
rect 27856 40282 27912 40284
rect 27616 40230 27662 40282
rect 27662 40230 27672 40282
rect 27696 40230 27726 40282
rect 27726 40230 27738 40282
rect 27738 40230 27752 40282
rect 27776 40230 27790 40282
rect 27790 40230 27802 40282
rect 27802 40230 27832 40282
rect 27856 40230 27866 40282
rect 27866 40230 27912 40282
rect 27616 40228 27672 40230
rect 27696 40228 27752 40230
rect 27776 40228 27832 40230
rect 27856 40228 27912 40230
rect 27616 39194 27672 39196
rect 27696 39194 27752 39196
rect 27776 39194 27832 39196
rect 27856 39194 27912 39196
rect 27616 39142 27662 39194
rect 27662 39142 27672 39194
rect 27696 39142 27726 39194
rect 27726 39142 27738 39194
rect 27738 39142 27752 39194
rect 27776 39142 27790 39194
rect 27790 39142 27802 39194
rect 27802 39142 27832 39194
rect 27856 39142 27866 39194
rect 27866 39142 27912 39194
rect 27616 39140 27672 39142
rect 27696 39140 27752 39142
rect 27776 39140 27832 39142
rect 27856 39140 27912 39142
rect 27616 38106 27672 38108
rect 27696 38106 27752 38108
rect 27776 38106 27832 38108
rect 27856 38106 27912 38108
rect 27616 38054 27662 38106
rect 27662 38054 27672 38106
rect 27696 38054 27726 38106
rect 27726 38054 27738 38106
rect 27738 38054 27752 38106
rect 27776 38054 27790 38106
rect 27790 38054 27802 38106
rect 27802 38054 27832 38106
rect 27856 38054 27866 38106
rect 27866 38054 27912 38106
rect 27616 38052 27672 38054
rect 27696 38052 27752 38054
rect 27776 38052 27832 38054
rect 27856 38052 27912 38054
rect 27616 37018 27672 37020
rect 27696 37018 27752 37020
rect 27776 37018 27832 37020
rect 27856 37018 27912 37020
rect 27616 36966 27662 37018
rect 27662 36966 27672 37018
rect 27696 36966 27726 37018
rect 27726 36966 27738 37018
rect 27738 36966 27752 37018
rect 27776 36966 27790 37018
rect 27790 36966 27802 37018
rect 27802 36966 27832 37018
rect 27856 36966 27866 37018
rect 27866 36966 27912 37018
rect 27616 36964 27672 36966
rect 27696 36964 27752 36966
rect 27776 36964 27832 36966
rect 27856 36964 27912 36966
rect 27616 35930 27672 35932
rect 27696 35930 27752 35932
rect 27776 35930 27832 35932
rect 27856 35930 27912 35932
rect 27616 35878 27662 35930
rect 27662 35878 27672 35930
rect 27696 35878 27726 35930
rect 27726 35878 27738 35930
rect 27738 35878 27752 35930
rect 27776 35878 27790 35930
rect 27790 35878 27802 35930
rect 27802 35878 27832 35930
rect 27856 35878 27866 35930
rect 27866 35878 27912 35930
rect 27616 35876 27672 35878
rect 27696 35876 27752 35878
rect 27776 35876 27832 35878
rect 27856 35876 27912 35878
rect 27616 34842 27672 34844
rect 27696 34842 27752 34844
rect 27776 34842 27832 34844
rect 27856 34842 27912 34844
rect 27616 34790 27662 34842
rect 27662 34790 27672 34842
rect 27696 34790 27726 34842
rect 27726 34790 27738 34842
rect 27738 34790 27752 34842
rect 27776 34790 27790 34842
rect 27790 34790 27802 34842
rect 27802 34790 27832 34842
rect 27856 34790 27866 34842
rect 27866 34790 27912 34842
rect 27616 34788 27672 34790
rect 27696 34788 27752 34790
rect 27776 34788 27832 34790
rect 27856 34788 27912 34790
rect 27616 33754 27672 33756
rect 27696 33754 27752 33756
rect 27776 33754 27832 33756
rect 27856 33754 27912 33756
rect 27616 33702 27662 33754
rect 27662 33702 27672 33754
rect 27696 33702 27726 33754
rect 27726 33702 27738 33754
rect 27738 33702 27752 33754
rect 27776 33702 27790 33754
rect 27790 33702 27802 33754
rect 27802 33702 27832 33754
rect 27856 33702 27866 33754
rect 27866 33702 27912 33754
rect 27616 33700 27672 33702
rect 27696 33700 27752 33702
rect 27776 33700 27832 33702
rect 27856 33700 27912 33702
rect 27616 32666 27672 32668
rect 27696 32666 27752 32668
rect 27776 32666 27832 32668
rect 27856 32666 27912 32668
rect 27616 32614 27662 32666
rect 27662 32614 27672 32666
rect 27696 32614 27726 32666
rect 27726 32614 27738 32666
rect 27738 32614 27752 32666
rect 27776 32614 27790 32666
rect 27790 32614 27802 32666
rect 27802 32614 27832 32666
rect 27856 32614 27866 32666
rect 27866 32614 27912 32666
rect 27616 32612 27672 32614
rect 27696 32612 27752 32614
rect 27776 32612 27832 32614
rect 27856 32612 27912 32614
rect 27616 31578 27672 31580
rect 27696 31578 27752 31580
rect 27776 31578 27832 31580
rect 27856 31578 27912 31580
rect 27616 31526 27662 31578
rect 27662 31526 27672 31578
rect 27696 31526 27726 31578
rect 27726 31526 27738 31578
rect 27738 31526 27752 31578
rect 27776 31526 27790 31578
rect 27790 31526 27802 31578
rect 27802 31526 27832 31578
rect 27856 31526 27866 31578
rect 27866 31526 27912 31578
rect 27616 31524 27672 31526
rect 27696 31524 27752 31526
rect 27776 31524 27832 31526
rect 27856 31524 27912 31526
rect 27616 30490 27672 30492
rect 27696 30490 27752 30492
rect 27776 30490 27832 30492
rect 27856 30490 27912 30492
rect 27616 30438 27662 30490
rect 27662 30438 27672 30490
rect 27696 30438 27726 30490
rect 27726 30438 27738 30490
rect 27738 30438 27752 30490
rect 27776 30438 27790 30490
rect 27790 30438 27802 30490
rect 27802 30438 27832 30490
rect 27856 30438 27866 30490
rect 27866 30438 27912 30490
rect 27616 30436 27672 30438
rect 27696 30436 27752 30438
rect 27776 30436 27832 30438
rect 27856 30436 27912 30438
rect 28814 45872 28870 45928
rect 27616 29402 27672 29404
rect 27696 29402 27752 29404
rect 27776 29402 27832 29404
rect 27856 29402 27912 29404
rect 27616 29350 27662 29402
rect 27662 29350 27672 29402
rect 27696 29350 27726 29402
rect 27726 29350 27738 29402
rect 27738 29350 27752 29402
rect 27776 29350 27790 29402
rect 27790 29350 27802 29402
rect 27802 29350 27832 29402
rect 27856 29350 27866 29402
rect 27866 29350 27912 29402
rect 27616 29348 27672 29350
rect 27696 29348 27752 29350
rect 27776 29348 27832 29350
rect 27856 29348 27912 29350
rect 27616 28314 27672 28316
rect 27696 28314 27752 28316
rect 27776 28314 27832 28316
rect 27856 28314 27912 28316
rect 27616 28262 27662 28314
rect 27662 28262 27672 28314
rect 27696 28262 27726 28314
rect 27726 28262 27738 28314
rect 27738 28262 27752 28314
rect 27776 28262 27790 28314
rect 27790 28262 27802 28314
rect 27802 28262 27832 28314
rect 27856 28262 27866 28314
rect 27866 28262 27912 28314
rect 27616 28260 27672 28262
rect 27696 28260 27752 28262
rect 27776 28260 27832 28262
rect 27856 28260 27912 28262
rect 27616 27226 27672 27228
rect 27696 27226 27752 27228
rect 27776 27226 27832 27228
rect 27856 27226 27912 27228
rect 27616 27174 27662 27226
rect 27662 27174 27672 27226
rect 27696 27174 27726 27226
rect 27726 27174 27738 27226
rect 27738 27174 27752 27226
rect 27776 27174 27790 27226
rect 27790 27174 27802 27226
rect 27802 27174 27832 27226
rect 27856 27174 27866 27226
rect 27866 27174 27912 27226
rect 27616 27172 27672 27174
rect 27696 27172 27752 27174
rect 27776 27172 27832 27174
rect 27856 27172 27912 27174
rect 27616 26138 27672 26140
rect 27696 26138 27752 26140
rect 27776 26138 27832 26140
rect 27856 26138 27912 26140
rect 27616 26086 27662 26138
rect 27662 26086 27672 26138
rect 27696 26086 27726 26138
rect 27726 26086 27738 26138
rect 27738 26086 27752 26138
rect 27776 26086 27790 26138
rect 27790 26086 27802 26138
rect 27802 26086 27832 26138
rect 27856 26086 27866 26138
rect 27866 26086 27912 26138
rect 27616 26084 27672 26086
rect 27696 26084 27752 26086
rect 27776 26084 27832 26086
rect 27856 26084 27912 26086
rect 27616 25050 27672 25052
rect 27696 25050 27752 25052
rect 27776 25050 27832 25052
rect 27856 25050 27912 25052
rect 27616 24998 27662 25050
rect 27662 24998 27672 25050
rect 27696 24998 27726 25050
rect 27726 24998 27738 25050
rect 27738 24998 27752 25050
rect 27776 24998 27790 25050
rect 27790 24998 27802 25050
rect 27802 24998 27832 25050
rect 27856 24998 27866 25050
rect 27866 24998 27912 25050
rect 27616 24996 27672 24998
rect 27696 24996 27752 24998
rect 27776 24996 27832 24998
rect 27856 24996 27912 24998
rect 27616 23962 27672 23964
rect 27696 23962 27752 23964
rect 27776 23962 27832 23964
rect 27856 23962 27912 23964
rect 27616 23910 27662 23962
rect 27662 23910 27672 23962
rect 27696 23910 27726 23962
rect 27726 23910 27738 23962
rect 27738 23910 27752 23962
rect 27776 23910 27790 23962
rect 27790 23910 27802 23962
rect 27802 23910 27832 23962
rect 27856 23910 27866 23962
rect 27866 23910 27912 23962
rect 27616 23908 27672 23910
rect 27696 23908 27752 23910
rect 27776 23908 27832 23910
rect 27856 23908 27912 23910
rect 26956 23418 27012 23420
rect 27036 23418 27092 23420
rect 27116 23418 27172 23420
rect 27196 23418 27252 23420
rect 26956 23366 27002 23418
rect 27002 23366 27012 23418
rect 27036 23366 27066 23418
rect 27066 23366 27078 23418
rect 27078 23366 27092 23418
rect 27116 23366 27130 23418
rect 27130 23366 27142 23418
rect 27142 23366 27172 23418
rect 27196 23366 27206 23418
rect 27206 23366 27252 23418
rect 26956 23364 27012 23366
rect 27036 23364 27092 23366
rect 27116 23364 27172 23366
rect 27196 23364 27252 23366
rect 27616 22874 27672 22876
rect 27696 22874 27752 22876
rect 27776 22874 27832 22876
rect 27856 22874 27912 22876
rect 27616 22822 27662 22874
rect 27662 22822 27672 22874
rect 27696 22822 27726 22874
rect 27726 22822 27738 22874
rect 27738 22822 27752 22874
rect 27776 22822 27790 22874
rect 27790 22822 27802 22874
rect 27802 22822 27832 22874
rect 27856 22822 27866 22874
rect 27866 22822 27912 22874
rect 27616 22820 27672 22822
rect 27696 22820 27752 22822
rect 27776 22820 27832 22822
rect 27856 22820 27912 22822
rect 26956 22330 27012 22332
rect 27036 22330 27092 22332
rect 27116 22330 27172 22332
rect 27196 22330 27252 22332
rect 26956 22278 27002 22330
rect 27002 22278 27012 22330
rect 27036 22278 27066 22330
rect 27066 22278 27078 22330
rect 27078 22278 27092 22330
rect 27116 22278 27130 22330
rect 27130 22278 27142 22330
rect 27142 22278 27172 22330
rect 27196 22278 27206 22330
rect 27206 22278 27252 22330
rect 26956 22276 27012 22278
rect 27036 22276 27092 22278
rect 27116 22276 27172 22278
rect 27196 22276 27252 22278
rect 27616 21786 27672 21788
rect 27696 21786 27752 21788
rect 27776 21786 27832 21788
rect 27856 21786 27912 21788
rect 27616 21734 27662 21786
rect 27662 21734 27672 21786
rect 27696 21734 27726 21786
rect 27726 21734 27738 21786
rect 27738 21734 27752 21786
rect 27776 21734 27790 21786
rect 27790 21734 27802 21786
rect 27802 21734 27832 21786
rect 27856 21734 27866 21786
rect 27866 21734 27912 21786
rect 27616 21732 27672 21734
rect 27696 21732 27752 21734
rect 27776 21732 27832 21734
rect 27856 21732 27912 21734
rect 26956 21242 27012 21244
rect 27036 21242 27092 21244
rect 27116 21242 27172 21244
rect 27196 21242 27252 21244
rect 26956 21190 27002 21242
rect 27002 21190 27012 21242
rect 27036 21190 27066 21242
rect 27066 21190 27078 21242
rect 27078 21190 27092 21242
rect 27116 21190 27130 21242
rect 27130 21190 27142 21242
rect 27142 21190 27172 21242
rect 27196 21190 27206 21242
rect 27206 21190 27252 21242
rect 26956 21188 27012 21190
rect 27036 21188 27092 21190
rect 27116 21188 27172 21190
rect 27196 21188 27252 21190
rect 26956 20154 27012 20156
rect 27036 20154 27092 20156
rect 27116 20154 27172 20156
rect 27196 20154 27252 20156
rect 26956 20102 27002 20154
rect 27002 20102 27012 20154
rect 27036 20102 27066 20154
rect 27066 20102 27078 20154
rect 27078 20102 27092 20154
rect 27116 20102 27130 20154
rect 27130 20102 27142 20154
rect 27142 20102 27172 20154
rect 27196 20102 27206 20154
rect 27206 20102 27252 20154
rect 26956 20100 27012 20102
rect 27036 20100 27092 20102
rect 27116 20100 27172 20102
rect 27196 20100 27252 20102
rect 26956 19066 27012 19068
rect 27036 19066 27092 19068
rect 27116 19066 27172 19068
rect 27196 19066 27252 19068
rect 26956 19014 27002 19066
rect 27002 19014 27012 19066
rect 27036 19014 27066 19066
rect 27066 19014 27078 19066
rect 27078 19014 27092 19066
rect 27116 19014 27130 19066
rect 27130 19014 27142 19066
rect 27142 19014 27172 19066
rect 27196 19014 27206 19066
rect 27206 19014 27252 19066
rect 26956 19012 27012 19014
rect 27036 19012 27092 19014
rect 27116 19012 27172 19014
rect 27196 19012 27252 19014
rect 26956 17978 27012 17980
rect 27036 17978 27092 17980
rect 27116 17978 27172 17980
rect 27196 17978 27252 17980
rect 26956 17926 27002 17978
rect 27002 17926 27012 17978
rect 27036 17926 27066 17978
rect 27066 17926 27078 17978
rect 27078 17926 27092 17978
rect 27116 17926 27130 17978
rect 27130 17926 27142 17978
rect 27142 17926 27172 17978
rect 27196 17926 27206 17978
rect 27206 17926 27252 17978
rect 26956 17924 27012 17926
rect 27036 17924 27092 17926
rect 27116 17924 27172 17926
rect 27196 17924 27252 17926
rect 26956 16890 27012 16892
rect 27036 16890 27092 16892
rect 27116 16890 27172 16892
rect 27196 16890 27252 16892
rect 26956 16838 27002 16890
rect 27002 16838 27012 16890
rect 27036 16838 27066 16890
rect 27066 16838 27078 16890
rect 27078 16838 27092 16890
rect 27116 16838 27130 16890
rect 27130 16838 27142 16890
rect 27142 16838 27172 16890
rect 27196 16838 27206 16890
rect 27206 16838 27252 16890
rect 26956 16836 27012 16838
rect 27036 16836 27092 16838
rect 27116 16836 27172 16838
rect 27196 16836 27252 16838
rect 26956 15802 27012 15804
rect 27036 15802 27092 15804
rect 27116 15802 27172 15804
rect 27196 15802 27252 15804
rect 26956 15750 27002 15802
rect 27002 15750 27012 15802
rect 27036 15750 27066 15802
rect 27066 15750 27078 15802
rect 27078 15750 27092 15802
rect 27116 15750 27130 15802
rect 27130 15750 27142 15802
rect 27142 15750 27172 15802
rect 27196 15750 27206 15802
rect 27206 15750 27252 15802
rect 26956 15748 27012 15750
rect 27036 15748 27092 15750
rect 27116 15748 27172 15750
rect 27196 15748 27252 15750
rect 26956 14714 27012 14716
rect 27036 14714 27092 14716
rect 27116 14714 27172 14716
rect 27196 14714 27252 14716
rect 26956 14662 27002 14714
rect 27002 14662 27012 14714
rect 27036 14662 27066 14714
rect 27066 14662 27078 14714
rect 27078 14662 27092 14714
rect 27116 14662 27130 14714
rect 27130 14662 27142 14714
rect 27142 14662 27172 14714
rect 27196 14662 27206 14714
rect 27206 14662 27252 14714
rect 26956 14660 27012 14662
rect 27036 14660 27092 14662
rect 27116 14660 27172 14662
rect 27196 14660 27252 14662
rect 26956 13626 27012 13628
rect 27036 13626 27092 13628
rect 27116 13626 27172 13628
rect 27196 13626 27252 13628
rect 26956 13574 27002 13626
rect 27002 13574 27012 13626
rect 27036 13574 27066 13626
rect 27066 13574 27078 13626
rect 27078 13574 27092 13626
rect 27116 13574 27130 13626
rect 27130 13574 27142 13626
rect 27142 13574 27172 13626
rect 27196 13574 27206 13626
rect 27206 13574 27252 13626
rect 26956 13572 27012 13574
rect 27036 13572 27092 13574
rect 27116 13572 27172 13574
rect 27196 13572 27252 13574
rect 27616 20698 27672 20700
rect 27696 20698 27752 20700
rect 27776 20698 27832 20700
rect 27856 20698 27912 20700
rect 27616 20646 27662 20698
rect 27662 20646 27672 20698
rect 27696 20646 27726 20698
rect 27726 20646 27738 20698
rect 27738 20646 27752 20698
rect 27776 20646 27790 20698
rect 27790 20646 27802 20698
rect 27802 20646 27832 20698
rect 27856 20646 27866 20698
rect 27866 20646 27912 20698
rect 27616 20644 27672 20646
rect 27696 20644 27752 20646
rect 27776 20644 27832 20646
rect 27856 20644 27912 20646
rect 27616 19610 27672 19612
rect 27696 19610 27752 19612
rect 27776 19610 27832 19612
rect 27856 19610 27912 19612
rect 27616 19558 27662 19610
rect 27662 19558 27672 19610
rect 27696 19558 27726 19610
rect 27726 19558 27738 19610
rect 27738 19558 27752 19610
rect 27776 19558 27790 19610
rect 27790 19558 27802 19610
rect 27802 19558 27832 19610
rect 27856 19558 27866 19610
rect 27866 19558 27912 19610
rect 27616 19556 27672 19558
rect 27696 19556 27752 19558
rect 27776 19556 27832 19558
rect 27856 19556 27912 19558
rect 27616 18522 27672 18524
rect 27696 18522 27752 18524
rect 27776 18522 27832 18524
rect 27856 18522 27912 18524
rect 27616 18470 27662 18522
rect 27662 18470 27672 18522
rect 27696 18470 27726 18522
rect 27726 18470 27738 18522
rect 27738 18470 27752 18522
rect 27776 18470 27790 18522
rect 27790 18470 27802 18522
rect 27802 18470 27832 18522
rect 27856 18470 27866 18522
rect 27866 18470 27912 18522
rect 27616 18468 27672 18470
rect 27696 18468 27752 18470
rect 27776 18468 27832 18470
rect 27856 18468 27912 18470
rect 27616 17434 27672 17436
rect 27696 17434 27752 17436
rect 27776 17434 27832 17436
rect 27856 17434 27912 17436
rect 27616 17382 27662 17434
rect 27662 17382 27672 17434
rect 27696 17382 27726 17434
rect 27726 17382 27738 17434
rect 27738 17382 27752 17434
rect 27776 17382 27790 17434
rect 27790 17382 27802 17434
rect 27802 17382 27832 17434
rect 27856 17382 27866 17434
rect 27866 17382 27912 17434
rect 27616 17380 27672 17382
rect 27696 17380 27752 17382
rect 27776 17380 27832 17382
rect 27856 17380 27912 17382
rect 27616 16346 27672 16348
rect 27696 16346 27752 16348
rect 27776 16346 27832 16348
rect 27856 16346 27912 16348
rect 27616 16294 27662 16346
rect 27662 16294 27672 16346
rect 27696 16294 27726 16346
rect 27726 16294 27738 16346
rect 27738 16294 27752 16346
rect 27776 16294 27790 16346
rect 27790 16294 27802 16346
rect 27802 16294 27832 16346
rect 27856 16294 27866 16346
rect 27866 16294 27912 16346
rect 27616 16292 27672 16294
rect 27696 16292 27752 16294
rect 27776 16292 27832 16294
rect 27856 16292 27912 16294
rect 27616 15258 27672 15260
rect 27696 15258 27752 15260
rect 27776 15258 27832 15260
rect 27856 15258 27912 15260
rect 27616 15206 27662 15258
rect 27662 15206 27672 15258
rect 27696 15206 27726 15258
rect 27726 15206 27738 15258
rect 27738 15206 27752 15258
rect 27776 15206 27790 15258
rect 27790 15206 27802 15258
rect 27802 15206 27832 15258
rect 27856 15206 27866 15258
rect 27866 15206 27912 15258
rect 27616 15204 27672 15206
rect 27696 15204 27752 15206
rect 27776 15204 27832 15206
rect 27856 15204 27912 15206
rect 27616 14170 27672 14172
rect 27696 14170 27752 14172
rect 27776 14170 27832 14172
rect 27856 14170 27912 14172
rect 27616 14118 27662 14170
rect 27662 14118 27672 14170
rect 27696 14118 27726 14170
rect 27726 14118 27738 14170
rect 27738 14118 27752 14170
rect 27776 14118 27790 14170
rect 27790 14118 27802 14170
rect 27802 14118 27832 14170
rect 27856 14118 27866 14170
rect 27866 14118 27912 14170
rect 27616 14116 27672 14118
rect 27696 14116 27752 14118
rect 27776 14116 27832 14118
rect 27856 14116 27912 14118
rect 27616 13082 27672 13084
rect 27696 13082 27752 13084
rect 27776 13082 27832 13084
rect 27856 13082 27912 13084
rect 27616 13030 27662 13082
rect 27662 13030 27672 13082
rect 27696 13030 27726 13082
rect 27726 13030 27738 13082
rect 27738 13030 27752 13082
rect 27776 13030 27790 13082
rect 27790 13030 27802 13082
rect 27802 13030 27832 13082
rect 27856 13030 27866 13082
rect 27866 13030 27912 13082
rect 27616 13028 27672 13030
rect 27696 13028 27752 13030
rect 27776 13028 27832 13030
rect 27856 13028 27912 13030
rect 26956 12538 27012 12540
rect 27036 12538 27092 12540
rect 27116 12538 27172 12540
rect 27196 12538 27252 12540
rect 26956 12486 27002 12538
rect 27002 12486 27012 12538
rect 27036 12486 27066 12538
rect 27066 12486 27078 12538
rect 27078 12486 27092 12538
rect 27116 12486 27130 12538
rect 27130 12486 27142 12538
rect 27142 12486 27172 12538
rect 27196 12486 27206 12538
rect 27206 12486 27252 12538
rect 26956 12484 27012 12486
rect 27036 12484 27092 12486
rect 27116 12484 27172 12486
rect 27196 12484 27252 12486
rect 27616 11994 27672 11996
rect 27696 11994 27752 11996
rect 27776 11994 27832 11996
rect 27856 11994 27912 11996
rect 27616 11942 27662 11994
rect 27662 11942 27672 11994
rect 27696 11942 27726 11994
rect 27726 11942 27738 11994
rect 27738 11942 27752 11994
rect 27776 11942 27790 11994
rect 27790 11942 27802 11994
rect 27802 11942 27832 11994
rect 27856 11942 27866 11994
rect 27866 11942 27912 11994
rect 27616 11940 27672 11942
rect 27696 11940 27752 11942
rect 27776 11940 27832 11942
rect 27856 11940 27912 11942
rect 26956 11450 27012 11452
rect 27036 11450 27092 11452
rect 27116 11450 27172 11452
rect 27196 11450 27252 11452
rect 26956 11398 27002 11450
rect 27002 11398 27012 11450
rect 27036 11398 27066 11450
rect 27066 11398 27078 11450
rect 27078 11398 27092 11450
rect 27116 11398 27130 11450
rect 27130 11398 27142 11450
rect 27142 11398 27172 11450
rect 27196 11398 27206 11450
rect 27206 11398 27252 11450
rect 26956 11396 27012 11398
rect 27036 11396 27092 11398
rect 27116 11396 27172 11398
rect 27196 11396 27252 11398
rect 27616 10906 27672 10908
rect 27696 10906 27752 10908
rect 27776 10906 27832 10908
rect 27856 10906 27912 10908
rect 27616 10854 27662 10906
rect 27662 10854 27672 10906
rect 27696 10854 27726 10906
rect 27726 10854 27738 10906
rect 27738 10854 27752 10906
rect 27776 10854 27790 10906
rect 27790 10854 27802 10906
rect 27802 10854 27832 10906
rect 27856 10854 27866 10906
rect 27866 10854 27912 10906
rect 27616 10852 27672 10854
rect 27696 10852 27752 10854
rect 27776 10852 27832 10854
rect 27856 10852 27912 10854
rect 26956 10362 27012 10364
rect 27036 10362 27092 10364
rect 27116 10362 27172 10364
rect 27196 10362 27252 10364
rect 26956 10310 27002 10362
rect 27002 10310 27012 10362
rect 27036 10310 27066 10362
rect 27066 10310 27078 10362
rect 27078 10310 27092 10362
rect 27116 10310 27130 10362
rect 27130 10310 27142 10362
rect 27142 10310 27172 10362
rect 27196 10310 27206 10362
rect 27206 10310 27252 10362
rect 26956 10308 27012 10310
rect 27036 10308 27092 10310
rect 27116 10308 27172 10310
rect 27196 10308 27252 10310
rect 27616 9818 27672 9820
rect 27696 9818 27752 9820
rect 27776 9818 27832 9820
rect 27856 9818 27912 9820
rect 27616 9766 27662 9818
rect 27662 9766 27672 9818
rect 27696 9766 27726 9818
rect 27726 9766 27738 9818
rect 27738 9766 27752 9818
rect 27776 9766 27790 9818
rect 27790 9766 27802 9818
rect 27802 9766 27832 9818
rect 27856 9766 27866 9818
rect 27866 9766 27912 9818
rect 27616 9764 27672 9766
rect 27696 9764 27752 9766
rect 27776 9764 27832 9766
rect 27856 9764 27912 9766
rect 26956 9274 27012 9276
rect 27036 9274 27092 9276
rect 27116 9274 27172 9276
rect 27196 9274 27252 9276
rect 26956 9222 27002 9274
rect 27002 9222 27012 9274
rect 27036 9222 27066 9274
rect 27066 9222 27078 9274
rect 27078 9222 27092 9274
rect 27116 9222 27130 9274
rect 27130 9222 27142 9274
rect 27142 9222 27172 9274
rect 27196 9222 27206 9274
rect 27206 9222 27252 9274
rect 26956 9220 27012 9222
rect 27036 9220 27092 9222
rect 27116 9220 27172 9222
rect 27196 9220 27252 9222
rect 27616 8730 27672 8732
rect 27696 8730 27752 8732
rect 27776 8730 27832 8732
rect 27856 8730 27912 8732
rect 27616 8678 27662 8730
rect 27662 8678 27672 8730
rect 27696 8678 27726 8730
rect 27726 8678 27738 8730
rect 27738 8678 27752 8730
rect 27776 8678 27790 8730
rect 27790 8678 27802 8730
rect 27802 8678 27832 8730
rect 27856 8678 27866 8730
rect 27866 8678 27912 8730
rect 27616 8676 27672 8678
rect 27696 8676 27752 8678
rect 27776 8676 27832 8678
rect 27856 8676 27912 8678
rect 26956 8186 27012 8188
rect 27036 8186 27092 8188
rect 27116 8186 27172 8188
rect 27196 8186 27252 8188
rect 26956 8134 27002 8186
rect 27002 8134 27012 8186
rect 27036 8134 27066 8186
rect 27066 8134 27078 8186
rect 27078 8134 27092 8186
rect 27116 8134 27130 8186
rect 27130 8134 27142 8186
rect 27142 8134 27172 8186
rect 27196 8134 27206 8186
rect 27206 8134 27252 8186
rect 26956 8132 27012 8134
rect 27036 8132 27092 8134
rect 27116 8132 27172 8134
rect 27196 8132 27252 8134
rect 27616 7642 27672 7644
rect 27696 7642 27752 7644
rect 27776 7642 27832 7644
rect 27856 7642 27912 7644
rect 27616 7590 27662 7642
rect 27662 7590 27672 7642
rect 27696 7590 27726 7642
rect 27726 7590 27738 7642
rect 27738 7590 27752 7642
rect 27776 7590 27790 7642
rect 27790 7590 27802 7642
rect 27802 7590 27832 7642
rect 27856 7590 27866 7642
rect 27866 7590 27912 7642
rect 27616 7588 27672 7590
rect 27696 7588 27752 7590
rect 27776 7588 27832 7590
rect 27856 7588 27912 7590
rect 26956 7098 27012 7100
rect 27036 7098 27092 7100
rect 27116 7098 27172 7100
rect 27196 7098 27252 7100
rect 26956 7046 27002 7098
rect 27002 7046 27012 7098
rect 27036 7046 27066 7098
rect 27066 7046 27078 7098
rect 27078 7046 27092 7098
rect 27116 7046 27130 7098
rect 27130 7046 27142 7098
rect 27142 7046 27172 7098
rect 27196 7046 27206 7098
rect 27206 7046 27252 7098
rect 26956 7044 27012 7046
rect 27036 7044 27092 7046
rect 27116 7044 27172 7046
rect 27196 7044 27252 7046
rect 27616 6554 27672 6556
rect 27696 6554 27752 6556
rect 27776 6554 27832 6556
rect 27856 6554 27912 6556
rect 27616 6502 27662 6554
rect 27662 6502 27672 6554
rect 27696 6502 27726 6554
rect 27726 6502 27738 6554
rect 27738 6502 27752 6554
rect 27776 6502 27790 6554
rect 27790 6502 27802 6554
rect 27802 6502 27832 6554
rect 27856 6502 27866 6554
rect 27866 6502 27912 6554
rect 27616 6500 27672 6502
rect 27696 6500 27752 6502
rect 27776 6500 27832 6502
rect 27856 6500 27912 6502
rect 26956 6010 27012 6012
rect 27036 6010 27092 6012
rect 27116 6010 27172 6012
rect 27196 6010 27252 6012
rect 26956 5958 27002 6010
rect 27002 5958 27012 6010
rect 27036 5958 27066 6010
rect 27066 5958 27078 6010
rect 27078 5958 27092 6010
rect 27116 5958 27130 6010
rect 27130 5958 27142 6010
rect 27142 5958 27172 6010
rect 27196 5958 27206 6010
rect 27206 5958 27252 6010
rect 26956 5956 27012 5958
rect 27036 5956 27092 5958
rect 27116 5956 27172 5958
rect 27196 5956 27252 5958
rect 27616 5466 27672 5468
rect 27696 5466 27752 5468
rect 27776 5466 27832 5468
rect 27856 5466 27912 5468
rect 27616 5414 27662 5466
rect 27662 5414 27672 5466
rect 27696 5414 27726 5466
rect 27726 5414 27738 5466
rect 27738 5414 27752 5466
rect 27776 5414 27790 5466
rect 27790 5414 27802 5466
rect 27802 5414 27832 5466
rect 27856 5414 27866 5466
rect 27866 5414 27912 5466
rect 27616 5412 27672 5414
rect 27696 5412 27752 5414
rect 27776 5412 27832 5414
rect 27856 5412 27912 5414
rect 26956 4922 27012 4924
rect 27036 4922 27092 4924
rect 27116 4922 27172 4924
rect 27196 4922 27252 4924
rect 26956 4870 27002 4922
rect 27002 4870 27012 4922
rect 27036 4870 27066 4922
rect 27066 4870 27078 4922
rect 27078 4870 27092 4922
rect 27116 4870 27130 4922
rect 27130 4870 27142 4922
rect 27142 4870 27172 4922
rect 27196 4870 27206 4922
rect 27206 4870 27252 4922
rect 26956 4868 27012 4870
rect 27036 4868 27092 4870
rect 27116 4868 27172 4870
rect 27196 4868 27252 4870
rect 22616 4378 22672 4380
rect 22696 4378 22752 4380
rect 22776 4378 22832 4380
rect 22856 4378 22912 4380
rect 22616 4326 22662 4378
rect 22662 4326 22672 4378
rect 22696 4326 22726 4378
rect 22726 4326 22738 4378
rect 22738 4326 22752 4378
rect 22776 4326 22790 4378
rect 22790 4326 22802 4378
rect 22802 4326 22832 4378
rect 22856 4326 22866 4378
rect 22866 4326 22912 4378
rect 22616 4324 22672 4326
rect 22696 4324 22752 4326
rect 22776 4324 22832 4326
rect 22856 4324 22912 4326
rect 27616 4378 27672 4380
rect 27696 4378 27752 4380
rect 27776 4378 27832 4380
rect 27856 4378 27912 4380
rect 27616 4326 27662 4378
rect 27662 4326 27672 4378
rect 27696 4326 27726 4378
rect 27726 4326 27738 4378
rect 27738 4326 27752 4378
rect 27776 4326 27790 4378
rect 27790 4326 27802 4378
rect 27802 4326 27832 4378
rect 27856 4326 27866 4378
rect 27866 4326 27912 4378
rect 27616 4324 27672 4326
rect 27696 4324 27752 4326
rect 27776 4324 27832 4326
rect 27856 4324 27912 4326
rect 21956 3834 22012 3836
rect 22036 3834 22092 3836
rect 22116 3834 22172 3836
rect 22196 3834 22252 3836
rect 21956 3782 22002 3834
rect 22002 3782 22012 3834
rect 22036 3782 22066 3834
rect 22066 3782 22078 3834
rect 22078 3782 22092 3834
rect 22116 3782 22130 3834
rect 22130 3782 22142 3834
rect 22142 3782 22172 3834
rect 22196 3782 22206 3834
rect 22206 3782 22252 3834
rect 21956 3780 22012 3782
rect 22036 3780 22092 3782
rect 22116 3780 22172 3782
rect 22196 3780 22252 3782
rect 26956 3834 27012 3836
rect 27036 3834 27092 3836
rect 27116 3834 27172 3836
rect 27196 3834 27252 3836
rect 26956 3782 27002 3834
rect 27002 3782 27012 3834
rect 27036 3782 27066 3834
rect 27066 3782 27078 3834
rect 27078 3782 27092 3834
rect 27116 3782 27130 3834
rect 27130 3782 27142 3834
rect 27142 3782 27172 3834
rect 27196 3782 27206 3834
rect 27206 3782 27252 3834
rect 26956 3780 27012 3782
rect 27036 3780 27092 3782
rect 27116 3780 27172 3782
rect 27196 3780 27252 3782
rect 22616 3290 22672 3292
rect 22696 3290 22752 3292
rect 22776 3290 22832 3292
rect 22856 3290 22912 3292
rect 22616 3238 22662 3290
rect 22662 3238 22672 3290
rect 22696 3238 22726 3290
rect 22726 3238 22738 3290
rect 22738 3238 22752 3290
rect 22776 3238 22790 3290
rect 22790 3238 22802 3290
rect 22802 3238 22832 3290
rect 22856 3238 22866 3290
rect 22866 3238 22912 3290
rect 22616 3236 22672 3238
rect 22696 3236 22752 3238
rect 22776 3236 22832 3238
rect 22856 3236 22912 3238
rect 27616 3290 27672 3292
rect 27696 3290 27752 3292
rect 27776 3290 27832 3292
rect 27856 3290 27912 3292
rect 27616 3238 27662 3290
rect 27662 3238 27672 3290
rect 27696 3238 27726 3290
rect 27726 3238 27738 3290
rect 27738 3238 27752 3290
rect 27776 3238 27790 3290
rect 27790 3238 27802 3290
rect 27802 3238 27832 3290
rect 27856 3238 27866 3290
rect 27866 3238 27912 3290
rect 27616 3236 27672 3238
rect 27696 3236 27752 3238
rect 27776 3236 27832 3238
rect 27856 3236 27912 3238
rect 30562 28736 30618 28792
rect 31956 68026 32012 68028
rect 32036 68026 32092 68028
rect 32116 68026 32172 68028
rect 32196 68026 32252 68028
rect 31956 67974 32002 68026
rect 32002 67974 32012 68026
rect 32036 67974 32066 68026
rect 32066 67974 32078 68026
rect 32078 67974 32092 68026
rect 32116 67974 32130 68026
rect 32130 67974 32142 68026
rect 32142 67974 32172 68026
rect 32196 67974 32206 68026
rect 32206 67974 32252 68026
rect 31956 67972 32012 67974
rect 32036 67972 32092 67974
rect 32116 67972 32172 67974
rect 32196 67972 32252 67974
rect 32402 67632 32458 67688
rect 32616 67482 32672 67484
rect 32696 67482 32752 67484
rect 32776 67482 32832 67484
rect 32856 67482 32912 67484
rect 32616 67430 32662 67482
rect 32662 67430 32672 67482
rect 32696 67430 32726 67482
rect 32726 67430 32738 67482
rect 32738 67430 32752 67482
rect 32776 67430 32790 67482
rect 32790 67430 32802 67482
rect 32802 67430 32832 67482
rect 32856 67430 32866 67482
rect 32866 67430 32912 67482
rect 32616 67428 32672 67430
rect 32696 67428 32752 67430
rect 32776 67428 32832 67430
rect 32856 67428 32912 67430
rect 31956 66938 32012 66940
rect 32036 66938 32092 66940
rect 32116 66938 32172 66940
rect 32196 66938 32252 66940
rect 31956 66886 32002 66938
rect 32002 66886 32012 66938
rect 32036 66886 32066 66938
rect 32066 66886 32078 66938
rect 32078 66886 32092 66938
rect 32116 66886 32130 66938
rect 32130 66886 32142 66938
rect 32142 66886 32172 66938
rect 32196 66886 32206 66938
rect 32206 66886 32252 66938
rect 31956 66884 32012 66886
rect 32036 66884 32092 66886
rect 32116 66884 32172 66886
rect 32196 66884 32252 66886
rect 32616 66394 32672 66396
rect 32696 66394 32752 66396
rect 32776 66394 32832 66396
rect 32856 66394 32912 66396
rect 32616 66342 32662 66394
rect 32662 66342 32672 66394
rect 32696 66342 32726 66394
rect 32726 66342 32738 66394
rect 32738 66342 32752 66394
rect 32776 66342 32790 66394
rect 32790 66342 32802 66394
rect 32802 66342 32832 66394
rect 32856 66342 32866 66394
rect 32866 66342 32912 66394
rect 32616 66340 32672 66342
rect 32696 66340 32752 66342
rect 32776 66340 32832 66342
rect 32856 66340 32912 66342
rect 31956 65850 32012 65852
rect 32036 65850 32092 65852
rect 32116 65850 32172 65852
rect 32196 65850 32252 65852
rect 31956 65798 32002 65850
rect 32002 65798 32012 65850
rect 32036 65798 32066 65850
rect 32066 65798 32078 65850
rect 32078 65798 32092 65850
rect 32116 65798 32130 65850
rect 32130 65798 32142 65850
rect 32142 65798 32172 65850
rect 32196 65798 32206 65850
rect 32206 65798 32252 65850
rect 31956 65796 32012 65798
rect 32036 65796 32092 65798
rect 32116 65796 32172 65798
rect 32196 65796 32252 65798
rect 32616 65306 32672 65308
rect 32696 65306 32752 65308
rect 32776 65306 32832 65308
rect 32856 65306 32912 65308
rect 32616 65254 32662 65306
rect 32662 65254 32672 65306
rect 32696 65254 32726 65306
rect 32726 65254 32738 65306
rect 32738 65254 32752 65306
rect 32776 65254 32790 65306
rect 32790 65254 32802 65306
rect 32802 65254 32832 65306
rect 32856 65254 32866 65306
rect 32866 65254 32912 65306
rect 32616 65252 32672 65254
rect 32696 65252 32752 65254
rect 32776 65252 32832 65254
rect 32856 65252 32912 65254
rect 31956 64762 32012 64764
rect 32036 64762 32092 64764
rect 32116 64762 32172 64764
rect 32196 64762 32252 64764
rect 31956 64710 32002 64762
rect 32002 64710 32012 64762
rect 32036 64710 32066 64762
rect 32066 64710 32078 64762
rect 32078 64710 32092 64762
rect 32116 64710 32130 64762
rect 32130 64710 32142 64762
rect 32142 64710 32172 64762
rect 32196 64710 32206 64762
rect 32206 64710 32252 64762
rect 31956 64708 32012 64710
rect 32036 64708 32092 64710
rect 32116 64708 32172 64710
rect 32196 64708 32252 64710
rect 32616 64218 32672 64220
rect 32696 64218 32752 64220
rect 32776 64218 32832 64220
rect 32856 64218 32912 64220
rect 32616 64166 32662 64218
rect 32662 64166 32672 64218
rect 32696 64166 32726 64218
rect 32726 64166 32738 64218
rect 32738 64166 32752 64218
rect 32776 64166 32790 64218
rect 32790 64166 32802 64218
rect 32802 64166 32832 64218
rect 32856 64166 32866 64218
rect 32866 64166 32912 64218
rect 32616 64164 32672 64166
rect 32696 64164 32752 64166
rect 32776 64164 32832 64166
rect 32856 64164 32912 64166
rect 31956 63674 32012 63676
rect 32036 63674 32092 63676
rect 32116 63674 32172 63676
rect 32196 63674 32252 63676
rect 31956 63622 32002 63674
rect 32002 63622 32012 63674
rect 32036 63622 32066 63674
rect 32066 63622 32078 63674
rect 32078 63622 32092 63674
rect 32116 63622 32130 63674
rect 32130 63622 32142 63674
rect 32142 63622 32172 63674
rect 32196 63622 32206 63674
rect 32206 63622 32252 63674
rect 31956 63620 32012 63622
rect 32036 63620 32092 63622
rect 32116 63620 32172 63622
rect 32196 63620 32252 63622
rect 31956 62586 32012 62588
rect 32036 62586 32092 62588
rect 32116 62586 32172 62588
rect 32196 62586 32252 62588
rect 31956 62534 32002 62586
rect 32002 62534 32012 62586
rect 32036 62534 32066 62586
rect 32066 62534 32078 62586
rect 32078 62534 32092 62586
rect 32116 62534 32130 62586
rect 32130 62534 32142 62586
rect 32142 62534 32172 62586
rect 32196 62534 32206 62586
rect 32206 62534 32252 62586
rect 31956 62532 32012 62534
rect 32036 62532 32092 62534
rect 32116 62532 32172 62534
rect 32196 62532 32252 62534
rect 31956 61498 32012 61500
rect 32036 61498 32092 61500
rect 32116 61498 32172 61500
rect 32196 61498 32252 61500
rect 31956 61446 32002 61498
rect 32002 61446 32012 61498
rect 32036 61446 32066 61498
rect 32066 61446 32078 61498
rect 32078 61446 32092 61498
rect 32116 61446 32130 61498
rect 32130 61446 32142 61498
rect 32142 61446 32172 61498
rect 32196 61446 32206 61498
rect 32206 61446 32252 61498
rect 31956 61444 32012 61446
rect 32036 61444 32092 61446
rect 32116 61444 32172 61446
rect 32196 61444 32252 61446
rect 31956 60410 32012 60412
rect 32036 60410 32092 60412
rect 32116 60410 32172 60412
rect 32196 60410 32252 60412
rect 31956 60358 32002 60410
rect 32002 60358 32012 60410
rect 32036 60358 32066 60410
rect 32066 60358 32078 60410
rect 32078 60358 32092 60410
rect 32116 60358 32130 60410
rect 32130 60358 32142 60410
rect 32142 60358 32172 60410
rect 32196 60358 32206 60410
rect 32206 60358 32252 60410
rect 31956 60356 32012 60358
rect 32036 60356 32092 60358
rect 32116 60356 32172 60358
rect 32196 60356 32252 60358
rect 31956 59322 32012 59324
rect 32036 59322 32092 59324
rect 32116 59322 32172 59324
rect 32196 59322 32252 59324
rect 31956 59270 32002 59322
rect 32002 59270 32012 59322
rect 32036 59270 32066 59322
rect 32066 59270 32078 59322
rect 32078 59270 32092 59322
rect 32116 59270 32130 59322
rect 32130 59270 32142 59322
rect 32142 59270 32172 59322
rect 32196 59270 32206 59322
rect 32206 59270 32252 59322
rect 31956 59268 32012 59270
rect 32036 59268 32092 59270
rect 32116 59268 32172 59270
rect 32196 59268 32252 59270
rect 31956 58234 32012 58236
rect 32036 58234 32092 58236
rect 32116 58234 32172 58236
rect 32196 58234 32252 58236
rect 31956 58182 32002 58234
rect 32002 58182 32012 58234
rect 32036 58182 32066 58234
rect 32066 58182 32078 58234
rect 32078 58182 32092 58234
rect 32116 58182 32130 58234
rect 32130 58182 32142 58234
rect 32142 58182 32172 58234
rect 32196 58182 32206 58234
rect 32206 58182 32252 58234
rect 31956 58180 32012 58182
rect 32036 58180 32092 58182
rect 32116 58180 32172 58182
rect 32196 58180 32252 58182
rect 31956 57146 32012 57148
rect 32036 57146 32092 57148
rect 32116 57146 32172 57148
rect 32196 57146 32252 57148
rect 31956 57094 32002 57146
rect 32002 57094 32012 57146
rect 32036 57094 32066 57146
rect 32066 57094 32078 57146
rect 32078 57094 32092 57146
rect 32116 57094 32130 57146
rect 32130 57094 32142 57146
rect 32142 57094 32172 57146
rect 32196 57094 32206 57146
rect 32206 57094 32252 57146
rect 31956 57092 32012 57094
rect 32036 57092 32092 57094
rect 32116 57092 32172 57094
rect 32196 57092 32252 57094
rect 31956 56058 32012 56060
rect 32036 56058 32092 56060
rect 32116 56058 32172 56060
rect 32196 56058 32252 56060
rect 31956 56006 32002 56058
rect 32002 56006 32012 56058
rect 32036 56006 32066 56058
rect 32066 56006 32078 56058
rect 32078 56006 32092 56058
rect 32116 56006 32130 56058
rect 32130 56006 32142 56058
rect 32142 56006 32172 56058
rect 32196 56006 32206 56058
rect 32206 56006 32252 56058
rect 31956 56004 32012 56006
rect 32036 56004 32092 56006
rect 32116 56004 32172 56006
rect 32196 56004 32252 56006
rect 31956 54970 32012 54972
rect 32036 54970 32092 54972
rect 32116 54970 32172 54972
rect 32196 54970 32252 54972
rect 31956 54918 32002 54970
rect 32002 54918 32012 54970
rect 32036 54918 32066 54970
rect 32066 54918 32078 54970
rect 32078 54918 32092 54970
rect 32116 54918 32130 54970
rect 32130 54918 32142 54970
rect 32142 54918 32172 54970
rect 32196 54918 32206 54970
rect 32206 54918 32252 54970
rect 31956 54916 32012 54918
rect 32036 54916 32092 54918
rect 32116 54916 32172 54918
rect 32196 54916 32252 54918
rect 31956 53882 32012 53884
rect 32036 53882 32092 53884
rect 32116 53882 32172 53884
rect 32196 53882 32252 53884
rect 31956 53830 32002 53882
rect 32002 53830 32012 53882
rect 32036 53830 32066 53882
rect 32066 53830 32078 53882
rect 32078 53830 32092 53882
rect 32116 53830 32130 53882
rect 32130 53830 32142 53882
rect 32142 53830 32172 53882
rect 32196 53830 32206 53882
rect 32206 53830 32252 53882
rect 31956 53828 32012 53830
rect 32036 53828 32092 53830
rect 32116 53828 32172 53830
rect 32196 53828 32252 53830
rect 31956 52794 32012 52796
rect 32036 52794 32092 52796
rect 32116 52794 32172 52796
rect 32196 52794 32252 52796
rect 31956 52742 32002 52794
rect 32002 52742 32012 52794
rect 32036 52742 32066 52794
rect 32066 52742 32078 52794
rect 32078 52742 32092 52794
rect 32116 52742 32130 52794
rect 32130 52742 32142 52794
rect 32142 52742 32172 52794
rect 32196 52742 32206 52794
rect 32206 52742 32252 52794
rect 31956 52740 32012 52742
rect 32036 52740 32092 52742
rect 32116 52740 32172 52742
rect 32196 52740 32252 52742
rect 31956 51706 32012 51708
rect 32036 51706 32092 51708
rect 32116 51706 32172 51708
rect 32196 51706 32252 51708
rect 31956 51654 32002 51706
rect 32002 51654 32012 51706
rect 32036 51654 32066 51706
rect 32066 51654 32078 51706
rect 32078 51654 32092 51706
rect 32116 51654 32130 51706
rect 32130 51654 32142 51706
rect 32142 51654 32172 51706
rect 32196 51654 32206 51706
rect 32206 51654 32252 51706
rect 31956 51652 32012 51654
rect 32036 51652 32092 51654
rect 32116 51652 32172 51654
rect 32196 51652 32252 51654
rect 31956 50618 32012 50620
rect 32036 50618 32092 50620
rect 32116 50618 32172 50620
rect 32196 50618 32252 50620
rect 31956 50566 32002 50618
rect 32002 50566 32012 50618
rect 32036 50566 32066 50618
rect 32066 50566 32078 50618
rect 32078 50566 32092 50618
rect 32116 50566 32130 50618
rect 32130 50566 32142 50618
rect 32142 50566 32172 50618
rect 32196 50566 32206 50618
rect 32206 50566 32252 50618
rect 31956 50564 32012 50566
rect 32036 50564 32092 50566
rect 32116 50564 32172 50566
rect 32196 50564 32252 50566
rect 31956 49530 32012 49532
rect 32036 49530 32092 49532
rect 32116 49530 32172 49532
rect 32196 49530 32252 49532
rect 31956 49478 32002 49530
rect 32002 49478 32012 49530
rect 32036 49478 32066 49530
rect 32066 49478 32078 49530
rect 32078 49478 32092 49530
rect 32116 49478 32130 49530
rect 32130 49478 32142 49530
rect 32142 49478 32172 49530
rect 32196 49478 32206 49530
rect 32206 49478 32252 49530
rect 31956 49476 32012 49478
rect 32036 49476 32092 49478
rect 32116 49476 32172 49478
rect 32196 49476 32252 49478
rect 31956 48442 32012 48444
rect 32036 48442 32092 48444
rect 32116 48442 32172 48444
rect 32196 48442 32252 48444
rect 31956 48390 32002 48442
rect 32002 48390 32012 48442
rect 32036 48390 32066 48442
rect 32066 48390 32078 48442
rect 32078 48390 32092 48442
rect 32116 48390 32130 48442
rect 32130 48390 32142 48442
rect 32142 48390 32172 48442
rect 32196 48390 32206 48442
rect 32206 48390 32252 48442
rect 31956 48388 32012 48390
rect 32036 48388 32092 48390
rect 32116 48388 32172 48390
rect 32196 48388 32252 48390
rect 31956 47354 32012 47356
rect 32036 47354 32092 47356
rect 32116 47354 32172 47356
rect 32196 47354 32252 47356
rect 31956 47302 32002 47354
rect 32002 47302 32012 47354
rect 32036 47302 32066 47354
rect 32066 47302 32078 47354
rect 32078 47302 32092 47354
rect 32116 47302 32130 47354
rect 32130 47302 32142 47354
rect 32142 47302 32172 47354
rect 32196 47302 32206 47354
rect 32206 47302 32252 47354
rect 31956 47300 32012 47302
rect 32036 47300 32092 47302
rect 32116 47300 32172 47302
rect 32196 47300 32252 47302
rect 31956 46266 32012 46268
rect 32036 46266 32092 46268
rect 32116 46266 32172 46268
rect 32196 46266 32252 46268
rect 31956 46214 32002 46266
rect 32002 46214 32012 46266
rect 32036 46214 32066 46266
rect 32066 46214 32078 46266
rect 32078 46214 32092 46266
rect 32116 46214 32130 46266
rect 32130 46214 32142 46266
rect 32142 46214 32172 46266
rect 32196 46214 32206 46266
rect 32206 46214 32252 46266
rect 31956 46212 32012 46214
rect 32036 46212 32092 46214
rect 32116 46212 32172 46214
rect 32196 46212 32252 46214
rect 31956 45178 32012 45180
rect 32036 45178 32092 45180
rect 32116 45178 32172 45180
rect 32196 45178 32252 45180
rect 31956 45126 32002 45178
rect 32002 45126 32012 45178
rect 32036 45126 32066 45178
rect 32066 45126 32078 45178
rect 32078 45126 32092 45178
rect 32116 45126 32130 45178
rect 32130 45126 32142 45178
rect 32142 45126 32172 45178
rect 32196 45126 32206 45178
rect 32206 45126 32252 45178
rect 31956 45124 32012 45126
rect 32036 45124 32092 45126
rect 32116 45124 32172 45126
rect 32196 45124 32252 45126
rect 31956 44090 32012 44092
rect 32036 44090 32092 44092
rect 32116 44090 32172 44092
rect 32196 44090 32252 44092
rect 31956 44038 32002 44090
rect 32002 44038 32012 44090
rect 32036 44038 32066 44090
rect 32066 44038 32078 44090
rect 32078 44038 32092 44090
rect 32116 44038 32130 44090
rect 32130 44038 32142 44090
rect 32142 44038 32172 44090
rect 32196 44038 32206 44090
rect 32206 44038 32252 44090
rect 31956 44036 32012 44038
rect 32036 44036 32092 44038
rect 32116 44036 32172 44038
rect 32196 44036 32252 44038
rect 31956 43002 32012 43004
rect 32036 43002 32092 43004
rect 32116 43002 32172 43004
rect 32196 43002 32252 43004
rect 31956 42950 32002 43002
rect 32002 42950 32012 43002
rect 32036 42950 32066 43002
rect 32066 42950 32078 43002
rect 32078 42950 32092 43002
rect 32116 42950 32130 43002
rect 32130 42950 32142 43002
rect 32142 42950 32172 43002
rect 32196 42950 32206 43002
rect 32206 42950 32252 43002
rect 31956 42948 32012 42950
rect 32036 42948 32092 42950
rect 32116 42948 32172 42950
rect 32196 42948 32252 42950
rect 31956 41914 32012 41916
rect 32036 41914 32092 41916
rect 32116 41914 32172 41916
rect 32196 41914 32252 41916
rect 31956 41862 32002 41914
rect 32002 41862 32012 41914
rect 32036 41862 32066 41914
rect 32066 41862 32078 41914
rect 32078 41862 32092 41914
rect 32116 41862 32130 41914
rect 32130 41862 32142 41914
rect 32142 41862 32172 41914
rect 32196 41862 32206 41914
rect 32206 41862 32252 41914
rect 31956 41860 32012 41862
rect 32036 41860 32092 41862
rect 32116 41860 32172 41862
rect 32196 41860 32252 41862
rect 31956 40826 32012 40828
rect 32036 40826 32092 40828
rect 32116 40826 32172 40828
rect 32196 40826 32252 40828
rect 31956 40774 32002 40826
rect 32002 40774 32012 40826
rect 32036 40774 32066 40826
rect 32066 40774 32078 40826
rect 32078 40774 32092 40826
rect 32116 40774 32130 40826
rect 32130 40774 32142 40826
rect 32142 40774 32172 40826
rect 32196 40774 32206 40826
rect 32206 40774 32252 40826
rect 31956 40772 32012 40774
rect 32036 40772 32092 40774
rect 32116 40772 32172 40774
rect 32196 40772 32252 40774
rect 31956 39738 32012 39740
rect 32036 39738 32092 39740
rect 32116 39738 32172 39740
rect 32196 39738 32252 39740
rect 31956 39686 32002 39738
rect 32002 39686 32012 39738
rect 32036 39686 32066 39738
rect 32066 39686 32078 39738
rect 32078 39686 32092 39738
rect 32116 39686 32130 39738
rect 32130 39686 32142 39738
rect 32142 39686 32172 39738
rect 32196 39686 32206 39738
rect 32206 39686 32252 39738
rect 31956 39684 32012 39686
rect 32036 39684 32092 39686
rect 32116 39684 32172 39686
rect 32196 39684 32252 39686
rect 31956 38650 32012 38652
rect 32036 38650 32092 38652
rect 32116 38650 32172 38652
rect 32196 38650 32252 38652
rect 31956 38598 32002 38650
rect 32002 38598 32012 38650
rect 32036 38598 32066 38650
rect 32066 38598 32078 38650
rect 32078 38598 32092 38650
rect 32116 38598 32130 38650
rect 32130 38598 32142 38650
rect 32142 38598 32172 38650
rect 32196 38598 32206 38650
rect 32206 38598 32252 38650
rect 31956 38596 32012 38598
rect 32036 38596 32092 38598
rect 32116 38596 32172 38598
rect 32196 38596 32252 38598
rect 31956 37562 32012 37564
rect 32036 37562 32092 37564
rect 32116 37562 32172 37564
rect 32196 37562 32252 37564
rect 31956 37510 32002 37562
rect 32002 37510 32012 37562
rect 32036 37510 32066 37562
rect 32066 37510 32078 37562
rect 32078 37510 32092 37562
rect 32116 37510 32130 37562
rect 32130 37510 32142 37562
rect 32142 37510 32172 37562
rect 32196 37510 32206 37562
rect 32206 37510 32252 37562
rect 31956 37508 32012 37510
rect 32036 37508 32092 37510
rect 32116 37508 32172 37510
rect 32196 37508 32252 37510
rect 31956 36474 32012 36476
rect 32036 36474 32092 36476
rect 32116 36474 32172 36476
rect 32196 36474 32252 36476
rect 31956 36422 32002 36474
rect 32002 36422 32012 36474
rect 32036 36422 32066 36474
rect 32066 36422 32078 36474
rect 32078 36422 32092 36474
rect 32116 36422 32130 36474
rect 32130 36422 32142 36474
rect 32142 36422 32172 36474
rect 32196 36422 32206 36474
rect 32206 36422 32252 36474
rect 31956 36420 32012 36422
rect 32036 36420 32092 36422
rect 32116 36420 32172 36422
rect 32196 36420 32252 36422
rect 31956 35386 32012 35388
rect 32036 35386 32092 35388
rect 32116 35386 32172 35388
rect 32196 35386 32252 35388
rect 31956 35334 32002 35386
rect 32002 35334 32012 35386
rect 32036 35334 32066 35386
rect 32066 35334 32078 35386
rect 32078 35334 32092 35386
rect 32116 35334 32130 35386
rect 32130 35334 32142 35386
rect 32142 35334 32172 35386
rect 32196 35334 32206 35386
rect 32206 35334 32252 35386
rect 31956 35332 32012 35334
rect 32036 35332 32092 35334
rect 32116 35332 32172 35334
rect 32196 35332 32252 35334
rect 31956 34298 32012 34300
rect 32036 34298 32092 34300
rect 32116 34298 32172 34300
rect 32196 34298 32252 34300
rect 31956 34246 32002 34298
rect 32002 34246 32012 34298
rect 32036 34246 32066 34298
rect 32066 34246 32078 34298
rect 32078 34246 32092 34298
rect 32116 34246 32130 34298
rect 32130 34246 32142 34298
rect 32142 34246 32172 34298
rect 32196 34246 32206 34298
rect 32206 34246 32252 34298
rect 31956 34244 32012 34246
rect 32036 34244 32092 34246
rect 32116 34244 32172 34246
rect 32196 34244 32252 34246
rect 31956 33210 32012 33212
rect 32036 33210 32092 33212
rect 32116 33210 32172 33212
rect 32196 33210 32252 33212
rect 31956 33158 32002 33210
rect 32002 33158 32012 33210
rect 32036 33158 32066 33210
rect 32066 33158 32078 33210
rect 32078 33158 32092 33210
rect 32116 33158 32130 33210
rect 32130 33158 32142 33210
rect 32142 33158 32172 33210
rect 32196 33158 32206 33210
rect 32206 33158 32252 33210
rect 31956 33156 32012 33158
rect 32036 33156 32092 33158
rect 32116 33156 32172 33158
rect 32196 33156 32252 33158
rect 31956 32122 32012 32124
rect 32036 32122 32092 32124
rect 32116 32122 32172 32124
rect 32196 32122 32252 32124
rect 31956 32070 32002 32122
rect 32002 32070 32012 32122
rect 32036 32070 32066 32122
rect 32066 32070 32078 32122
rect 32078 32070 32092 32122
rect 32116 32070 32130 32122
rect 32130 32070 32142 32122
rect 32142 32070 32172 32122
rect 32196 32070 32206 32122
rect 32206 32070 32252 32122
rect 31956 32068 32012 32070
rect 32036 32068 32092 32070
rect 32116 32068 32172 32070
rect 32196 32068 32252 32070
rect 31956 31034 32012 31036
rect 32036 31034 32092 31036
rect 32116 31034 32172 31036
rect 32196 31034 32252 31036
rect 31956 30982 32002 31034
rect 32002 30982 32012 31034
rect 32036 30982 32066 31034
rect 32066 30982 32078 31034
rect 32078 30982 32092 31034
rect 32116 30982 32130 31034
rect 32130 30982 32142 31034
rect 32142 30982 32172 31034
rect 32196 30982 32206 31034
rect 32206 30982 32252 31034
rect 31956 30980 32012 30982
rect 32036 30980 32092 30982
rect 32116 30980 32172 30982
rect 32196 30980 32252 30982
rect 31956 29946 32012 29948
rect 32036 29946 32092 29948
rect 32116 29946 32172 29948
rect 32196 29946 32252 29948
rect 31956 29894 32002 29946
rect 32002 29894 32012 29946
rect 32036 29894 32066 29946
rect 32066 29894 32078 29946
rect 32078 29894 32092 29946
rect 32116 29894 32130 29946
rect 32130 29894 32142 29946
rect 32142 29894 32172 29946
rect 32196 29894 32206 29946
rect 32206 29894 32252 29946
rect 31956 29892 32012 29894
rect 32036 29892 32092 29894
rect 32116 29892 32172 29894
rect 32196 29892 32252 29894
rect 31956 28858 32012 28860
rect 32036 28858 32092 28860
rect 32116 28858 32172 28860
rect 32196 28858 32252 28860
rect 31956 28806 32002 28858
rect 32002 28806 32012 28858
rect 32036 28806 32066 28858
rect 32066 28806 32078 28858
rect 32078 28806 32092 28858
rect 32116 28806 32130 28858
rect 32130 28806 32142 28858
rect 32142 28806 32172 28858
rect 32196 28806 32206 28858
rect 32206 28806 32252 28858
rect 31956 28804 32012 28806
rect 32036 28804 32092 28806
rect 32116 28804 32172 28806
rect 32196 28804 32252 28806
rect 31956 27770 32012 27772
rect 32036 27770 32092 27772
rect 32116 27770 32172 27772
rect 32196 27770 32252 27772
rect 31956 27718 32002 27770
rect 32002 27718 32012 27770
rect 32036 27718 32066 27770
rect 32066 27718 32078 27770
rect 32078 27718 32092 27770
rect 32116 27718 32130 27770
rect 32130 27718 32142 27770
rect 32142 27718 32172 27770
rect 32196 27718 32206 27770
rect 32206 27718 32252 27770
rect 31956 27716 32012 27718
rect 32036 27716 32092 27718
rect 32116 27716 32172 27718
rect 32196 27716 32252 27718
rect 31956 26682 32012 26684
rect 32036 26682 32092 26684
rect 32116 26682 32172 26684
rect 32196 26682 32252 26684
rect 31956 26630 32002 26682
rect 32002 26630 32012 26682
rect 32036 26630 32066 26682
rect 32066 26630 32078 26682
rect 32078 26630 32092 26682
rect 32116 26630 32130 26682
rect 32130 26630 32142 26682
rect 32142 26630 32172 26682
rect 32196 26630 32206 26682
rect 32206 26630 32252 26682
rect 31956 26628 32012 26630
rect 32036 26628 32092 26630
rect 32116 26628 32172 26630
rect 32196 26628 32252 26630
rect 32616 63130 32672 63132
rect 32696 63130 32752 63132
rect 32776 63130 32832 63132
rect 32856 63130 32912 63132
rect 32616 63078 32662 63130
rect 32662 63078 32672 63130
rect 32696 63078 32726 63130
rect 32726 63078 32738 63130
rect 32738 63078 32752 63130
rect 32776 63078 32790 63130
rect 32790 63078 32802 63130
rect 32802 63078 32832 63130
rect 32856 63078 32866 63130
rect 32866 63078 32912 63130
rect 32616 63076 32672 63078
rect 32696 63076 32752 63078
rect 32776 63076 32832 63078
rect 32856 63076 32912 63078
rect 32616 62042 32672 62044
rect 32696 62042 32752 62044
rect 32776 62042 32832 62044
rect 32856 62042 32912 62044
rect 32616 61990 32662 62042
rect 32662 61990 32672 62042
rect 32696 61990 32726 62042
rect 32726 61990 32738 62042
rect 32738 61990 32752 62042
rect 32776 61990 32790 62042
rect 32790 61990 32802 62042
rect 32802 61990 32832 62042
rect 32856 61990 32866 62042
rect 32866 61990 32912 62042
rect 32616 61988 32672 61990
rect 32696 61988 32752 61990
rect 32776 61988 32832 61990
rect 32856 61988 32912 61990
rect 32616 60954 32672 60956
rect 32696 60954 32752 60956
rect 32776 60954 32832 60956
rect 32856 60954 32912 60956
rect 32616 60902 32662 60954
rect 32662 60902 32672 60954
rect 32696 60902 32726 60954
rect 32726 60902 32738 60954
rect 32738 60902 32752 60954
rect 32776 60902 32790 60954
rect 32790 60902 32802 60954
rect 32802 60902 32832 60954
rect 32856 60902 32866 60954
rect 32866 60902 32912 60954
rect 32616 60900 32672 60902
rect 32696 60900 32752 60902
rect 32776 60900 32832 60902
rect 32856 60900 32912 60902
rect 32616 59866 32672 59868
rect 32696 59866 32752 59868
rect 32776 59866 32832 59868
rect 32856 59866 32912 59868
rect 32616 59814 32662 59866
rect 32662 59814 32672 59866
rect 32696 59814 32726 59866
rect 32726 59814 32738 59866
rect 32738 59814 32752 59866
rect 32776 59814 32790 59866
rect 32790 59814 32802 59866
rect 32802 59814 32832 59866
rect 32856 59814 32866 59866
rect 32866 59814 32912 59866
rect 32616 59812 32672 59814
rect 32696 59812 32752 59814
rect 32776 59812 32832 59814
rect 32856 59812 32912 59814
rect 32616 58778 32672 58780
rect 32696 58778 32752 58780
rect 32776 58778 32832 58780
rect 32856 58778 32912 58780
rect 32616 58726 32662 58778
rect 32662 58726 32672 58778
rect 32696 58726 32726 58778
rect 32726 58726 32738 58778
rect 32738 58726 32752 58778
rect 32776 58726 32790 58778
rect 32790 58726 32802 58778
rect 32802 58726 32832 58778
rect 32856 58726 32866 58778
rect 32866 58726 32912 58778
rect 32616 58724 32672 58726
rect 32696 58724 32752 58726
rect 32776 58724 32832 58726
rect 32856 58724 32912 58726
rect 32616 57690 32672 57692
rect 32696 57690 32752 57692
rect 32776 57690 32832 57692
rect 32856 57690 32912 57692
rect 32616 57638 32662 57690
rect 32662 57638 32672 57690
rect 32696 57638 32726 57690
rect 32726 57638 32738 57690
rect 32738 57638 32752 57690
rect 32776 57638 32790 57690
rect 32790 57638 32802 57690
rect 32802 57638 32832 57690
rect 32856 57638 32866 57690
rect 32866 57638 32912 57690
rect 32616 57636 32672 57638
rect 32696 57636 32752 57638
rect 32776 57636 32832 57638
rect 32856 57636 32912 57638
rect 32616 56602 32672 56604
rect 32696 56602 32752 56604
rect 32776 56602 32832 56604
rect 32856 56602 32912 56604
rect 32616 56550 32662 56602
rect 32662 56550 32672 56602
rect 32696 56550 32726 56602
rect 32726 56550 32738 56602
rect 32738 56550 32752 56602
rect 32776 56550 32790 56602
rect 32790 56550 32802 56602
rect 32802 56550 32832 56602
rect 32856 56550 32866 56602
rect 32866 56550 32912 56602
rect 32616 56548 32672 56550
rect 32696 56548 32752 56550
rect 32776 56548 32832 56550
rect 32856 56548 32912 56550
rect 32616 55514 32672 55516
rect 32696 55514 32752 55516
rect 32776 55514 32832 55516
rect 32856 55514 32912 55516
rect 32616 55462 32662 55514
rect 32662 55462 32672 55514
rect 32696 55462 32726 55514
rect 32726 55462 32738 55514
rect 32738 55462 32752 55514
rect 32776 55462 32790 55514
rect 32790 55462 32802 55514
rect 32802 55462 32832 55514
rect 32856 55462 32866 55514
rect 32866 55462 32912 55514
rect 32616 55460 32672 55462
rect 32696 55460 32752 55462
rect 32776 55460 32832 55462
rect 32856 55460 32912 55462
rect 32616 54426 32672 54428
rect 32696 54426 32752 54428
rect 32776 54426 32832 54428
rect 32856 54426 32912 54428
rect 32616 54374 32662 54426
rect 32662 54374 32672 54426
rect 32696 54374 32726 54426
rect 32726 54374 32738 54426
rect 32738 54374 32752 54426
rect 32776 54374 32790 54426
rect 32790 54374 32802 54426
rect 32802 54374 32832 54426
rect 32856 54374 32866 54426
rect 32866 54374 32912 54426
rect 32616 54372 32672 54374
rect 32696 54372 32752 54374
rect 32776 54372 32832 54374
rect 32856 54372 32912 54374
rect 32616 53338 32672 53340
rect 32696 53338 32752 53340
rect 32776 53338 32832 53340
rect 32856 53338 32912 53340
rect 32616 53286 32662 53338
rect 32662 53286 32672 53338
rect 32696 53286 32726 53338
rect 32726 53286 32738 53338
rect 32738 53286 32752 53338
rect 32776 53286 32790 53338
rect 32790 53286 32802 53338
rect 32802 53286 32832 53338
rect 32856 53286 32866 53338
rect 32866 53286 32912 53338
rect 32616 53284 32672 53286
rect 32696 53284 32752 53286
rect 32776 53284 32832 53286
rect 32856 53284 32912 53286
rect 36956 69114 37012 69116
rect 37036 69114 37092 69116
rect 37116 69114 37172 69116
rect 37196 69114 37252 69116
rect 36956 69062 37002 69114
rect 37002 69062 37012 69114
rect 37036 69062 37066 69114
rect 37066 69062 37078 69114
rect 37078 69062 37092 69114
rect 37116 69062 37130 69114
rect 37130 69062 37142 69114
rect 37142 69062 37172 69114
rect 37196 69062 37206 69114
rect 37206 69062 37252 69114
rect 36956 69060 37012 69062
rect 37036 69060 37092 69062
rect 37116 69060 37172 69062
rect 37196 69060 37252 69062
rect 33230 58284 33232 58304
rect 33232 58284 33284 58304
rect 33284 58284 33286 58304
rect 33230 58248 33286 58284
rect 33506 55664 33562 55720
rect 32616 52250 32672 52252
rect 32696 52250 32752 52252
rect 32776 52250 32832 52252
rect 32856 52250 32912 52252
rect 32616 52198 32662 52250
rect 32662 52198 32672 52250
rect 32696 52198 32726 52250
rect 32726 52198 32738 52250
rect 32738 52198 32752 52250
rect 32776 52198 32790 52250
rect 32790 52198 32802 52250
rect 32802 52198 32832 52250
rect 32856 52198 32866 52250
rect 32866 52198 32912 52250
rect 32616 52196 32672 52198
rect 32696 52196 32752 52198
rect 32776 52196 32832 52198
rect 32856 52196 32912 52198
rect 32616 51162 32672 51164
rect 32696 51162 32752 51164
rect 32776 51162 32832 51164
rect 32856 51162 32912 51164
rect 32616 51110 32662 51162
rect 32662 51110 32672 51162
rect 32696 51110 32726 51162
rect 32726 51110 32738 51162
rect 32738 51110 32752 51162
rect 32776 51110 32790 51162
rect 32790 51110 32802 51162
rect 32802 51110 32832 51162
rect 32856 51110 32866 51162
rect 32866 51110 32912 51162
rect 32616 51108 32672 51110
rect 32696 51108 32752 51110
rect 32776 51108 32832 51110
rect 32856 51108 32912 51110
rect 32616 50074 32672 50076
rect 32696 50074 32752 50076
rect 32776 50074 32832 50076
rect 32856 50074 32912 50076
rect 32616 50022 32662 50074
rect 32662 50022 32672 50074
rect 32696 50022 32726 50074
rect 32726 50022 32738 50074
rect 32738 50022 32752 50074
rect 32776 50022 32790 50074
rect 32790 50022 32802 50074
rect 32802 50022 32832 50074
rect 32856 50022 32866 50074
rect 32866 50022 32912 50074
rect 32616 50020 32672 50022
rect 32696 50020 32752 50022
rect 32776 50020 32832 50022
rect 32856 50020 32912 50022
rect 32616 48986 32672 48988
rect 32696 48986 32752 48988
rect 32776 48986 32832 48988
rect 32856 48986 32912 48988
rect 32616 48934 32662 48986
rect 32662 48934 32672 48986
rect 32696 48934 32726 48986
rect 32726 48934 32738 48986
rect 32738 48934 32752 48986
rect 32776 48934 32790 48986
rect 32790 48934 32802 48986
rect 32802 48934 32832 48986
rect 32856 48934 32866 48986
rect 32866 48934 32912 48986
rect 32616 48932 32672 48934
rect 32696 48932 32752 48934
rect 32776 48932 32832 48934
rect 32856 48932 32912 48934
rect 32616 47898 32672 47900
rect 32696 47898 32752 47900
rect 32776 47898 32832 47900
rect 32856 47898 32912 47900
rect 32616 47846 32662 47898
rect 32662 47846 32672 47898
rect 32696 47846 32726 47898
rect 32726 47846 32738 47898
rect 32738 47846 32752 47898
rect 32776 47846 32790 47898
rect 32790 47846 32802 47898
rect 32802 47846 32832 47898
rect 32856 47846 32866 47898
rect 32866 47846 32912 47898
rect 32616 47844 32672 47846
rect 32696 47844 32752 47846
rect 32776 47844 32832 47846
rect 32856 47844 32912 47846
rect 33138 51212 33140 51232
rect 33140 51212 33192 51232
rect 33192 51212 33194 51232
rect 33138 51176 33194 51212
rect 32616 46810 32672 46812
rect 32696 46810 32752 46812
rect 32776 46810 32832 46812
rect 32856 46810 32912 46812
rect 32616 46758 32662 46810
rect 32662 46758 32672 46810
rect 32696 46758 32726 46810
rect 32726 46758 32738 46810
rect 32738 46758 32752 46810
rect 32776 46758 32790 46810
rect 32790 46758 32802 46810
rect 32802 46758 32832 46810
rect 32856 46758 32866 46810
rect 32866 46758 32912 46810
rect 32616 46756 32672 46758
rect 32696 46756 32752 46758
rect 32776 46756 32832 46758
rect 32856 46756 32912 46758
rect 32616 45722 32672 45724
rect 32696 45722 32752 45724
rect 32776 45722 32832 45724
rect 32856 45722 32912 45724
rect 32616 45670 32662 45722
rect 32662 45670 32672 45722
rect 32696 45670 32726 45722
rect 32726 45670 32738 45722
rect 32738 45670 32752 45722
rect 32776 45670 32790 45722
rect 32790 45670 32802 45722
rect 32802 45670 32832 45722
rect 32856 45670 32866 45722
rect 32866 45670 32912 45722
rect 32616 45668 32672 45670
rect 32696 45668 32752 45670
rect 32776 45668 32832 45670
rect 32856 45668 32912 45670
rect 32616 44634 32672 44636
rect 32696 44634 32752 44636
rect 32776 44634 32832 44636
rect 32856 44634 32912 44636
rect 32616 44582 32662 44634
rect 32662 44582 32672 44634
rect 32696 44582 32726 44634
rect 32726 44582 32738 44634
rect 32738 44582 32752 44634
rect 32776 44582 32790 44634
rect 32790 44582 32802 44634
rect 32802 44582 32832 44634
rect 32856 44582 32866 44634
rect 32866 44582 32912 44634
rect 32616 44580 32672 44582
rect 32696 44580 32752 44582
rect 32776 44580 32832 44582
rect 32856 44580 32912 44582
rect 32616 43546 32672 43548
rect 32696 43546 32752 43548
rect 32776 43546 32832 43548
rect 32856 43546 32912 43548
rect 32616 43494 32662 43546
rect 32662 43494 32672 43546
rect 32696 43494 32726 43546
rect 32726 43494 32738 43546
rect 32738 43494 32752 43546
rect 32776 43494 32790 43546
rect 32790 43494 32802 43546
rect 32802 43494 32832 43546
rect 32856 43494 32866 43546
rect 32866 43494 32912 43546
rect 32616 43492 32672 43494
rect 32696 43492 32752 43494
rect 32776 43492 32832 43494
rect 32856 43492 32912 43494
rect 32616 42458 32672 42460
rect 32696 42458 32752 42460
rect 32776 42458 32832 42460
rect 32856 42458 32912 42460
rect 32616 42406 32662 42458
rect 32662 42406 32672 42458
rect 32696 42406 32726 42458
rect 32726 42406 32738 42458
rect 32738 42406 32752 42458
rect 32776 42406 32790 42458
rect 32790 42406 32802 42458
rect 32802 42406 32832 42458
rect 32856 42406 32866 42458
rect 32866 42406 32912 42458
rect 32616 42404 32672 42406
rect 32696 42404 32752 42406
rect 32776 42404 32832 42406
rect 32856 42404 32912 42406
rect 32616 41370 32672 41372
rect 32696 41370 32752 41372
rect 32776 41370 32832 41372
rect 32856 41370 32912 41372
rect 32616 41318 32662 41370
rect 32662 41318 32672 41370
rect 32696 41318 32726 41370
rect 32726 41318 32738 41370
rect 32738 41318 32752 41370
rect 32776 41318 32790 41370
rect 32790 41318 32802 41370
rect 32802 41318 32832 41370
rect 32856 41318 32866 41370
rect 32866 41318 32912 41370
rect 32616 41316 32672 41318
rect 32696 41316 32752 41318
rect 32776 41316 32832 41318
rect 32856 41316 32912 41318
rect 32616 40282 32672 40284
rect 32696 40282 32752 40284
rect 32776 40282 32832 40284
rect 32856 40282 32912 40284
rect 32616 40230 32662 40282
rect 32662 40230 32672 40282
rect 32696 40230 32726 40282
rect 32726 40230 32738 40282
rect 32738 40230 32752 40282
rect 32776 40230 32790 40282
rect 32790 40230 32802 40282
rect 32802 40230 32832 40282
rect 32856 40230 32866 40282
rect 32866 40230 32912 40282
rect 32616 40228 32672 40230
rect 32696 40228 32752 40230
rect 32776 40228 32832 40230
rect 32856 40228 32912 40230
rect 32616 39194 32672 39196
rect 32696 39194 32752 39196
rect 32776 39194 32832 39196
rect 32856 39194 32912 39196
rect 32616 39142 32662 39194
rect 32662 39142 32672 39194
rect 32696 39142 32726 39194
rect 32726 39142 32738 39194
rect 32738 39142 32752 39194
rect 32776 39142 32790 39194
rect 32790 39142 32802 39194
rect 32802 39142 32832 39194
rect 32856 39142 32866 39194
rect 32866 39142 32912 39194
rect 32616 39140 32672 39142
rect 32696 39140 32752 39142
rect 32776 39140 32832 39142
rect 32856 39140 32912 39142
rect 32616 38106 32672 38108
rect 32696 38106 32752 38108
rect 32776 38106 32832 38108
rect 32856 38106 32912 38108
rect 32616 38054 32662 38106
rect 32662 38054 32672 38106
rect 32696 38054 32726 38106
rect 32726 38054 32738 38106
rect 32738 38054 32752 38106
rect 32776 38054 32790 38106
rect 32790 38054 32802 38106
rect 32802 38054 32832 38106
rect 32856 38054 32866 38106
rect 32866 38054 32912 38106
rect 32616 38052 32672 38054
rect 32696 38052 32752 38054
rect 32776 38052 32832 38054
rect 32856 38052 32912 38054
rect 32616 37018 32672 37020
rect 32696 37018 32752 37020
rect 32776 37018 32832 37020
rect 32856 37018 32912 37020
rect 32616 36966 32662 37018
rect 32662 36966 32672 37018
rect 32696 36966 32726 37018
rect 32726 36966 32738 37018
rect 32738 36966 32752 37018
rect 32776 36966 32790 37018
rect 32790 36966 32802 37018
rect 32802 36966 32832 37018
rect 32856 36966 32866 37018
rect 32866 36966 32912 37018
rect 32616 36964 32672 36966
rect 32696 36964 32752 36966
rect 32776 36964 32832 36966
rect 32856 36964 32912 36966
rect 32616 35930 32672 35932
rect 32696 35930 32752 35932
rect 32776 35930 32832 35932
rect 32856 35930 32912 35932
rect 32616 35878 32662 35930
rect 32662 35878 32672 35930
rect 32696 35878 32726 35930
rect 32726 35878 32738 35930
rect 32738 35878 32752 35930
rect 32776 35878 32790 35930
rect 32790 35878 32802 35930
rect 32802 35878 32832 35930
rect 32856 35878 32866 35930
rect 32866 35878 32912 35930
rect 32616 35876 32672 35878
rect 32696 35876 32752 35878
rect 32776 35876 32832 35878
rect 32856 35876 32912 35878
rect 32616 34842 32672 34844
rect 32696 34842 32752 34844
rect 32776 34842 32832 34844
rect 32856 34842 32912 34844
rect 32616 34790 32662 34842
rect 32662 34790 32672 34842
rect 32696 34790 32726 34842
rect 32726 34790 32738 34842
rect 32738 34790 32752 34842
rect 32776 34790 32790 34842
rect 32790 34790 32802 34842
rect 32802 34790 32832 34842
rect 32856 34790 32866 34842
rect 32866 34790 32912 34842
rect 32616 34788 32672 34790
rect 32696 34788 32752 34790
rect 32776 34788 32832 34790
rect 32856 34788 32912 34790
rect 32616 33754 32672 33756
rect 32696 33754 32752 33756
rect 32776 33754 32832 33756
rect 32856 33754 32912 33756
rect 32616 33702 32662 33754
rect 32662 33702 32672 33754
rect 32696 33702 32726 33754
rect 32726 33702 32738 33754
rect 32738 33702 32752 33754
rect 32776 33702 32790 33754
rect 32790 33702 32802 33754
rect 32802 33702 32832 33754
rect 32856 33702 32866 33754
rect 32866 33702 32912 33754
rect 32616 33700 32672 33702
rect 32696 33700 32752 33702
rect 32776 33700 32832 33702
rect 32856 33700 32912 33702
rect 32616 32666 32672 32668
rect 32696 32666 32752 32668
rect 32776 32666 32832 32668
rect 32856 32666 32912 32668
rect 32616 32614 32662 32666
rect 32662 32614 32672 32666
rect 32696 32614 32726 32666
rect 32726 32614 32738 32666
rect 32738 32614 32752 32666
rect 32776 32614 32790 32666
rect 32790 32614 32802 32666
rect 32802 32614 32832 32666
rect 32856 32614 32866 32666
rect 32866 32614 32912 32666
rect 32616 32612 32672 32614
rect 32696 32612 32752 32614
rect 32776 32612 32832 32614
rect 32856 32612 32912 32614
rect 32616 31578 32672 31580
rect 32696 31578 32752 31580
rect 32776 31578 32832 31580
rect 32856 31578 32912 31580
rect 32616 31526 32662 31578
rect 32662 31526 32672 31578
rect 32696 31526 32726 31578
rect 32726 31526 32738 31578
rect 32738 31526 32752 31578
rect 32776 31526 32790 31578
rect 32790 31526 32802 31578
rect 32802 31526 32832 31578
rect 32856 31526 32866 31578
rect 32866 31526 32912 31578
rect 32616 31524 32672 31526
rect 32696 31524 32752 31526
rect 32776 31524 32832 31526
rect 32856 31524 32912 31526
rect 32616 30490 32672 30492
rect 32696 30490 32752 30492
rect 32776 30490 32832 30492
rect 32856 30490 32912 30492
rect 32616 30438 32662 30490
rect 32662 30438 32672 30490
rect 32696 30438 32726 30490
rect 32726 30438 32738 30490
rect 32738 30438 32752 30490
rect 32776 30438 32790 30490
rect 32790 30438 32802 30490
rect 32802 30438 32832 30490
rect 32856 30438 32866 30490
rect 32866 30438 32912 30490
rect 32616 30436 32672 30438
rect 32696 30436 32752 30438
rect 32776 30436 32832 30438
rect 32856 30436 32912 30438
rect 32616 29402 32672 29404
rect 32696 29402 32752 29404
rect 32776 29402 32832 29404
rect 32856 29402 32912 29404
rect 32616 29350 32662 29402
rect 32662 29350 32672 29402
rect 32696 29350 32726 29402
rect 32726 29350 32738 29402
rect 32738 29350 32752 29402
rect 32776 29350 32790 29402
rect 32790 29350 32802 29402
rect 32802 29350 32832 29402
rect 32856 29350 32866 29402
rect 32866 29350 32912 29402
rect 32616 29348 32672 29350
rect 32696 29348 32752 29350
rect 32776 29348 32832 29350
rect 32856 29348 32912 29350
rect 32616 28314 32672 28316
rect 32696 28314 32752 28316
rect 32776 28314 32832 28316
rect 32856 28314 32912 28316
rect 32616 28262 32662 28314
rect 32662 28262 32672 28314
rect 32696 28262 32726 28314
rect 32726 28262 32738 28314
rect 32738 28262 32752 28314
rect 32776 28262 32790 28314
rect 32790 28262 32802 28314
rect 32802 28262 32832 28314
rect 32856 28262 32866 28314
rect 32866 28262 32912 28314
rect 32616 28260 32672 28262
rect 32696 28260 32752 28262
rect 32776 28260 32832 28262
rect 32856 28260 32912 28262
rect 32616 27226 32672 27228
rect 32696 27226 32752 27228
rect 32776 27226 32832 27228
rect 32856 27226 32912 27228
rect 32616 27174 32662 27226
rect 32662 27174 32672 27226
rect 32696 27174 32726 27226
rect 32726 27174 32738 27226
rect 32738 27174 32752 27226
rect 32776 27174 32790 27226
rect 32790 27174 32802 27226
rect 32802 27174 32832 27226
rect 32856 27174 32866 27226
rect 32866 27174 32912 27226
rect 32616 27172 32672 27174
rect 32696 27172 32752 27174
rect 32776 27172 32832 27174
rect 32856 27172 32912 27174
rect 32616 26138 32672 26140
rect 32696 26138 32752 26140
rect 32776 26138 32832 26140
rect 32856 26138 32912 26140
rect 32616 26086 32662 26138
rect 32662 26086 32672 26138
rect 32696 26086 32726 26138
rect 32726 26086 32738 26138
rect 32738 26086 32752 26138
rect 32776 26086 32790 26138
rect 32790 26086 32802 26138
rect 32802 26086 32832 26138
rect 32856 26086 32866 26138
rect 32866 26086 32912 26138
rect 32616 26084 32672 26086
rect 32696 26084 32752 26086
rect 32776 26084 32832 26086
rect 32856 26084 32912 26086
rect 31956 25594 32012 25596
rect 32036 25594 32092 25596
rect 32116 25594 32172 25596
rect 32196 25594 32252 25596
rect 31956 25542 32002 25594
rect 32002 25542 32012 25594
rect 32036 25542 32066 25594
rect 32066 25542 32078 25594
rect 32078 25542 32092 25594
rect 32116 25542 32130 25594
rect 32130 25542 32142 25594
rect 32142 25542 32172 25594
rect 32196 25542 32206 25594
rect 32206 25542 32252 25594
rect 31956 25540 32012 25542
rect 32036 25540 32092 25542
rect 32116 25540 32172 25542
rect 32196 25540 32252 25542
rect 32616 25050 32672 25052
rect 32696 25050 32752 25052
rect 32776 25050 32832 25052
rect 32856 25050 32912 25052
rect 32616 24998 32662 25050
rect 32662 24998 32672 25050
rect 32696 24998 32726 25050
rect 32726 24998 32738 25050
rect 32738 24998 32752 25050
rect 32776 24998 32790 25050
rect 32790 24998 32802 25050
rect 32802 24998 32832 25050
rect 32856 24998 32866 25050
rect 32866 24998 32912 25050
rect 32616 24996 32672 24998
rect 32696 24996 32752 24998
rect 32776 24996 32832 24998
rect 32856 24996 32912 24998
rect 31956 24506 32012 24508
rect 32036 24506 32092 24508
rect 32116 24506 32172 24508
rect 32196 24506 32252 24508
rect 31956 24454 32002 24506
rect 32002 24454 32012 24506
rect 32036 24454 32066 24506
rect 32066 24454 32078 24506
rect 32078 24454 32092 24506
rect 32116 24454 32130 24506
rect 32130 24454 32142 24506
rect 32142 24454 32172 24506
rect 32196 24454 32206 24506
rect 32206 24454 32252 24506
rect 31956 24452 32012 24454
rect 32036 24452 32092 24454
rect 32116 24452 32172 24454
rect 32196 24452 32252 24454
rect 32616 23962 32672 23964
rect 32696 23962 32752 23964
rect 32776 23962 32832 23964
rect 32856 23962 32912 23964
rect 32616 23910 32662 23962
rect 32662 23910 32672 23962
rect 32696 23910 32726 23962
rect 32726 23910 32738 23962
rect 32738 23910 32752 23962
rect 32776 23910 32790 23962
rect 32790 23910 32802 23962
rect 32802 23910 32832 23962
rect 32856 23910 32866 23962
rect 32866 23910 32912 23962
rect 32616 23908 32672 23910
rect 32696 23908 32752 23910
rect 32776 23908 32832 23910
rect 32856 23908 32912 23910
rect 31956 23418 32012 23420
rect 32036 23418 32092 23420
rect 32116 23418 32172 23420
rect 32196 23418 32252 23420
rect 31956 23366 32002 23418
rect 32002 23366 32012 23418
rect 32036 23366 32066 23418
rect 32066 23366 32078 23418
rect 32078 23366 32092 23418
rect 32116 23366 32130 23418
rect 32130 23366 32142 23418
rect 32142 23366 32172 23418
rect 32196 23366 32206 23418
rect 32206 23366 32252 23418
rect 31956 23364 32012 23366
rect 32036 23364 32092 23366
rect 32116 23364 32172 23366
rect 32196 23364 32252 23366
rect 32616 22874 32672 22876
rect 32696 22874 32752 22876
rect 32776 22874 32832 22876
rect 32856 22874 32912 22876
rect 32616 22822 32662 22874
rect 32662 22822 32672 22874
rect 32696 22822 32726 22874
rect 32726 22822 32738 22874
rect 32738 22822 32752 22874
rect 32776 22822 32790 22874
rect 32790 22822 32802 22874
rect 32802 22822 32832 22874
rect 32856 22822 32866 22874
rect 32866 22822 32912 22874
rect 32616 22820 32672 22822
rect 32696 22820 32752 22822
rect 32776 22820 32832 22822
rect 32856 22820 32912 22822
rect 31956 22330 32012 22332
rect 32036 22330 32092 22332
rect 32116 22330 32172 22332
rect 32196 22330 32252 22332
rect 31956 22278 32002 22330
rect 32002 22278 32012 22330
rect 32036 22278 32066 22330
rect 32066 22278 32078 22330
rect 32078 22278 32092 22330
rect 32116 22278 32130 22330
rect 32130 22278 32142 22330
rect 32142 22278 32172 22330
rect 32196 22278 32206 22330
rect 32206 22278 32252 22330
rect 31956 22276 32012 22278
rect 32036 22276 32092 22278
rect 32116 22276 32172 22278
rect 32196 22276 32252 22278
rect 32616 21786 32672 21788
rect 32696 21786 32752 21788
rect 32776 21786 32832 21788
rect 32856 21786 32912 21788
rect 32616 21734 32662 21786
rect 32662 21734 32672 21786
rect 32696 21734 32726 21786
rect 32726 21734 32738 21786
rect 32738 21734 32752 21786
rect 32776 21734 32790 21786
rect 32790 21734 32802 21786
rect 32802 21734 32832 21786
rect 32856 21734 32866 21786
rect 32866 21734 32912 21786
rect 32616 21732 32672 21734
rect 32696 21732 32752 21734
rect 32776 21732 32832 21734
rect 32856 21732 32912 21734
rect 31956 21242 32012 21244
rect 32036 21242 32092 21244
rect 32116 21242 32172 21244
rect 32196 21242 32252 21244
rect 31956 21190 32002 21242
rect 32002 21190 32012 21242
rect 32036 21190 32066 21242
rect 32066 21190 32078 21242
rect 32078 21190 32092 21242
rect 32116 21190 32130 21242
rect 32130 21190 32142 21242
rect 32142 21190 32172 21242
rect 32196 21190 32206 21242
rect 32206 21190 32252 21242
rect 31956 21188 32012 21190
rect 32036 21188 32092 21190
rect 32116 21188 32172 21190
rect 32196 21188 32252 21190
rect 31956 20154 32012 20156
rect 32036 20154 32092 20156
rect 32116 20154 32172 20156
rect 32196 20154 32252 20156
rect 31956 20102 32002 20154
rect 32002 20102 32012 20154
rect 32036 20102 32066 20154
rect 32066 20102 32078 20154
rect 32078 20102 32092 20154
rect 32116 20102 32130 20154
rect 32130 20102 32142 20154
rect 32142 20102 32172 20154
rect 32196 20102 32206 20154
rect 32206 20102 32252 20154
rect 31956 20100 32012 20102
rect 32036 20100 32092 20102
rect 32116 20100 32172 20102
rect 32196 20100 32252 20102
rect 31956 19066 32012 19068
rect 32036 19066 32092 19068
rect 32116 19066 32172 19068
rect 32196 19066 32252 19068
rect 31956 19014 32002 19066
rect 32002 19014 32012 19066
rect 32036 19014 32066 19066
rect 32066 19014 32078 19066
rect 32078 19014 32092 19066
rect 32116 19014 32130 19066
rect 32130 19014 32142 19066
rect 32142 19014 32172 19066
rect 32196 19014 32206 19066
rect 32206 19014 32252 19066
rect 31956 19012 32012 19014
rect 32036 19012 32092 19014
rect 32116 19012 32172 19014
rect 32196 19012 32252 19014
rect 31956 17978 32012 17980
rect 32036 17978 32092 17980
rect 32116 17978 32172 17980
rect 32196 17978 32252 17980
rect 31956 17926 32002 17978
rect 32002 17926 32012 17978
rect 32036 17926 32066 17978
rect 32066 17926 32078 17978
rect 32078 17926 32092 17978
rect 32116 17926 32130 17978
rect 32130 17926 32142 17978
rect 32142 17926 32172 17978
rect 32196 17926 32206 17978
rect 32206 17926 32252 17978
rect 31956 17924 32012 17926
rect 32036 17924 32092 17926
rect 32116 17924 32172 17926
rect 32196 17924 32252 17926
rect 31956 16890 32012 16892
rect 32036 16890 32092 16892
rect 32116 16890 32172 16892
rect 32196 16890 32252 16892
rect 31956 16838 32002 16890
rect 32002 16838 32012 16890
rect 32036 16838 32066 16890
rect 32066 16838 32078 16890
rect 32078 16838 32092 16890
rect 32116 16838 32130 16890
rect 32130 16838 32142 16890
rect 32142 16838 32172 16890
rect 32196 16838 32206 16890
rect 32206 16838 32252 16890
rect 31956 16836 32012 16838
rect 32036 16836 32092 16838
rect 32116 16836 32172 16838
rect 32196 16836 32252 16838
rect 31956 15802 32012 15804
rect 32036 15802 32092 15804
rect 32116 15802 32172 15804
rect 32196 15802 32252 15804
rect 31956 15750 32002 15802
rect 32002 15750 32012 15802
rect 32036 15750 32066 15802
rect 32066 15750 32078 15802
rect 32078 15750 32092 15802
rect 32116 15750 32130 15802
rect 32130 15750 32142 15802
rect 32142 15750 32172 15802
rect 32196 15750 32206 15802
rect 32206 15750 32252 15802
rect 31956 15748 32012 15750
rect 32036 15748 32092 15750
rect 32116 15748 32172 15750
rect 32196 15748 32252 15750
rect 32616 20698 32672 20700
rect 32696 20698 32752 20700
rect 32776 20698 32832 20700
rect 32856 20698 32912 20700
rect 32616 20646 32662 20698
rect 32662 20646 32672 20698
rect 32696 20646 32726 20698
rect 32726 20646 32738 20698
rect 32738 20646 32752 20698
rect 32776 20646 32790 20698
rect 32790 20646 32802 20698
rect 32802 20646 32832 20698
rect 32856 20646 32866 20698
rect 32866 20646 32912 20698
rect 32616 20644 32672 20646
rect 32696 20644 32752 20646
rect 32776 20644 32832 20646
rect 32856 20644 32912 20646
rect 32616 19610 32672 19612
rect 32696 19610 32752 19612
rect 32776 19610 32832 19612
rect 32856 19610 32912 19612
rect 32616 19558 32662 19610
rect 32662 19558 32672 19610
rect 32696 19558 32726 19610
rect 32726 19558 32738 19610
rect 32738 19558 32752 19610
rect 32776 19558 32790 19610
rect 32790 19558 32802 19610
rect 32802 19558 32832 19610
rect 32856 19558 32866 19610
rect 32866 19558 32912 19610
rect 32616 19556 32672 19558
rect 32696 19556 32752 19558
rect 32776 19556 32832 19558
rect 32856 19556 32912 19558
rect 32616 18522 32672 18524
rect 32696 18522 32752 18524
rect 32776 18522 32832 18524
rect 32856 18522 32912 18524
rect 32616 18470 32662 18522
rect 32662 18470 32672 18522
rect 32696 18470 32726 18522
rect 32726 18470 32738 18522
rect 32738 18470 32752 18522
rect 32776 18470 32790 18522
rect 32790 18470 32802 18522
rect 32802 18470 32832 18522
rect 32856 18470 32866 18522
rect 32866 18470 32912 18522
rect 32616 18468 32672 18470
rect 32696 18468 32752 18470
rect 32776 18468 32832 18470
rect 32856 18468 32912 18470
rect 32616 17434 32672 17436
rect 32696 17434 32752 17436
rect 32776 17434 32832 17436
rect 32856 17434 32912 17436
rect 32616 17382 32662 17434
rect 32662 17382 32672 17434
rect 32696 17382 32726 17434
rect 32726 17382 32738 17434
rect 32738 17382 32752 17434
rect 32776 17382 32790 17434
rect 32790 17382 32802 17434
rect 32802 17382 32832 17434
rect 32856 17382 32866 17434
rect 32866 17382 32912 17434
rect 32616 17380 32672 17382
rect 32696 17380 32752 17382
rect 32776 17380 32832 17382
rect 32856 17380 32912 17382
rect 32616 16346 32672 16348
rect 32696 16346 32752 16348
rect 32776 16346 32832 16348
rect 32856 16346 32912 16348
rect 32616 16294 32662 16346
rect 32662 16294 32672 16346
rect 32696 16294 32726 16346
rect 32726 16294 32738 16346
rect 32738 16294 32752 16346
rect 32776 16294 32790 16346
rect 32790 16294 32802 16346
rect 32802 16294 32832 16346
rect 32856 16294 32866 16346
rect 32866 16294 32912 16346
rect 32616 16292 32672 16294
rect 32696 16292 32752 16294
rect 32776 16292 32832 16294
rect 32856 16292 32912 16294
rect 32616 15258 32672 15260
rect 32696 15258 32752 15260
rect 32776 15258 32832 15260
rect 32856 15258 32912 15260
rect 32616 15206 32662 15258
rect 32662 15206 32672 15258
rect 32696 15206 32726 15258
rect 32726 15206 32738 15258
rect 32738 15206 32752 15258
rect 32776 15206 32790 15258
rect 32790 15206 32802 15258
rect 32802 15206 32832 15258
rect 32856 15206 32866 15258
rect 32866 15206 32912 15258
rect 32616 15204 32672 15206
rect 32696 15204 32752 15206
rect 32776 15204 32832 15206
rect 32856 15204 32912 15206
rect 31956 14714 32012 14716
rect 32036 14714 32092 14716
rect 32116 14714 32172 14716
rect 32196 14714 32252 14716
rect 31956 14662 32002 14714
rect 32002 14662 32012 14714
rect 32036 14662 32066 14714
rect 32066 14662 32078 14714
rect 32078 14662 32092 14714
rect 32116 14662 32130 14714
rect 32130 14662 32142 14714
rect 32142 14662 32172 14714
rect 32196 14662 32206 14714
rect 32206 14662 32252 14714
rect 31956 14660 32012 14662
rect 32036 14660 32092 14662
rect 32116 14660 32172 14662
rect 32196 14660 32252 14662
rect 32616 14170 32672 14172
rect 32696 14170 32752 14172
rect 32776 14170 32832 14172
rect 32856 14170 32912 14172
rect 32616 14118 32662 14170
rect 32662 14118 32672 14170
rect 32696 14118 32726 14170
rect 32726 14118 32738 14170
rect 32738 14118 32752 14170
rect 32776 14118 32790 14170
rect 32790 14118 32802 14170
rect 32802 14118 32832 14170
rect 32856 14118 32866 14170
rect 32866 14118 32912 14170
rect 32616 14116 32672 14118
rect 32696 14116 32752 14118
rect 32776 14116 32832 14118
rect 32856 14116 32912 14118
rect 31956 13626 32012 13628
rect 32036 13626 32092 13628
rect 32116 13626 32172 13628
rect 32196 13626 32252 13628
rect 31956 13574 32002 13626
rect 32002 13574 32012 13626
rect 32036 13574 32066 13626
rect 32066 13574 32078 13626
rect 32078 13574 32092 13626
rect 32116 13574 32130 13626
rect 32130 13574 32142 13626
rect 32142 13574 32172 13626
rect 32196 13574 32206 13626
rect 32206 13574 32252 13626
rect 31956 13572 32012 13574
rect 32036 13572 32092 13574
rect 32116 13572 32172 13574
rect 32196 13572 32252 13574
rect 32616 13082 32672 13084
rect 32696 13082 32752 13084
rect 32776 13082 32832 13084
rect 32856 13082 32912 13084
rect 32616 13030 32662 13082
rect 32662 13030 32672 13082
rect 32696 13030 32726 13082
rect 32726 13030 32738 13082
rect 32738 13030 32752 13082
rect 32776 13030 32790 13082
rect 32790 13030 32802 13082
rect 32802 13030 32832 13082
rect 32856 13030 32866 13082
rect 32866 13030 32912 13082
rect 32616 13028 32672 13030
rect 32696 13028 32752 13030
rect 32776 13028 32832 13030
rect 32856 13028 32912 13030
rect 31956 12538 32012 12540
rect 32036 12538 32092 12540
rect 32116 12538 32172 12540
rect 32196 12538 32252 12540
rect 31956 12486 32002 12538
rect 32002 12486 32012 12538
rect 32036 12486 32066 12538
rect 32066 12486 32078 12538
rect 32078 12486 32092 12538
rect 32116 12486 32130 12538
rect 32130 12486 32142 12538
rect 32142 12486 32172 12538
rect 32196 12486 32206 12538
rect 32206 12486 32252 12538
rect 31956 12484 32012 12486
rect 32036 12484 32092 12486
rect 32116 12484 32172 12486
rect 32196 12484 32252 12486
rect 32616 11994 32672 11996
rect 32696 11994 32752 11996
rect 32776 11994 32832 11996
rect 32856 11994 32912 11996
rect 32616 11942 32662 11994
rect 32662 11942 32672 11994
rect 32696 11942 32726 11994
rect 32726 11942 32738 11994
rect 32738 11942 32752 11994
rect 32776 11942 32790 11994
rect 32790 11942 32802 11994
rect 32802 11942 32832 11994
rect 32856 11942 32866 11994
rect 32866 11942 32912 11994
rect 32616 11940 32672 11942
rect 32696 11940 32752 11942
rect 32776 11940 32832 11942
rect 32856 11940 32912 11942
rect 31956 11450 32012 11452
rect 32036 11450 32092 11452
rect 32116 11450 32172 11452
rect 32196 11450 32252 11452
rect 31956 11398 32002 11450
rect 32002 11398 32012 11450
rect 32036 11398 32066 11450
rect 32066 11398 32078 11450
rect 32078 11398 32092 11450
rect 32116 11398 32130 11450
rect 32130 11398 32142 11450
rect 32142 11398 32172 11450
rect 32196 11398 32206 11450
rect 32206 11398 32252 11450
rect 31956 11396 32012 11398
rect 32036 11396 32092 11398
rect 32116 11396 32172 11398
rect 32196 11396 32252 11398
rect 33874 55800 33930 55856
rect 33138 10920 33194 10976
rect 32616 10906 32672 10908
rect 32696 10906 32752 10908
rect 32776 10906 32832 10908
rect 32856 10906 32912 10908
rect 32616 10854 32662 10906
rect 32662 10854 32672 10906
rect 32696 10854 32726 10906
rect 32726 10854 32738 10906
rect 32738 10854 32752 10906
rect 32776 10854 32790 10906
rect 32790 10854 32802 10906
rect 32802 10854 32832 10906
rect 32856 10854 32866 10906
rect 32866 10854 32912 10906
rect 32616 10852 32672 10854
rect 32696 10852 32752 10854
rect 32776 10852 32832 10854
rect 32856 10852 32912 10854
rect 31956 10362 32012 10364
rect 32036 10362 32092 10364
rect 32116 10362 32172 10364
rect 32196 10362 32252 10364
rect 31956 10310 32002 10362
rect 32002 10310 32012 10362
rect 32036 10310 32066 10362
rect 32066 10310 32078 10362
rect 32078 10310 32092 10362
rect 32116 10310 32130 10362
rect 32130 10310 32142 10362
rect 32142 10310 32172 10362
rect 32196 10310 32206 10362
rect 32206 10310 32252 10362
rect 31956 10308 32012 10310
rect 32036 10308 32092 10310
rect 32116 10308 32172 10310
rect 32196 10308 32252 10310
rect 32616 9818 32672 9820
rect 32696 9818 32752 9820
rect 32776 9818 32832 9820
rect 32856 9818 32912 9820
rect 32616 9766 32662 9818
rect 32662 9766 32672 9818
rect 32696 9766 32726 9818
rect 32726 9766 32738 9818
rect 32738 9766 32752 9818
rect 32776 9766 32790 9818
rect 32790 9766 32802 9818
rect 32802 9766 32832 9818
rect 32856 9766 32866 9818
rect 32866 9766 32912 9818
rect 32616 9764 32672 9766
rect 32696 9764 32752 9766
rect 32776 9764 32832 9766
rect 32856 9764 32912 9766
rect 31956 9274 32012 9276
rect 32036 9274 32092 9276
rect 32116 9274 32172 9276
rect 32196 9274 32252 9276
rect 31956 9222 32002 9274
rect 32002 9222 32012 9274
rect 32036 9222 32066 9274
rect 32066 9222 32078 9274
rect 32078 9222 32092 9274
rect 32116 9222 32130 9274
rect 32130 9222 32142 9274
rect 32142 9222 32172 9274
rect 32196 9222 32206 9274
rect 32206 9222 32252 9274
rect 31956 9220 32012 9222
rect 32036 9220 32092 9222
rect 32116 9220 32172 9222
rect 32196 9220 32252 9222
rect 36956 68026 37012 68028
rect 37036 68026 37092 68028
rect 37116 68026 37172 68028
rect 37196 68026 37252 68028
rect 36956 67974 37002 68026
rect 37002 67974 37012 68026
rect 37036 67974 37066 68026
rect 37066 67974 37078 68026
rect 37078 67974 37092 68026
rect 37116 67974 37130 68026
rect 37130 67974 37142 68026
rect 37142 67974 37172 68026
rect 37196 67974 37206 68026
rect 37206 67974 37252 68026
rect 36956 67972 37012 67974
rect 37036 67972 37092 67974
rect 37116 67972 37172 67974
rect 37196 67972 37252 67974
rect 36956 66938 37012 66940
rect 37036 66938 37092 66940
rect 37116 66938 37172 66940
rect 37196 66938 37252 66940
rect 36956 66886 37002 66938
rect 37002 66886 37012 66938
rect 37036 66886 37066 66938
rect 37066 66886 37078 66938
rect 37078 66886 37092 66938
rect 37116 66886 37130 66938
rect 37130 66886 37142 66938
rect 37142 66886 37172 66938
rect 37196 66886 37206 66938
rect 37206 66886 37252 66938
rect 36956 66884 37012 66886
rect 37036 66884 37092 66886
rect 37116 66884 37172 66886
rect 37196 66884 37252 66886
rect 36956 65850 37012 65852
rect 37036 65850 37092 65852
rect 37116 65850 37172 65852
rect 37196 65850 37252 65852
rect 36956 65798 37002 65850
rect 37002 65798 37012 65850
rect 37036 65798 37066 65850
rect 37066 65798 37078 65850
rect 37078 65798 37092 65850
rect 37116 65798 37130 65850
rect 37130 65798 37142 65850
rect 37142 65798 37172 65850
rect 37196 65798 37206 65850
rect 37206 65798 37252 65850
rect 36956 65796 37012 65798
rect 37036 65796 37092 65798
rect 37116 65796 37172 65798
rect 37196 65796 37252 65798
rect 36956 64762 37012 64764
rect 37036 64762 37092 64764
rect 37116 64762 37172 64764
rect 37196 64762 37252 64764
rect 36956 64710 37002 64762
rect 37002 64710 37012 64762
rect 37036 64710 37066 64762
rect 37066 64710 37078 64762
rect 37078 64710 37092 64762
rect 37116 64710 37130 64762
rect 37130 64710 37142 64762
rect 37142 64710 37172 64762
rect 37196 64710 37206 64762
rect 37206 64710 37252 64762
rect 36956 64708 37012 64710
rect 37036 64708 37092 64710
rect 37116 64708 37172 64710
rect 37196 64708 37252 64710
rect 36956 63674 37012 63676
rect 37036 63674 37092 63676
rect 37116 63674 37172 63676
rect 37196 63674 37252 63676
rect 36956 63622 37002 63674
rect 37002 63622 37012 63674
rect 37036 63622 37066 63674
rect 37066 63622 37078 63674
rect 37078 63622 37092 63674
rect 37116 63622 37130 63674
rect 37130 63622 37142 63674
rect 37142 63622 37172 63674
rect 37196 63622 37206 63674
rect 37206 63622 37252 63674
rect 36956 63620 37012 63622
rect 37036 63620 37092 63622
rect 37116 63620 37172 63622
rect 37196 63620 37252 63622
rect 36956 62586 37012 62588
rect 37036 62586 37092 62588
rect 37116 62586 37172 62588
rect 37196 62586 37252 62588
rect 36956 62534 37002 62586
rect 37002 62534 37012 62586
rect 37036 62534 37066 62586
rect 37066 62534 37078 62586
rect 37078 62534 37092 62586
rect 37116 62534 37130 62586
rect 37130 62534 37142 62586
rect 37142 62534 37172 62586
rect 37196 62534 37206 62586
rect 37206 62534 37252 62586
rect 36956 62532 37012 62534
rect 37036 62532 37092 62534
rect 37116 62532 37172 62534
rect 37196 62532 37252 62534
rect 36956 61498 37012 61500
rect 37036 61498 37092 61500
rect 37116 61498 37172 61500
rect 37196 61498 37252 61500
rect 36956 61446 37002 61498
rect 37002 61446 37012 61498
rect 37036 61446 37066 61498
rect 37066 61446 37078 61498
rect 37078 61446 37092 61498
rect 37116 61446 37130 61498
rect 37130 61446 37142 61498
rect 37142 61446 37172 61498
rect 37196 61446 37206 61498
rect 37206 61446 37252 61498
rect 36956 61444 37012 61446
rect 37036 61444 37092 61446
rect 37116 61444 37172 61446
rect 37196 61444 37252 61446
rect 36956 60410 37012 60412
rect 37036 60410 37092 60412
rect 37116 60410 37172 60412
rect 37196 60410 37252 60412
rect 36956 60358 37002 60410
rect 37002 60358 37012 60410
rect 37036 60358 37066 60410
rect 37066 60358 37078 60410
rect 37078 60358 37092 60410
rect 37116 60358 37130 60410
rect 37130 60358 37142 60410
rect 37142 60358 37172 60410
rect 37196 60358 37206 60410
rect 37206 60358 37252 60410
rect 36956 60356 37012 60358
rect 37036 60356 37092 60358
rect 37116 60356 37172 60358
rect 37196 60356 37252 60358
rect 36956 59322 37012 59324
rect 37036 59322 37092 59324
rect 37116 59322 37172 59324
rect 37196 59322 37252 59324
rect 36956 59270 37002 59322
rect 37002 59270 37012 59322
rect 37036 59270 37066 59322
rect 37066 59270 37078 59322
rect 37078 59270 37092 59322
rect 37116 59270 37130 59322
rect 37130 59270 37142 59322
rect 37142 59270 37172 59322
rect 37196 59270 37206 59322
rect 37206 59270 37252 59322
rect 36956 59268 37012 59270
rect 37036 59268 37092 59270
rect 37116 59268 37172 59270
rect 37196 59268 37252 59270
rect 36956 58234 37012 58236
rect 37036 58234 37092 58236
rect 37116 58234 37172 58236
rect 37196 58234 37252 58236
rect 36956 58182 37002 58234
rect 37002 58182 37012 58234
rect 37036 58182 37066 58234
rect 37066 58182 37078 58234
rect 37078 58182 37092 58234
rect 37116 58182 37130 58234
rect 37130 58182 37142 58234
rect 37142 58182 37172 58234
rect 37196 58182 37206 58234
rect 37206 58182 37252 58234
rect 36956 58180 37012 58182
rect 37036 58180 37092 58182
rect 37116 58180 37172 58182
rect 37196 58180 37252 58182
rect 36956 57146 37012 57148
rect 37036 57146 37092 57148
rect 37116 57146 37172 57148
rect 37196 57146 37252 57148
rect 36956 57094 37002 57146
rect 37002 57094 37012 57146
rect 37036 57094 37066 57146
rect 37066 57094 37078 57146
rect 37078 57094 37092 57146
rect 37116 57094 37130 57146
rect 37130 57094 37142 57146
rect 37142 57094 37172 57146
rect 37196 57094 37206 57146
rect 37206 57094 37252 57146
rect 36956 57092 37012 57094
rect 37036 57092 37092 57094
rect 37116 57092 37172 57094
rect 37196 57092 37252 57094
rect 36956 56058 37012 56060
rect 37036 56058 37092 56060
rect 37116 56058 37172 56060
rect 37196 56058 37252 56060
rect 36956 56006 37002 56058
rect 37002 56006 37012 56058
rect 37036 56006 37066 56058
rect 37066 56006 37078 56058
rect 37078 56006 37092 56058
rect 37116 56006 37130 56058
rect 37130 56006 37142 56058
rect 37142 56006 37172 56058
rect 37196 56006 37206 56058
rect 37206 56006 37252 56058
rect 36956 56004 37012 56006
rect 37036 56004 37092 56006
rect 37116 56004 37172 56006
rect 37196 56004 37252 56006
rect 36956 54970 37012 54972
rect 37036 54970 37092 54972
rect 37116 54970 37172 54972
rect 37196 54970 37252 54972
rect 36956 54918 37002 54970
rect 37002 54918 37012 54970
rect 37036 54918 37066 54970
rect 37066 54918 37078 54970
rect 37078 54918 37092 54970
rect 37116 54918 37130 54970
rect 37130 54918 37142 54970
rect 37142 54918 37172 54970
rect 37196 54918 37206 54970
rect 37206 54918 37252 54970
rect 36956 54916 37012 54918
rect 37036 54916 37092 54918
rect 37116 54916 37172 54918
rect 37196 54916 37252 54918
rect 36956 53882 37012 53884
rect 37036 53882 37092 53884
rect 37116 53882 37172 53884
rect 37196 53882 37252 53884
rect 36956 53830 37002 53882
rect 37002 53830 37012 53882
rect 37036 53830 37066 53882
rect 37066 53830 37078 53882
rect 37078 53830 37092 53882
rect 37116 53830 37130 53882
rect 37130 53830 37142 53882
rect 37142 53830 37172 53882
rect 37196 53830 37206 53882
rect 37206 53830 37252 53882
rect 36956 53828 37012 53830
rect 37036 53828 37092 53830
rect 37116 53828 37172 53830
rect 37196 53828 37252 53830
rect 36956 52794 37012 52796
rect 37036 52794 37092 52796
rect 37116 52794 37172 52796
rect 37196 52794 37252 52796
rect 36956 52742 37002 52794
rect 37002 52742 37012 52794
rect 37036 52742 37066 52794
rect 37066 52742 37078 52794
rect 37078 52742 37092 52794
rect 37116 52742 37130 52794
rect 37130 52742 37142 52794
rect 37142 52742 37172 52794
rect 37196 52742 37206 52794
rect 37206 52742 37252 52794
rect 36956 52740 37012 52742
rect 37036 52740 37092 52742
rect 37116 52740 37172 52742
rect 37196 52740 37252 52742
rect 36956 51706 37012 51708
rect 37036 51706 37092 51708
rect 37116 51706 37172 51708
rect 37196 51706 37252 51708
rect 36956 51654 37002 51706
rect 37002 51654 37012 51706
rect 37036 51654 37066 51706
rect 37066 51654 37078 51706
rect 37078 51654 37092 51706
rect 37116 51654 37130 51706
rect 37130 51654 37142 51706
rect 37142 51654 37172 51706
rect 37196 51654 37206 51706
rect 37206 51654 37252 51706
rect 36956 51652 37012 51654
rect 37036 51652 37092 51654
rect 37116 51652 37172 51654
rect 37196 51652 37252 51654
rect 36956 50618 37012 50620
rect 37036 50618 37092 50620
rect 37116 50618 37172 50620
rect 37196 50618 37252 50620
rect 36956 50566 37002 50618
rect 37002 50566 37012 50618
rect 37036 50566 37066 50618
rect 37066 50566 37078 50618
rect 37078 50566 37092 50618
rect 37116 50566 37130 50618
rect 37130 50566 37142 50618
rect 37142 50566 37172 50618
rect 37196 50566 37206 50618
rect 37206 50566 37252 50618
rect 36956 50564 37012 50566
rect 37036 50564 37092 50566
rect 37116 50564 37172 50566
rect 37196 50564 37252 50566
rect 36956 49530 37012 49532
rect 37036 49530 37092 49532
rect 37116 49530 37172 49532
rect 37196 49530 37252 49532
rect 36956 49478 37002 49530
rect 37002 49478 37012 49530
rect 37036 49478 37066 49530
rect 37066 49478 37078 49530
rect 37078 49478 37092 49530
rect 37116 49478 37130 49530
rect 37130 49478 37142 49530
rect 37142 49478 37172 49530
rect 37196 49478 37206 49530
rect 37206 49478 37252 49530
rect 36956 49476 37012 49478
rect 37036 49476 37092 49478
rect 37116 49476 37172 49478
rect 37196 49476 37252 49478
rect 36956 48442 37012 48444
rect 37036 48442 37092 48444
rect 37116 48442 37172 48444
rect 37196 48442 37252 48444
rect 36956 48390 37002 48442
rect 37002 48390 37012 48442
rect 37036 48390 37066 48442
rect 37066 48390 37078 48442
rect 37078 48390 37092 48442
rect 37116 48390 37130 48442
rect 37130 48390 37142 48442
rect 37142 48390 37172 48442
rect 37196 48390 37206 48442
rect 37206 48390 37252 48442
rect 36956 48388 37012 48390
rect 37036 48388 37092 48390
rect 37116 48388 37172 48390
rect 37196 48388 37252 48390
rect 36956 47354 37012 47356
rect 37036 47354 37092 47356
rect 37116 47354 37172 47356
rect 37196 47354 37252 47356
rect 36956 47302 37002 47354
rect 37002 47302 37012 47354
rect 37036 47302 37066 47354
rect 37066 47302 37078 47354
rect 37078 47302 37092 47354
rect 37116 47302 37130 47354
rect 37130 47302 37142 47354
rect 37142 47302 37172 47354
rect 37196 47302 37206 47354
rect 37206 47302 37252 47354
rect 36956 47300 37012 47302
rect 37036 47300 37092 47302
rect 37116 47300 37172 47302
rect 37196 47300 37252 47302
rect 36956 46266 37012 46268
rect 37036 46266 37092 46268
rect 37116 46266 37172 46268
rect 37196 46266 37252 46268
rect 36956 46214 37002 46266
rect 37002 46214 37012 46266
rect 37036 46214 37066 46266
rect 37066 46214 37078 46266
rect 37078 46214 37092 46266
rect 37116 46214 37130 46266
rect 37130 46214 37142 46266
rect 37142 46214 37172 46266
rect 37196 46214 37206 46266
rect 37206 46214 37252 46266
rect 36956 46212 37012 46214
rect 37036 46212 37092 46214
rect 37116 46212 37172 46214
rect 37196 46212 37252 46214
rect 36956 45178 37012 45180
rect 37036 45178 37092 45180
rect 37116 45178 37172 45180
rect 37196 45178 37252 45180
rect 36956 45126 37002 45178
rect 37002 45126 37012 45178
rect 37036 45126 37066 45178
rect 37066 45126 37078 45178
rect 37078 45126 37092 45178
rect 37116 45126 37130 45178
rect 37130 45126 37142 45178
rect 37142 45126 37172 45178
rect 37196 45126 37206 45178
rect 37206 45126 37252 45178
rect 36956 45124 37012 45126
rect 37036 45124 37092 45126
rect 37116 45124 37172 45126
rect 37196 45124 37252 45126
rect 36956 44090 37012 44092
rect 37036 44090 37092 44092
rect 37116 44090 37172 44092
rect 37196 44090 37252 44092
rect 36956 44038 37002 44090
rect 37002 44038 37012 44090
rect 37036 44038 37066 44090
rect 37066 44038 37078 44090
rect 37078 44038 37092 44090
rect 37116 44038 37130 44090
rect 37130 44038 37142 44090
rect 37142 44038 37172 44090
rect 37196 44038 37206 44090
rect 37206 44038 37252 44090
rect 36956 44036 37012 44038
rect 37036 44036 37092 44038
rect 37116 44036 37172 44038
rect 37196 44036 37252 44038
rect 36956 43002 37012 43004
rect 37036 43002 37092 43004
rect 37116 43002 37172 43004
rect 37196 43002 37252 43004
rect 36956 42950 37002 43002
rect 37002 42950 37012 43002
rect 37036 42950 37066 43002
rect 37066 42950 37078 43002
rect 37078 42950 37092 43002
rect 37116 42950 37130 43002
rect 37130 42950 37142 43002
rect 37142 42950 37172 43002
rect 37196 42950 37206 43002
rect 37206 42950 37252 43002
rect 36956 42948 37012 42950
rect 37036 42948 37092 42950
rect 37116 42948 37172 42950
rect 37196 42948 37252 42950
rect 36956 41914 37012 41916
rect 37036 41914 37092 41916
rect 37116 41914 37172 41916
rect 37196 41914 37252 41916
rect 36956 41862 37002 41914
rect 37002 41862 37012 41914
rect 37036 41862 37066 41914
rect 37066 41862 37078 41914
rect 37078 41862 37092 41914
rect 37116 41862 37130 41914
rect 37130 41862 37142 41914
rect 37142 41862 37172 41914
rect 37196 41862 37206 41914
rect 37206 41862 37252 41914
rect 36956 41860 37012 41862
rect 37036 41860 37092 41862
rect 37116 41860 37172 41862
rect 37196 41860 37252 41862
rect 36956 40826 37012 40828
rect 37036 40826 37092 40828
rect 37116 40826 37172 40828
rect 37196 40826 37252 40828
rect 36956 40774 37002 40826
rect 37002 40774 37012 40826
rect 37036 40774 37066 40826
rect 37066 40774 37078 40826
rect 37078 40774 37092 40826
rect 37116 40774 37130 40826
rect 37130 40774 37142 40826
rect 37142 40774 37172 40826
rect 37196 40774 37206 40826
rect 37206 40774 37252 40826
rect 36956 40772 37012 40774
rect 37036 40772 37092 40774
rect 37116 40772 37172 40774
rect 37196 40772 37252 40774
rect 36956 39738 37012 39740
rect 37036 39738 37092 39740
rect 37116 39738 37172 39740
rect 37196 39738 37252 39740
rect 36956 39686 37002 39738
rect 37002 39686 37012 39738
rect 37036 39686 37066 39738
rect 37066 39686 37078 39738
rect 37078 39686 37092 39738
rect 37116 39686 37130 39738
rect 37130 39686 37142 39738
rect 37142 39686 37172 39738
rect 37196 39686 37206 39738
rect 37206 39686 37252 39738
rect 36956 39684 37012 39686
rect 37036 39684 37092 39686
rect 37116 39684 37172 39686
rect 37196 39684 37252 39686
rect 36956 38650 37012 38652
rect 37036 38650 37092 38652
rect 37116 38650 37172 38652
rect 37196 38650 37252 38652
rect 36956 38598 37002 38650
rect 37002 38598 37012 38650
rect 37036 38598 37066 38650
rect 37066 38598 37078 38650
rect 37078 38598 37092 38650
rect 37116 38598 37130 38650
rect 37130 38598 37142 38650
rect 37142 38598 37172 38650
rect 37196 38598 37206 38650
rect 37206 38598 37252 38650
rect 36956 38596 37012 38598
rect 37036 38596 37092 38598
rect 37116 38596 37172 38598
rect 37196 38596 37252 38598
rect 36956 37562 37012 37564
rect 37036 37562 37092 37564
rect 37116 37562 37172 37564
rect 37196 37562 37252 37564
rect 36956 37510 37002 37562
rect 37002 37510 37012 37562
rect 37036 37510 37066 37562
rect 37066 37510 37078 37562
rect 37078 37510 37092 37562
rect 37116 37510 37130 37562
rect 37130 37510 37142 37562
rect 37142 37510 37172 37562
rect 37196 37510 37206 37562
rect 37206 37510 37252 37562
rect 36956 37508 37012 37510
rect 37036 37508 37092 37510
rect 37116 37508 37172 37510
rect 37196 37508 37252 37510
rect 36956 36474 37012 36476
rect 37036 36474 37092 36476
rect 37116 36474 37172 36476
rect 37196 36474 37252 36476
rect 36956 36422 37002 36474
rect 37002 36422 37012 36474
rect 37036 36422 37066 36474
rect 37066 36422 37078 36474
rect 37078 36422 37092 36474
rect 37116 36422 37130 36474
rect 37130 36422 37142 36474
rect 37142 36422 37172 36474
rect 37196 36422 37206 36474
rect 37206 36422 37252 36474
rect 36956 36420 37012 36422
rect 37036 36420 37092 36422
rect 37116 36420 37172 36422
rect 37196 36420 37252 36422
rect 36956 35386 37012 35388
rect 37036 35386 37092 35388
rect 37116 35386 37172 35388
rect 37196 35386 37252 35388
rect 36956 35334 37002 35386
rect 37002 35334 37012 35386
rect 37036 35334 37066 35386
rect 37066 35334 37078 35386
rect 37078 35334 37092 35386
rect 37116 35334 37130 35386
rect 37130 35334 37142 35386
rect 37142 35334 37172 35386
rect 37196 35334 37206 35386
rect 37206 35334 37252 35386
rect 36956 35332 37012 35334
rect 37036 35332 37092 35334
rect 37116 35332 37172 35334
rect 37196 35332 37252 35334
rect 36956 34298 37012 34300
rect 37036 34298 37092 34300
rect 37116 34298 37172 34300
rect 37196 34298 37252 34300
rect 36956 34246 37002 34298
rect 37002 34246 37012 34298
rect 37036 34246 37066 34298
rect 37066 34246 37078 34298
rect 37078 34246 37092 34298
rect 37116 34246 37130 34298
rect 37130 34246 37142 34298
rect 37142 34246 37172 34298
rect 37196 34246 37206 34298
rect 37206 34246 37252 34298
rect 36956 34244 37012 34246
rect 37036 34244 37092 34246
rect 37116 34244 37172 34246
rect 37196 34244 37252 34246
rect 36956 33210 37012 33212
rect 37036 33210 37092 33212
rect 37116 33210 37172 33212
rect 37196 33210 37252 33212
rect 36956 33158 37002 33210
rect 37002 33158 37012 33210
rect 37036 33158 37066 33210
rect 37066 33158 37078 33210
rect 37078 33158 37092 33210
rect 37116 33158 37130 33210
rect 37130 33158 37142 33210
rect 37142 33158 37172 33210
rect 37196 33158 37206 33210
rect 37206 33158 37252 33210
rect 36956 33156 37012 33158
rect 37036 33156 37092 33158
rect 37116 33156 37172 33158
rect 37196 33156 37252 33158
rect 36956 32122 37012 32124
rect 37036 32122 37092 32124
rect 37116 32122 37172 32124
rect 37196 32122 37252 32124
rect 36956 32070 37002 32122
rect 37002 32070 37012 32122
rect 37036 32070 37066 32122
rect 37066 32070 37078 32122
rect 37078 32070 37092 32122
rect 37116 32070 37130 32122
rect 37130 32070 37142 32122
rect 37142 32070 37172 32122
rect 37196 32070 37206 32122
rect 37206 32070 37252 32122
rect 36956 32068 37012 32070
rect 37036 32068 37092 32070
rect 37116 32068 37172 32070
rect 37196 32068 37252 32070
rect 36956 31034 37012 31036
rect 37036 31034 37092 31036
rect 37116 31034 37172 31036
rect 37196 31034 37252 31036
rect 36956 30982 37002 31034
rect 37002 30982 37012 31034
rect 37036 30982 37066 31034
rect 37066 30982 37078 31034
rect 37078 30982 37092 31034
rect 37116 30982 37130 31034
rect 37130 30982 37142 31034
rect 37142 30982 37172 31034
rect 37196 30982 37206 31034
rect 37206 30982 37252 31034
rect 36956 30980 37012 30982
rect 37036 30980 37092 30982
rect 37116 30980 37172 30982
rect 37196 30980 37252 30982
rect 36956 29946 37012 29948
rect 37036 29946 37092 29948
rect 37116 29946 37172 29948
rect 37196 29946 37252 29948
rect 36956 29894 37002 29946
rect 37002 29894 37012 29946
rect 37036 29894 37066 29946
rect 37066 29894 37078 29946
rect 37078 29894 37092 29946
rect 37116 29894 37130 29946
rect 37130 29894 37142 29946
rect 37142 29894 37172 29946
rect 37196 29894 37206 29946
rect 37206 29894 37252 29946
rect 36956 29892 37012 29894
rect 37036 29892 37092 29894
rect 37116 29892 37172 29894
rect 37196 29892 37252 29894
rect 36956 28858 37012 28860
rect 37036 28858 37092 28860
rect 37116 28858 37172 28860
rect 37196 28858 37252 28860
rect 36956 28806 37002 28858
rect 37002 28806 37012 28858
rect 37036 28806 37066 28858
rect 37066 28806 37078 28858
rect 37078 28806 37092 28858
rect 37116 28806 37130 28858
rect 37130 28806 37142 28858
rect 37142 28806 37172 28858
rect 37196 28806 37206 28858
rect 37206 28806 37252 28858
rect 36956 28804 37012 28806
rect 37036 28804 37092 28806
rect 37116 28804 37172 28806
rect 37196 28804 37252 28806
rect 36956 27770 37012 27772
rect 37036 27770 37092 27772
rect 37116 27770 37172 27772
rect 37196 27770 37252 27772
rect 36956 27718 37002 27770
rect 37002 27718 37012 27770
rect 37036 27718 37066 27770
rect 37066 27718 37078 27770
rect 37078 27718 37092 27770
rect 37116 27718 37130 27770
rect 37130 27718 37142 27770
rect 37142 27718 37172 27770
rect 37196 27718 37206 27770
rect 37206 27718 37252 27770
rect 36956 27716 37012 27718
rect 37036 27716 37092 27718
rect 37116 27716 37172 27718
rect 37196 27716 37252 27718
rect 36956 26682 37012 26684
rect 37036 26682 37092 26684
rect 37116 26682 37172 26684
rect 37196 26682 37252 26684
rect 36956 26630 37002 26682
rect 37002 26630 37012 26682
rect 37036 26630 37066 26682
rect 37066 26630 37078 26682
rect 37078 26630 37092 26682
rect 37116 26630 37130 26682
rect 37130 26630 37142 26682
rect 37142 26630 37172 26682
rect 37196 26630 37206 26682
rect 37206 26630 37252 26682
rect 36956 26628 37012 26630
rect 37036 26628 37092 26630
rect 37116 26628 37172 26630
rect 37196 26628 37252 26630
rect 36956 25594 37012 25596
rect 37036 25594 37092 25596
rect 37116 25594 37172 25596
rect 37196 25594 37252 25596
rect 36956 25542 37002 25594
rect 37002 25542 37012 25594
rect 37036 25542 37066 25594
rect 37066 25542 37078 25594
rect 37078 25542 37092 25594
rect 37116 25542 37130 25594
rect 37130 25542 37142 25594
rect 37142 25542 37172 25594
rect 37196 25542 37206 25594
rect 37206 25542 37252 25594
rect 36956 25540 37012 25542
rect 37036 25540 37092 25542
rect 37116 25540 37172 25542
rect 37196 25540 37252 25542
rect 36956 24506 37012 24508
rect 37036 24506 37092 24508
rect 37116 24506 37172 24508
rect 37196 24506 37252 24508
rect 36956 24454 37002 24506
rect 37002 24454 37012 24506
rect 37036 24454 37066 24506
rect 37066 24454 37078 24506
rect 37078 24454 37092 24506
rect 37116 24454 37130 24506
rect 37130 24454 37142 24506
rect 37142 24454 37172 24506
rect 37196 24454 37206 24506
rect 37206 24454 37252 24506
rect 36956 24452 37012 24454
rect 37036 24452 37092 24454
rect 37116 24452 37172 24454
rect 37196 24452 37252 24454
rect 36956 23418 37012 23420
rect 37036 23418 37092 23420
rect 37116 23418 37172 23420
rect 37196 23418 37252 23420
rect 36956 23366 37002 23418
rect 37002 23366 37012 23418
rect 37036 23366 37066 23418
rect 37066 23366 37078 23418
rect 37078 23366 37092 23418
rect 37116 23366 37130 23418
rect 37130 23366 37142 23418
rect 37142 23366 37172 23418
rect 37196 23366 37206 23418
rect 37206 23366 37252 23418
rect 36956 23364 37012 23366
rect 37036 23364 37092 23366
rect 37116 23364 37172 23366
rect 37196 23364 37252 23366
rect 36956 22330 37012 22332
rect 37036 22330 37092 22332
rect 37116 22330 37172 22332
rect 37196 22330 37252 22332
rect 36956 22278 37002 22330
rect 37002 22278 37012 22330
rect 37036 22278 37066 22330
rect 37066 22278 37078 22330
rect 37078 22278 37092 22330
rect 37116 22278 37130 22330
rect 37130 22278 37142 22330
rect 37142 22278 37172 22330
rect 37196 22278 37206 22330
rect 37206 22278 37252 22330
rect 36956 22276 37012 22278
rect 37036 22276 37092 22278
rect 37116 22276 37172 22278
rect 37196 22276 37252 22278
rect 37616 68570 37672 68572
rect 37696 68570 37752 68572
rect 37776 68570 37832 68572
rect 37856 68570 37912 68572
rect 37616 68518 37662 68570
rect 37662 68518 37672 68570
rect 37696 68518 37726 68570
rect 37726 68518 37738 68570
rect 37738 68518 37752 68570
rect 37776 68518 37790 68570
rect 37790 68518 37802 68570
rect 37802 68518 37832 68570
rect 37856 68518 37866 68570
rect 37866 68518 37912 68570
rect 37616 68516 37672 68518
rect 37696 68516 37752 68518
rect 37776 68516 37832 68518
rect 37856 68516 37912 68518
rect 37616 67482 37672 67484
rect 37696 67482 37752 67484
rect 37776 67482 37832 67484
rect 37856 67482 37912 67484
rect 37616 67430 37662 67482
rect 37662 67430 37672 67482
rect 37696 67430 37726 67482
rect 37726 67430 37738 67482
rect 37738 67430 37752 67482
rect 37776 67430 37790 67482
rect 37790 67430 37802 67482
rect 37802 67430 37832 67482
rect 37856 67430 37866 67482
rect 37866 67430 37912 67482
rect 37616 67428 37672 67430
rect 37696 67428 37752 67430
rect 37776 67428 37832 67430
rect 37856 67428 37912 67430
rect 37616 66394 37672 66396
rect 37696 66394 37752 66396
rect 37776 66394 37832 66396
rect 37856 66394 37912 66396
rect 37616 66342 37662 66394
rect 37662 66342 37672 66394
rect 37696 66342 37726 66394
rect 37726 66342 37738 66394
rect 37738 66342 37752 66394
rect 37776 66342 37790 66394
rect 37790 66342 37802 66394
rect 37802 66342 37832 66394
rect 37856 66342 37866 66394
rect 37866 66342 37912 66394
rect 37616 66340 37672 66342
rect 37696 66340 37752 66342
rect 37776 66340 37832 66342
rect 37856 66340 37912 66342
rect 37616 65306 37672 65308
rect 37696 65306 37752 65308
rect 37776 65306 37832 65308
rect 37856 65306 37912 65308
rect 37616 65254 37662 65306
rect 37662 65254 37672 65306
rect 37696 65254 37726 65306
rect 37726 65254 37738 65306
rect 37738 65254 37752 65306
rect 37776 65254 37790 65306
rect 37790 65254 37802 65306
rect 37802 65254 37832 65306
rect 37856 65254 37866 65306
rect 37866 65254 37912 65306
rect 37616 65252 37672 65254
rect 37696 65252 37752 65254
rect 37776 65252 37832 65254
rect 37856 65252 37912 65254
rect 37616 64218 37672 64220
rect 37696 64218 37752 64220
rect 37776 64218 37832 64220
rect 37856 64218 37912 64220
rect 37616 64166 37662 64218
rect 37662 64166 37672 64218
rect 37696 64166 37726 64218
rect 37726 64166 37738 64218
rect 37738 64166 37752 64218
rect 37776 64166 37790 64218
rect 37790 64166 37802 64218
rect 37802 64166 37832 64218
rect 37856 64166 37866 64218
rect 37866 64166 37912 64218
rect 37616 64164 37672 64166
rect 37696 64164 37752 64166
rect 37776 64164 37832 64166
rect 37856 64164 37912 64166
rect 37616 63130 37672 63132
rect 37696 63130 37752 63132
rect 37776 63130 37832 63132
rect 37856 63130 37912 63132
rect 37616 63078 37662 63130
rect 37662 63078 37672 63130
rect 37696 63078 37726 63130
rect 37726 63078 37738 63130
rect 37738 63078 37752 63130
rect 37776 63078 37790 63130
rect 37790 63078 37802 63130
rect 37802 63078 37832 63130
rect 37856 63078 37866 63130
rect 37866 63078 37912 63130
rect 37616 63076 37672 63078
rect 37696 63076 37752 63078
rect 37776 63076 37832 63078
rect 37856 63076 37912 63078
rect 37616 62042 37672 62044
rect 37696 62042 37752 62044
rect 37776 62042 37832 62044
rect 37856 62042 37912 62044
rect 37616 61990 37662 62042
rect 37662 61990 37672 62042
rect 37696 61990 37726 62042
rect 37726 61990 37738 62042
rect 37738 61990 37752 62042
rect 37776 61990 37790 62042
rect 37790 61990 37802 62042
rect 37802 61990 37832 62042
rect 37856 61990 37866 62042
rect 37866 61990 37912 62042
rect 37616 61988 37672 61990
rect 37696 61988 37752 61990
rect 37776 61988 37832 61990
rect 37856 61988 37912 61990
rect 37616 60954 37672 60956
rect 37696 60954 37752 60956
rect 37776 60954 37832 60956
rect 37856 60954 37912 60956
rect 37616 60902 37662 60954
rect 37662 60902 37672 60954
rect 37696 60902 37726 60954
rect 37726 60902 37738 60954
rect 37738 60902 37752 60954
rect 37776 60902 37790 60954
rect 37790 60902 37802 60954
rect 37802 60902 37832 60954
rect 37856 60902 37866 60954
rect 37866 60902 37912 60954
rect 37616 60900 37672 60902
rect 37696 60900 37752 60902
rect 37776 60900 37832 60902
rect 37856 60900 37912 60902
rect 37616 59866 37672 59868
rect 37696 59866 37752 59868
rect 37776 59866 37832 59868
rect 37856 59866 37912 59868
rect 37616 59814 37662 59866
rect 37662 59814 37672 59866
rect 37696 59814 37726 59866
rect 37726 59814 37738 59866
rect 37738 59814 37752 59866
rect 37776 59814 37790 59866
rect 37790 59814 37802 59866
rect 37802 59814 37832 59866
rect 37856 59814 37866 59866
rect 37866 59814 37912 59866
rect 37616 59812 37672 59814
rect 37696 59812 37752 59814
rect 37776 59812 37832 59814
rect 37856 59812 37912 59814
rect 37616 58778 37672 58780
rect 37696 58778 37752 58780
rect 37776 58778 37832 58780
rect 37856 58778 37912 58780
rect 37616 58726 37662 58778
rect 37662 58726 37672 58778
rect 37696 58726 37726 58778
rect 37726 58726 37738 58778
rect 37738 58726 37752 58778
rect 37776 58726 37790 58778
rect 37790 58726 37802 58778
rect 37802 58726 37832 58778
rect 37856 58726 37866 58778
rect 37866 58726 37912 58778
rect 37616 58724 37672 58726
rect 37696 58724 37752 58726
rect 37776 58724 37832 58726
rect 37856 58724 37912 58726
rect 37616 57690 37672 57692
rect 37696 57690 37752 57692
rect 37776 57690 37832 57692
rect 37856 57690 37912 57692
rect 37616 57638 37662 57690
rect 37662 57638 37672 57690
rect 37696 57638 37726 57690
rect 37726 57638 37738 57690
rect 37738 57638 37752 57690
rect 37776 57638 37790 57690
rect 37790 57638 37802 57690
rect 37802 57638 37832 57690
rect 37856 57638 37866 57690
rect 37866 57638 37912 57690
rect 37616 57636 37672 57638
rect 37696 57636 37752 57638
rect 37776 57636 37832 57638
rect 37856 57636 37912 57638
rect 37616 56602 37672 56604
rect 37696 56602 37752 56604
rect 37776 56602 37832 56604
rect 37856 56602 37912 56604
rect 37616 56550 37662 56602
rect 37662 56550 37672 56602
rect 37696 56550 37726 56602
rect 37726 56550 37738 56602
rect 37738 56550 37752 56602
rect 37776 56550 37790 56602
rect 37790 56550 37802 56602
rect 37802 56550 37832 56602
rect 37856 56550 37866 56602
rect 37866 56550 37912 56602
rect 37616 56548 37672 56550
rect 37696 56548 37752 56550
rect 37776 56548 37832 56550
rect 37856 56548 37912 56550
rect 37616 55514 37672 55516
rect 37696 55514 37752 55516
rect 37776 55514 37832 55516
rect 37856 55514 37912 55516
rect 37616 55462 37662 55514
rect 37662 55462 37672 55514
rect 37696 55462 37726 55514
rect 37726 55462 37738 55514
rect 37738 55462 37752 55514
rect 37776 55462 37790 55514
rect 37790 55462 37802 55514
rect 37802 55462 37832 55514
rect 37856 55462 37866 55514
rect 37866 55462 37912 55514
rect 37616 55460 37672 55462
rect 37696 55460 37752 55462
rect 37776 55460 37832 55462
rect 37856 55460 37912 55462
rect 37616 54426 37672 54428
rect 37696 54426 37752 54428
rect 37776 54426 37832 54428
rect 37856 54426 37912 54428
rect 37616 54374 37662 54426
rect 37662 54374 37672 54426
rect 37696 54374 37726 54426
rect 37726 54374 37738 54426
rect 37738 54374 37752 54426
rect 37776 54374 37790 54426
rect 37790 54374 37802 54426
rect 37802 54374 37832 54426
rect 37856 54374 37866 54426
rect 37866 54374 37912 54426
rect 37616 54372 37672 54374
rect 37696 54372 37752 54374
rect 37776 54372 37832 54374
rect 37856 54372 37912 54374
rect 37616 53338 37672 53340
rect 37696 53338 37752 53340
rect 37776 53338 37832 53340
rect 37856 53338 37912 53340
rect 37616 53286 37662 53338
rect 37662 53286 37672 53338
rect 37696 53286 37726 53338
rect 37726 53286 37738 53338
rect 37738 53286 37752 53338
rect 37776 53286 37790 53338
rect 37790 53286 37802 53338
rect 37802 53286 37832 53338
rect 37856 53286 37866 53338
rect 37866 53286 37912 53338
rect 37616 53284 37672 53286
rect 37696 53284 37752 53286
rect 37776 53284 37832 53286
rect 37856 53284 37912 53286
rect 37616 52250 37672 52252
rect 37696 52250 37752 52252
rect 37776 52250 37832 52252
rect 37856 52250 37912 52252
rect 37616 52198 37662 52250
rect 37662 52198 37672 52250
rect 37696 52198 37726 52250
rect 37726 52198 37738 52250
rect 37738 52198 37752 52250
rect 37776 52198 37790 52250
rect 37790 52198 37802 52250
rect 37802 52198 37832 52250
rect 37856 52198 37866 52250
rect 37866 52198 37912 52250
rect 37616 52196 37672 52198
rect 37696 52196 37752 52198
rect 37776 52196 37832 52198
rect 37856 52196 37912 52198
rect 37616 51162 37672 51164
rect 37696 51162 37752 51164
rect 37776 51162 37832 51164
rect 37856 51162 37912 51164
rect 37616 51110 37662 51162
rect 37662 51110 37672 51162
rect 37696 51110 37726 51162
rect 37726 51110 37738 51162
rect 37738 51110 37752 51162
rect 37776 51110 37790 51162
rect 37790 51110 37802 51162
rect 37802 51110 37832 51162
rect 37856 51110 37866 51162
rect 37866 51110 37912 51162
rect 37616 51108 37672 51110
rect 37696 51108 37752 51110
rect 37776 51108 37832 51110
rect 37856 51108 37912 51110
rect 37616 50074 37672 50076
rect 37696 50074 37752 50076
rect 37776 50074 37832 50076
rect 37856 50074 37912 50076
rect 37616 50022 37662 50074
rect 37662 50022 37672 50074
rect 37696 50022 37726 50074
rect 37726 50022 37738 50074
rect 37738 50022 37752 50074
rect 37776 50022 37790 50074
rect 37790 50022 37802 50074
rect 37802 50022 37832 50074
rect 37856 50022 37866 50074
rect 37866 50022 37912 50074
rect 37616 50020 37672 50022
rect 37696 50020 37752 50022
rect 37776 50020 37832 50022
rect 37856 50020 37912 50022
rect 37616 48986 37672 48988
rect 37696 48986 37752 48988
rect 37776 48986 37832 48988
rect 37856 48986 37912 48988
rect 37616 48934 37662 48986
rect 37662 48934 37672 48986
rect 37696 48934 37726 48986
rect 37726 48934 37738 48986
rect 37738 48934 37752 48986
rect 37776 48934 37790 48986
rect 37790 48934 37802 48986
rect 37802 48934 37832 48986
rect 37856 48934 37866 48986
rect 37866 48934 37912 48986
rect 37616 48932 37672 48934
rect 37696 48932 37752 48934
rect 37776 48932 37832 48934
rect 37856 48932 37912 48934
rect 37616 47898 37672 47900
rect 37696 47898 37752 47900
rect 37776 47898 37832 47900
rect 37856 47898 37912 47900
rect 37616 47846 37662 47898
rect 37662 47846 37672 47898
rect 37696 47846 37726 47898
rect 37726 47846 37738 47898
rect 37738 47846 37752 47898
rect 37776 47846 37790 47898
rect 37790 47846 37802 47898
rect 37802 47846 37832 47898
rect 37856 47846 37866 47898
rect 37866 47846 37912 47898
rect 37616 47844 37672 47846
rect 37696 47844 37752 47846
rect 37776 47844 37832 47846
rect 37856 47844 37912 47846
rect 37616 46810 37672 46812
rect 37696 46810 37752 46812
rect 37776 46810 37832 46812
rect 37856 46810 37912 46812
rect 37616 46758 37662 46810
rect 37662 46758 37672 46810
rect 37696 46758 37726 46810
rect 37726 46758 37738 46810
rect 37738 46758 37752 46810
rect 37776 46758 37790 46810
rect 37790 46758 37802 46810
rect 37802 46758 37832 46810
rect 37856 46758 37866 46810
rect 37866 46758 37912 46810
rect 37616 46756 37672 46758
rect 37696 46756 37752 46758
rect 37776 46756 37832 46758
rect 37856 46756 37912 46758
rect 37616 45722 37672 45724
rect 37696 45722 37752 45724
rect 37776 45722 37832 45724
rect 37856 45722 37912 45724
rect 37616 45670 37662 45722
rect 37662 45670 37672 45722
rect 37696 45670 37726 45722
rect 37726 45670 37738 45722
rect 37738 45670 37752 45722
rect 37776 45670 37790 45722
rect 37790 45670 37802 45722
rect 37802 45670 37832 45722
rect 37856 45670 37866 45722
rect 37866 45670 37912 45722
rect 37616 45668 37672 45670
rect 37696 45668 37752 45670
rect 37776 45668 37832 45670
rect 37856 45668 37912 45670
rect 37616 44634 37672 44636
rect 37696 44634 37752 44636
rect 37776 44634 37832 44636
rect 37856 44634 37912 44636
rect 37616 44582 37662 44634
rect 37662 44582 37672 44634
rect 37696 44582 37726 44634
rect 37726 44582 37738 44634
rect 37738 44582 37752 44634
rect 37776 44582 37790 44634
rect 37790 44582 37802 44634
rect 37802 44582 37832 44634
rect 37856 44582 37866 44634
rect 37866 44582 37912 44634
rect 37616 44580 37672 44582
rect 37696 44580 37752 44582
rect 37776 44580 37832 44582
rect 37856 44580 37912 44582
rect 37616 43546 37672 43548
rect 37696 43546 37752 43548
rect 37776 43546 37832 43548
rect 37856 43546 37912 43548
rect 37616 43494 37662 43546
rect 37662 43494 37672 43546
rect 37696 43494 37726 43546
rect 37726 43494 37738 43546
rect 37738 43494 37752 43546
rect 37776 43494 37790 43546
rect 37790 43494 37802 43546
rect 37802 43494 37832 43546
rect 37856 43494 37866 43546
rect 37866 43494 37912 43546
rect 37616 43492 37672 43494
rect 37696 43492 37752 43494
rect 37776 43492 37832 43494
rect 37856 43492 37912 43494
rect 37616 42458 37672 42460
rect 37696 42458 37752 42460
rect 37776 42458 37832 42460
rect 37856 42458 37912 42460
rect 37616 42406 37662 42458
rect 37662 42406 37672 42458
rect 37696 42406 37726 42458
rect 37726 42406 37738 42458
rect 37738 42406 37752 42458
rect 37776 42406 37790 42458
rect 37790 42406 37802 42458
rect 37802 42406 37832 42458
rect 37856 42406 37866 42458
rect 37866 42406 37912 42458
rect 37616 42404 37672 42406
rect 37696 42404 37752 42406
rect 37776 42404 37832 42406
rect 37856 42404 37912 42406
rect 37616 41370 37672 41372
rect 37696 41370 37752 41372
rect 37776 41370 37832 41372
rect 37856 41370 37912 41372
rect 37616 41318 37662 41370
rect 37662 41318 37672 41370
rect 37696 41318 37726 41370
rect 37726 41318 37738 41370
rect 37738 41318 37752 41370
rect 37776 41318 37790 41370
rect 37790 41318 37802 41370
rect 37802 41318 37832 41370
rect 37856 41318 37866 41370
rect 37866 41318 37912 41370
rect 37616 41316 37672 41318
rect 37696 41316 37752 41318
rect 37776 41316 37832 41318
rect 37856 41316 37912 41318
rect 37616 40282 37672 40284
rect 37696 40282 37752 40284
rect 37776 40282 37832 40284
rect 37856 40282 37912 40284
rect 37616 40230 37662 40282
rect 37662 40230 37672 40282
rect 37696 40230 37726 40282
rect 37726 40230 37738 40282
rect 37738 40230 37752 40282
rect 37776 40230 37790 40282
rect 37790 40230 37802 40282
rect 37802 40230 37832 40282
rect 37856 40230 37866 40282
rect 37866 40230 37912 40282
rect 37616 40228 37672 40230
rect 37696 40228 37752 40230
rect 37776 40228 37832 40230
rect 37856 40228 37912 40230
rect 37616 39194 37672 39196
rect 37696 39194 37752 39196
rect 37776 39194 37832 39196
rect 37856 39194 37912 39196
rect 37616 39142 37662 39194
rect 37662 39142 37672 39194
rect 37696 39142 37726 39194
rect 37726 39142 37738 39194
rect 37738 39142 37752 39194
rect 37776 39142 37790 39194
rect 37790 39142 37802 39194
rect 37802 39142 37832 39194
rect 37856 39142 37866 39194
rect 37866 39142 37912 39194
rect 37616 39140 37672 39142
rect 37696 39140 37752 39142
rect 37776 39140 37832 39142
rect 37856 39140 37912 39142
rect 37616 38106 37672 38108
rect 37696 38106 37752 38108
rect 37776 38106 37832 38108
rect 37856 38106 37912 38108
rect 37616 38054 37662 38106
rect 37662 38054 37672 38106
rect 37696 38054 37726 38106
rect 37726 38054 37738 38106
rect 37738 38054 37752 38106
rect 37776 38054 37790 38106
rect 37790 38054 37802 38106
rect 37802 38054 37832 38106
rect 37856 38054 37866 38106
rect 37866 38054 37912 38106
rect 37616 38052 37672 38054
rect 37696 38052 37752 38054
rect 37776 38052 37832 38054
rect 37856 38052 37912 38054
rect 37616 37018 37672 37020
rect 37696 37018 37752 37020
rect 37776 37018 37832 37020
rect 37856 37018 37912 37020
rect 37616 36966 37662 37018
rect 37662 36966 37672 37018
rect 37696 36966 37726 37018
rect 37726 36966 37738 37018
rect 37738 36966 37752 37018
rect 37776 36966 37790 37018
rect 37790 36966 37802 37018
rect 37802 36966 37832 37018
rect 37856 36966 37866 37018
rect 37866 36966 37912 37018
rect 37616 36964 37672 36966
rect 37696 36964 37752 36966
rect 37776 36964 37832 36966
rect 37856 36964 37912 36966
rect 37616 35930 37672 35932
rect 37696 35930 37752 35932
rect 37776 35930 37832 35932
rect 37856 35930 37912 35932
rect 37616 35878 37662 35930
rect 37662 35878 37672 35930
rect 37696 35878 37726 35930
rect 37726 35878 37738 35930
rect 37738 35878 37752 35930
rect 37776 35878 37790 35930
rect 37790 35878 37802 35930
rect 37802 35878 37832 35930
rect 37856 35878 37866 35930
rect 37866 35878 37912 35930
rect 37616 35876 37672 35878
rect 37696 35876 37752 35878
rect 37776 35876 37832 35878
rect 37856 35876 37912 35878
rect 37616 34842 37672 34844
rect 37696 34842 37752 34844
rect 37776 34842 37832 34844
rect 37856 34842 37912 34844
rect 37616 34790 37662 34842
rect 37662 34790 37672 34842
rect 37696 34790 37726 34842
rect 37726 34790 37738 34842
rect 37738 34790 37752 34842
rect 37776 34790 37790 34842
rect 37790 34790 37802 34842
rect 37802 34790 37832 34842
rect 37856 34790 37866 34842
rect 37866 34790 37912 34842
rect 37616 34788 37672 34790
rect 37696 34788 37752 34790
rect 37776 34788 37832 34790
rect 37856 34788 37912 34790
rect 37616 33754 37672 33756
rect 37696 33754 37752 33756
rect 37776 33754 37832 33756
rect 37856 33754 37912 33756
rect 37616 33702 37662 33754
rect 37662 33702 37672 33754
rect 37696 33702 37726 33754
rect 37726 33702 37738 33754
rect 37738 33702 37752 33754
rect 37776 33702 37790 33754
rect 37790 33702 37802 33754
rect 37802 33702 37832 33754
rect 37856 33702 37866 33754
rect 37866 33702 37912 33754
rect 37616 33700 37672 33702
rect 37696 33700 37752 33702
rect 37776 33700 37832 33702
rect 37856 33700 37912 33702
rect 37616 32666 37672 32668
rect 37696 32666 37752 32668
rect 37776 32666 37832 32668
rect 37856 32666 37912 32668
rect 37616 32614 37662 32666
rect 37662 32614 37672 32666
rect 37696 32614 37726 32666
rect 37726 32614 37738 32666
rect 37738 32614 37752 32666
rect 37776 32614 37790 32666
rect 37790 32614 37802 32666
rect 37802 32614 37832 32666
rect 37856 32614 37866 32666
rect 37866 32614 37912 32666
rect 37616 32612 37672 32614
rect 37696 32612 37752 32614
rect 37776 32612 37832 32614
rect 37856 32612 37912 32614
rect 37616 31578 37672 31580
rect 37696 31578 37752 31580
rect 37776 31578 37832 31580
rect 37856 31578 37912 31580
rect 37616 31526 37662 31578
rect 37662 31526 37672 31578
rect 37696 31526 37726 31578
rect 37726 31526 37738 31578
rect 37738 31526 37752 31578
rect 37776 31526 37790 31578
rect 37790 31526 37802 31578
rect 37802 31526 37832 31578
rect 37856 31526 37866 31578
rect 37866 31526 37912 31578
rect 37616 31524 37672 31526
rect 37696 31524 37752 31526
rect 37776 31524 37832 31526
rect 37856 31524 37912 31526
rect 37616 30490 37672 30492
rect 37696 30490 37752 30492
rect 37776 30490 37832 30492
rect 37856 30490 37912 30492
rect 37616 30438 37662 30490
rect 37662 30438 37672 30490
rect 37696 30438 37726 30490
rect 37726 30438 37738 30490
rect 37738 30438 37752 30490
rect 37776 30438 37790 30490
rect 37790 30438 37802 30490
rect 37802 30438 37832 30490
rect 37856 30438 37866 30490
rect 37866 30438 37912 30490
rect 37616 30436 37672 30438
rect 37696 30436 37752 30438
rect 37776 30436 37832 30438
rect 37856 30436 37912 30438
rect 37616 29402 37672 29404
rect 37696 29402 37752 29404
rect 37776 29402 37832 29404
rect 37856 29402 37912 29404
rect 37616 29350 37662 29402
rect 37662 29350 37672 29402
rect 37696 29350 37726 29402
rect 37726 29350 37738 29402
rect 37738 29350 37752 29402
rect 37776 29350 37790 29402
rect 37790 29350 37802 29402
rect 37802 29350 37832 29402
rect 37856 29350 37866 29402
rect 37866 29350 37912 29402
rect 37616 29348 37672 29350
rect 37696 29348 37752 29350
rect 37776 29348 37832 29350
rect 37856 29348 37912 29350
rect 37616 28314 37672 28316
rect 37696 28314 37752 28316
rect 37776 28314 37832 28316
rect 37856 28314 37912 28316
rect 37616 28262 37662 28314
rect 37662 28262 37672 28314
rect 37696 28262 37726 28314
rect 37726 28262 37738 28314
rect 37738 28262 37752 28314
rect 37776 28262 37790 28314
rect 37790 28262 37802 28314
rect 37802 28262 37832 28314
rect 37856 28262 37866 28314
rect 37866 28262 37912 28314
rect 37616 28260 37672 28262
rect 37696 28260 37752 28262
rect 37776 28260 37832 28262
rect 37856 28260 37912 28262
rect 37616 27226 37672 27228
rect 37696 27226 37752 27228
rect 37776 27226 37832 27228
rect 37856 27226 37912 27228
rect 37616 27174 37662 27226
rect 37662 27174 37672 27226
rect 37696 27174 37726 27226
rect 37726 27174 37738 27226
rect 37738 27174 37752 27226
rect 37776 27174 37790 27226
rect 37790 27174 37802 27226
rect 37802 27174 37832 27226
rect 37856 27174 37866 27226
rect 37866 27174 37912 27226
rect 37616 27172 37672 27174
rect 37696 27172 37752 27174
rect 37776 27172 37832 27174
rect 37856 27172 37912 27174
rect 37616 26138 37672 26140
rect 37696 26138 37752 26140
rect 37776 26138 37832 26140
rect 37856 26138 37912 26140
rect 37616 26086 37662 26138
rect 37662 26086 37672 26138
rect 37696 26086 37726 26138
rect 37726 26086 37738 26138
rect 37738 26086 37752 26138
rect 37776 26086 37790 26138
rect 37790 26086 37802 26138
rect 37802 26086 37832 26138
rect 37856 26086 37866 26138
rect 37866 26086 37912 26138
rect 37616 26084 37672 26086
rect 37696 26084 37752 26086
rect 37776 26084 37832 26086
rect 37856 26084 37912 26086
rect 37616 25050 37672 25052
rect 37696 25050 37752 25052
rect 37776 25050 37832 25052
rect 37856 25050 37912 25052
rect 37616 24998 37662 25050
rect 37662 24998 37672 25050
rect 37696 24998 37726 25050
rect 37726 24998 37738 25050
rect 37738 24998 37752 25050
rect 37776 24998 37790 25050
rect 37790 24998 37802 25050
rect 37802 24998 37832 25050
rect 37856 24998 37866 25050
rect 37866 24998 37912 25050
rect 37616 24996 37672 24998
rect 37696 24996 37752 24998
rect 37776 24996 37832 24998
rect 37856 24996 37912 24998
rect 37616 23962 37672 23964
rect 37696 23962 37752 23964
rect 37776 23962 37832 23964
rect 37856 23962 37912 23964
rect 37616 23910 37662 23962
rect 37662 23910 37672 23962
rect 37696 23910 37726 23962
rect 37726 23910 37738 23962
rect 37738 23910 37752 23962
rect 37776 23910 37790 23962
rect 37790 23910 37802 23962
rect 37802 23910 37832 23962
rect 37856 23910 37866 23962
rect 37866 23910 37912 23962
rect 37616 23908 37672 23910
rect 37696 23908 37752 23910
rect 37776 23908 37832 23910
rect 37856 23908 37912 23910
rect 37616 22874 37672 22876
rect 37696 22874 37752 22876
rect 37776 22874 37832 22876
rect 37856 22874 37912 22876
rect 37616 22822 37662 22874
rect 37662 22822 37672 22874
rect 37696 22822 37726 22874
rect 37726 22822 37738 22874
rect 37738 22822 37752 22874
rect 37776 22822 37790 22874
rect 37790 22822 37802 22874
rect 37802 22822 37832 22874
rect 37856 22822 37866 22874
rect 37866 22822 37912 22874
rect 37616 22820 37672 22822
rect 37696 22820 37752 22822
rect 37776 22820 37832 22822
rect 37856 22820 37912 22822
rect 37616 21786 37672 21788
rect 37696 21786 37752 21788
rect 37776 21786 37832 21788
rect 37856 21786 37912 21788
rect 37616 21734 37662 21786
rect 37662 21734 37672 21786
rect 37696 21734 37726 21786
rect 37726 21734 37738 21786
rect 37738 21734 37752 21786
rect 37776 21734 37790 21786
rect 37790 21734 37802 21786
rect 37802 21734 37832 21786
rect 37856 21734 37866 21786
rect 37866 21734 37912 21786
rect 37616 21732 37672 21734
rect 37696 21732 37752 21734
rect 37776 21732 37832 21734
rect 37856 21732 37912 21734
rect 36956 21242 37012 21244
rect 37036 21242 37092 21244
rect 37116 21242 37172 21244
rect 37196 21242 37252 21244
rect 36956 21190 37002 21242
rect 37002 21190 37012 21242
rect 37036 21190 37066 21242
rect 37066 21190 37078 21242
rect 37078 21190 37092 21242
rect 37116 21190 37130 21242
rect 37130 21190 37142 21242
rect 37142 21190 37172 21242
rect 37196 21190 37206 21242
rect 37206 21190 37252 21242
rect 36956 21188 37012 21190
rect 37036 21188 37092 21190
rect 37116 21188 37172 21190
rect 37196 21188 37252 21190
rect 37616 20698 37672 20700
rect 37696 20698 37752 20700
rect 37776 20698 37832 20700
rect 37856 20698 37912 20700
rect 37616 20646 37662 20698
rect 37662 20646 37672 20698
rect 37696 20646 37726 20698
rect 37726 20646 37738 20698
rect 37738 20646 37752 20698
rect 37776 20646 37790 20698
rect 37790 20646 37802 20698
rect 37802 20646 37832 20698
rect 37856 20646 37866 20698
rect 37866 20646 37912 20698
rect 37616 20644 37672 20646
rect 37696 20644 37752 20646
rect 37776 20644 37832 20646
rect 37856 20644 37912 20646
rect 36956 20154 37012 20156
rect 37036 20154 37092 20156
rect 37116 20154 37172 20156
rect 37196 20154 37252 20156
rect 36956 20102 37002 20154
rect 37002 20102 37012 20154
rect 37036 20102 37066 20154
rect 37066 20102 37078 20154
rect 37078 20102 37092 20154
rect 37116 20102 37130 20154
rect 37130 20102 37142 20154
rect 37142 20102 37172 20154
rect 37196 20102 37206 20154
rect 37206 20102 37252 20154
rect 36956 20100 37012 20102
rect 37036 20100 37092 20102
rect 37116 20100 37172 20102
rect 37196 20100 37252 20102
rect 37616 19610 37672 19612
rect 37696 19610 37752 19612
rect 37776 19610 37832 19612
rect 37856 19610 37912 19612
rect 37616 19558 37662 19610
rect 37662 19558 37672 19610
rect 37696 19558 37726 19610
rect 37726 19558 37738 19610
rect 37738 19558 37752 19610
rect 37776 19558 37790 19610
rect 37790 19558 37802 19610
rect 37802 19558 37832 19610
rect 37856 19558 37866 19610
rect 37866 19558 37912 19610
rect 37616 19556 37672 19558
rect 37696 19556 37752 19558
rect 37776 19556 37832 19558
rect 37856 19556 37912 19558
rect 36956 19066 37012 19068
rect 37036 19066 37092 19068
rect 37116 19066 37172 19068
rect 37196 19066 37252 19068
rect 36956 19014 37002 19066
rect 37002 19014 37012 19066
rect 37036 19014 37066 19066
rect 37066 19014 37078 19066
rect 37078 19014 37092 19066
rect 37116 19014 37130 19066
rect 37130 19014 37142 19066
rect 37142 19014 37172 19066
rect 37196 19014 37206 19066
rect 37206 19014 37252 19066
rect 36956 19012 37012 19014
rect 37036 19012 37092 19014
rect 37116 19012 37172 19014
rect 37196 19012 37252 19014
rect 37616 18522 37672 18524
rect 37696 18522 37752 18524
rect 37776 18522 37832 18524
rect 37856 18522 37912 18524
rect 37616 18470 37662 18522
rect 37662 18470 37672 18522
rect 37696 18470 37726 18522
rect 37726 18470 37738 18522
rect 37738 18470 37752 18522
rect 37776 18470 37790 18522
rect 37790 18470 37802 18522
rect 37802 18470 37832 18522
rect 37856 18470 37866 18522
rect 37866 18470 37912 18522
rect 37616 18468 37672 18470
rect 37696 18468 37752 18470
rect 37776 18468 37832 18470
rect 37856 18468 37912 18470
rect 32616 8730 32672 8732
rect 32696 8730 32752 8732
rect 32776 8730 32832 8732
rect 32856 8730 32912 8732
rect 32616 8678 32662 8730
rect 32662 8678 32672 8730
rect 32696 8678 32726 8730
rect 32726 8678 32738 8730
rect 32738 8678 32752 8730
rect 32776 8678 32790 8730
rect 32790 8678 32802 8730
rect 32802 8678 32832 8730
rect 32856 8678 32866 8730
rect 32866 8678 32912 8730
rect 32616 8676 32672 8678
rect 32696 8676 32752 8678
rect 32776 8676 32832 8678
rect 32856 8676 32912 8678
rect 31956 8186 32012 8188
rect 32036 8186 32092 8188
rect 32116 8186 32172 8188
rect 32196 8186 32252 8188
rect 31956 8134 32002 8186
rect 32002 8134 32012 8186
rect 32036 8134 32066 8186
rect 32066 8134 32078 8186
rect 32078 8134 32092 8186
rect 32116 8134 32130 8186
rect 32130 8134 32142 8186
rect 32142 8134 32172 8186
rect 32196 8134 32206 8186
rect 32206 8134 32252 8186
rect 31956 8132 32012 8134
rect 32036 8132 32092 8134
rect 32116 8132 32172 8134
rect 32196 8132 32252 8134
rect 32616 7642 32672 7644
rect 32696 7642 32752 7644
rect 32776 7642 32832 7644
rect 32856 7642 32912 7644
rect 32616 7590 32662 7642
rect 32662 7590 32672 7642
rect 32696 7590 32726 7642
rect 32726 7590 32738 7642
rect 32738 7590 32752 7642
rect 32776 7590 32790 7642
rect 32790 7590 32802 7642
rect 32802 7590 32832 7642
rect 32856 7590 32866 7642
rect 32866 7590 32912 7642
rect 32616 7588 32672 7590
rect 32696 7588 32752 7590
rect 32776 7588 32832 7590
rect 32856 7588 32912 7590
rect 31956 7098 32012 7100
rect 32036 7098 32092 7100
rect 32116 7098 32172 7100
rect 32196 7098 32252 7100
rect 31956 7046 32002 7098
rect 32002 7046 32012 7098
rect 32036 7046 32066 7098
rect 32066 7046 32078 7098
rect 32078 7046 32092 7098
rect 32116 7046 32130 7098
rect 32130 7046 32142 7098
rect 32142 7046 32172 7098
rect 32196 7046 32206 7098
rect 32206 7046 32252 7098
rect 31956 7044 32012 7046
rect 32036 7044 32092 7046
rect 32116 7044 32172 7046
rect 32196 7044 32252 7046
rect 32616 6554 32672 6556
rect 32696 6554 32752 6556
rect 32776 6554 32832 6556
rect 32856 6554 32912 6556
rect 32616 6502 32662 6554
rect 32662 6502 32672 6554
rect 32696 6502 32726 6554
rect 32726 6502 32738 6554
rect 32738 6502 32752 6554
rect 32776 6502 32790 6554
rect 32790 6502 32802 6554
rect 32802 6502 32832 6554
rect 32856 6502 32866 6554
rect 32866 6502 32912 6554
rect 32616 6500 32672 6502
rect 32696 6500 32752 6502
rect 32776 6500 32832 6502
rect 32856 6500 32912 6502
rect 31956 6010 32012 6012
rect 32036 6010 32092 6012
rect 32116 6010 32172 6012
rect 32196 6010 32252 6012
rect 31956 5958 32002 6010
rect 32002 5958 32012 6010
rect 32036 5958 32066 6010
rect 32066 5958 32078 6010
rect 32078 5958 32092 6010
rect 32116 5958 32130 6010
rect 32130 5958 32142 6010
rect 32142 5958 32172 6010
rect 32196 5958 32206 6010
rect 32206 5958 32252 6010
rect 31956 5956 32012 5958
rect 32036 5956 32092 5958
rect 32116 5956 32172 5958
rect 32196 5956 32252 5958
rect 32616 5466 32672 5468
rect 32696 5466 32752 5468
rect 32776 5466 32832 5468
rect 32856 5466 32912 5468
rect 32616 5414 32662 5466
rect 32662 5414 32672 5466
rect 32696 5414 32726 5466
rect 32726 5414 32738 5466
rect 32738 5414 32752 5466
rect 32776 5414 32790 5466
rect 32790 5414 32802 5466
rect 32802 5414 32832 5466
rect 32856 5414 32866 5466
rect 32866 5414 32912 5466
rect 32616 5412 32672 5414
rect 32696 5412 32752 5414
rect 32776 5412 32832 5414
rect 32856 5412 32912 5414
rect 31956 4922 32012 4924
rect 32036 4922 32092 4924
rect 32116 4922 32172 4924
rect 32196 4922 32252 4924
rect 31956 4870 32002 4922
rect 32002 4870 32012 4922
rect 32036 4870 32066 4922
rect 32066 4870 32078 4922
rect 32078 4870 32092 4922
rect 32116 4870 32130 4922
rect 32130 4870 32142 4922
rect 32142 4870 32172 4922
rect 32196 4870 32206 4922
rect 32206 4870 32252 4922
rect 31956 4868 32012 4870
rect 32036 4868 32092 4870
rect 32116 4868 32172 4870
rect 32196 4868 32252 4870
rect 32616 4378 32672 4380
rect 32696 4378 32752 4380
rect 32776 4378 32832 4380
rect 32856 4378 32912 4380
rect 32616 4326 32662 4378
rect 32662 4326 32672 4378
rect 32696 4326 32726 4378
rect 32726 4326 32738 4378
rect 32738 4326 32752 4378
rect 32776 4326 32790 4378
rect 32790 4326 32802 4378
rect 32802 4326 32832 4378
rect 32856 4326 32866 4378
rect 32866 4326 32912 4378
rect 32616 4324 32672 4326
rect 32696 4324 32752 4326
rect 32776 4324 32832 4326
rect 32856 4324 32912 4326
rect 31956 3834 32012 3836
rect 32036 3834 32092 3836
rect 32116 3834 32172 3836
rect 32196 3834 32252 3836
rect 31956 3782 32002 3834
rect 32002 3782 32012 3834
rect 32036 3782 32066 3834
rect 32066 3782 32078 3834
rect 32078 3782 32092 3834
rect 32116 3782 32130 3834
rect 32130 3782 32142 3834
rect 32142 3782 32172 3834
rect 32196 3782 32206 3834
rect 32206 3782 32252 3834
rect 31956 3780 32012 3782
rect 32036 3780 32092 3782
rect 32116 3780 32172 3782
rect 32196 3780 32252 3782
rect 32616 3290 32672 3292
rect 32696 3290 32752 3292
rect 32776 3290 32832 3292
rect 32856 3290 32912 3292
rect 32616 3238 32662 3290
rect 32662 3238 32672 3290
rect 32696 3238 32726 3290
rect 32726 3238 32738 3290
rect 32738 3238 32752 3290
rect 32776 3238 32790 3290
rect 32790 3238 32802 3290
rect 32802 3238 32832 3290
rect 32856 3238 32866 3290
rect 32866 3238 32912 3290
rect 32616 3236 32672 3238
rect 32696 3236 32752 3238
rect 32776 3236 32832 3238
rect 32856 3236 32912 3238
rect 21956 2746 22012 2748
rect 22036 2746 22092 2748
rect 22116 2746 22172 2748
rect 22196 2746 22252 2748
rect 21956 2694 22002 2746
rect 22002 2694 22012 2746
rect 22036 2694 22066 2746
rect 22066 2694 22078 2746
rect 22078 2694 22092 2746
rect 22116 2694 22130 2746
rect 22130 2694 22142 2746
rect 22142 2694 22172 2746
rect 22196 2694 22206 2746
rect 22206 2694 22252 2746
rect 21956 2692 22012 2694
rect 22036 2692 22092 2694
rect 22116 2692 22172 2694
rect 22196 2692 22252 2694
rect 26956 2746 27012 2748
rect 27036 2746 27092 2748
rect 27116 2746 27172 2748
rect 27196 2746 27252 2748
rect 26956 2694 27002 2746
rect 27002 2694 27012 2746
rect 27036 2694 27066 2746
rect 27066 2694 27078 2746
rect 27078 2694 27092 2746
rect 27116 2694 27130 2746
rect 27130 2694 27142 2746
rect 27142 2694 27172 2746
rect 27196 2694 27206 2746
rect 27206 2694 27252 2746
rect 26956 2692 27012 2694
rect 27036 2692 27092 2694
rect 27116 2692 27172 2694
rect 27196 2692 27252 2694
rect 31956 2746 32012 2748
rect 32036 2746 32092 2748
rect 32116 2746 32172 2748
rect 32196 2746 32252 2748
rect 31956 2694 32002 2746
rect 32002 2694 32012 2746
rect 32036 2694 32066 2746
rect 32066 2694 32078 2746
rect 32078 2694 32092 2746
rect 32116 2694 32130 2746
rect 32130 2694 32142 2746
rect 32142 2694 32172 2746
rect 32196 2694 32206 2746
rect 32206 2694 32252 2746
rect 31956 2692 32012 2694
rect 32036 2692 32092 2694
rect 32116 2692 32172 2694
rect 32196 2692 32252 2694
rect 36956 17978 37012 17980
rect 37036 17978 37092 17980
rect 37116 17978 37172 17980
rect 37196 17978 37252 17980
rect 36956 17926 37002 17978
rect 37002 17926 37012 17978
rect 37036 17926 37066 17978
rect 37066 17926 37078 17978
rect 37078 17926 37092 17978
rect 37116 17926 37130 17978
rect 37130 17926 37142 17978
rect 37142 17926 37172 17978
rect 37196 17926 37206 17978
rect 37206 17926 37252 17978
rect 36956 17924 37012 17926
rect 37036 17924 37092 17926
rect 37116 17924 37172 17926
rect 37196 17924 37252 17926
rect 37616 17434 37672 17436
rect 37696 17434 37752 17436
rect 37776 17434 37832 17436
rect 37856 17434 37912 17436
rect 37616 17382 37662 17434
rect 37662 17382 37672 17434
rect 37696 17382 37726 17434
rect 37726 17382 37738 17434
rect 37738 17382 37752 17434
rect 37776 17382 37790 17434
rect 37790 17382 37802 17434
rect 37802 17382 37832 17434
rect 37856 17382 37866 17434
rect 37866 17382 37912 17434
rect 37616 17380 37672 17382
rect 37696 17380 37752 17382
rect 37776 17380 37832 17382
rect 37856 17380 37912 17382
rect 36956 16890 37012 16892
rect 37036 16890 37092 16892
rect 37116 16890 37172 16892
rect 37196 16890 37252 16892
rect 36956 16838 37002 16890
rect 37002 16838 37012 16890
rect 37036 16838 37066 16890
rect 37066 16838 37078 16890
rect 37078 16838 37092 16890
rect 37116 16838 37130 16890
rect 37130 16838 37142 16890
rect 37142 16838 37172 16890
rect 37196 16838 37206 16890
rect 37206 16838 37252 16890
rect 36956 16836 37012 16838
rect 37036 16836 37092 16838
rect 37116 16836 37172 16838
rect 37196 16836 37252 16838
rect 37616 16346 37672 16348
rect 37696 16346 37752 16348
rect 37776 16346 37832 16348
rect 37856 16346 37912 16348
rect 37616 16294 37662 16346
rect 37662 16294 37672 16346
rect 37696 16294 37726 16346
rect 37726 16294 37738 16346
rect 37738 16294 37752 16346
rect 37776 16294 37790 16346
rect 37790 16294 37802 16346
rect 37802 16294 37832 16346
rect 37856 16294 37866 16346
rect 37866 16294 37912 16346
rect 37616 16292 37672 16294
rect 37696 16292 37752 16294
rect 37776 16292 37832 16294
rect 37856 16292 37912 16294
rect 36956 15802 37012 15804
rect 37036 15802 37092 15804
rect 37116 15802 37172 15804
rect 37196 15802 37252 15804
rect 36956 15750 37002 15802
rect 37002 15750 37012 15802
rect 37036 15750 37066 15802
rect 37066 15750 37078 15802
rect 37078 15750 37092 15802
rect 37116 15750 37130 15802
rect 37130 15750 37142 15802
rect 37142 15750 37172 15802
rect 37196 15750 37206 15802
rect 37206 15750 37252 15802
rect 36956 15748 37012 15750
rect 37036 15748 37092 15750
rect 37116 15748 37172 15750
rect 37196 15748 37252 15750
rect 37616 15258 37672 15260
rect 37696 15258 37752 15260
rect 37776 15258 37832 15260
rect 37856 15258 37912 15260
rect 37616 15206 37662 15258
rect 37662 15206 37672 15258
rect 37696 15206 37726 15258
rect 37726 15206 37738 15258
rect 37738 15206 37752 15258
rect 37776 15206 37790 15258
rect 37790 15206 37802 15258
rect 37802 15206 37832 15258
rect 37856 15206 37866 15258
rect 37866 15206 37912 15258
rect 37616 15204 37672 15206
rect 37696 15204 37752 15206
rect 37776 15204 37832 15206
rect 37856 15204 37912 15206
rect 36956 14714 37012 14716
rect 37036 14714 37092 14716
rect 37116 14714 37172 14716
rect 37196 14714 37252 14716
rect 36956 14662 37002 14714
rect 37002 14662 37012 14714
rect 37036 14662 37066 14714
rect 37066 14662 37078 14714
rect 37078 14662 37092 14714
rect 37116 14662 37130 14714
rect 37130 14662 37142 14714
rect 37142 14662 37172 14714
rect 37196 14662 37206 14714
rect 37206 14662 37252 14714
rect 36956 14660 37012 14662
rect 37036 14660 37092 14662
rect 37116 14660 37172 14662
rect 37196 14660 37252 14662
rect 37616 14170 37672 14172
rect 37696 14170 37752 14172
rect 37776 14170 37832 14172
rect 37856 14170 37912 14172
rect 37616 14118 37662 14170
rect 37662 14118 37672 14170
rect 37696 14118 37726 14170
rect 37726 14118 37738 14170
rect 37738 14118 37752 14170
rect 37776 14118 37790 14170
rect 37790 14118 37802 14170
rect 37802 14118 37832 14170
rect 37856 14118 37866 14170
rect 37866 14118 37912 14170
rect 37616 14116 37672 14118
rect 37696 14116 37752 14118
rect 37776 14116 37832 14118
rect 37856 14116 37912 14118
rect 36956 13626 37012 13628
rect 37036 13626 37092 13628
rect 37116 13626 37172 13628
rect 37196 13626 37252 13628
rect 36956 13574 37002 13626
rect 37002 13574 37012 13626
rect 37036 13574 37066 13626
rect 37066 13574 37078 13626
rect 37078 13574 37092 13626
rect 37116 13574 37130 13626
rect 37130 13574 37142 13626
rect 37142 13574 37172 13626
rect 37196 13574 37206 13626
rect 37206 13574 37252 13626
rect 36956 13572 37012 13574
rect 37036 13572 37092 13574
rect 37116 13572 37172 13574
rect 37196 13572 37252 13574
rect 37616 13082 37672 13084
rect 37696 13082 37752 13084
rect 37776 13082 37832 13084
rect 37856 13082 37912 13084
rect 37616 13030 37662 13082
rect 37662 13030 37672 13082
rect 37696 13030 37726 13082
rect 37726 13030 37738 13082
rect 37738 13030 37752 13082
rect 37776 13030 37790 13082
rect 37790 13030 37802 13082
rect 37802 13030 37832 13082
rect 37856 13030 37866 13082
rect 37866 13030 37912 13082
rect 37616 13028 37672 13030
rect 37696 13028 37752 13030
rect 37776 13028 37832 13030
rect 37856 13028 37912 13030
rect 36956 12538 37012 12540
rect 37036 12538 37092 12540
rect 37116 12538 37172 12540
rect 37196 12538 37252 12540
rect 36956 12486 37002 12538
rect 37002 12486 37012 12538
rect 37036 12486 37066 12538
rect 37066 12486 37078 12538
rect 37078 12486 37092 12538
rect 37116 12486 37130 12538
rect 37130 12486 37142 12538
rect 37142 12486 37172 12538
rect 37196 12486 37206 12538
rect 37206 12486 37252 12538
rect 36956 12484 37012 12486
rect 37036 12484 37092 12486
rect 37116 12484 37172 12486
rect 37196 12484 37252 12486
rect 37616 11994 37672 11996
rect 37696 11994 37752 11996
rect 37776 11994 37832 11996
rect 37856 11994 37912 11996
rect 37616 11942 37662 11994
rect 37662 11942 37672 11994
rect 37696 11942 37726 11994
rect 37726 11942 37738 11994
rect 37738 11942 37752 11994
rect 37776 11942 37790 11994
rect 37790 11942 37802 11994
rect 37802 11942 37832 11994
rect 37856 11942 37866 11994
rect 37866 11942 37912 11994
rect 37616 11940 37672 11942
rect 37696 11940 37752 11942
rect 37776 11940 37832 11942
rect 37856 11940 37912 11942
rect 36956 11450 37012 11452
rect 37036 11450 37092 11452
rect 37116 11450 37172 11452
rect 37196 11450 37252 11452
rect 36956 11398 37002 11450
rect 37002 11398 37012 11450
rect 37036 11398 37066 11450
rect 37066 11398 37078 11450
rect 37078 11398 37092 11450
rect 37116 11398 37130 11450
rect 37130 11398 37142 11450
rect 37142 11398 37172 11450
rect 37196 11398 37206 11450
rect 37206 11398 37252 11450
rect 36956 11396 37012 11398
rect 37036 11396 37092 11398
rect 37116 11396 37172 11398
rect 37196 11396 37252 11398
rect 37616 10906 37672 10908
rect 37696 10906 37752 10908
rect 37776 10906 37832 10908
rect 37856 10906 37912 10908
rect 37616 10854 37662 10906
rect 37662 10854 37672 10906
rect 37696 10854 37726 10906
rect 37726 10854 37738 10906
rect 37738 10854 37752 10906
rect 37776 10854 37790 10906
rect 37790 10854 37802 10906
rect 37802 10854 37832 10906
rect 37856 10854 37866 10906
rect 37866 10854 37912 10906
rect 37616 10852 37672 10854
rect 37696 10852 37752 10854
rect 37776 10852 37832 10854
rect 37856 10852 37912 10854
rect 36956 10362 37012 10364
rect 37036 10362 37092 10364
rect 37116 10362 37172 10364
rect 37196 10362 37252 10364
rect 36956 10310 37002 10362
rect 37002 10310 37012 10362
rect 37036 10310 37066 10362
rect 37066 10310 37078 10362
rect 37078 10310 37092 10362
rect 37116 10310 37130 10362
rect 37130 10310 37142 10362
rect 37142 10310 37172 10362
rect 37196 10310 37206 10362
rect 37206 10310 37252 10362
rect 36956 10308 37012 10310
rect 37036 10308 37092 10310
rect 37116 10308 37172 10310
rect 37196 10308 37252 10310
rect 37616 9818 37672 9820
rect 37696 9818 37752 9820
rect 37776 9818 37832 9820
rect 37856 9818 37912 9820
rect 37616 9766 37662 9818
rect 37662 9766 37672 9818
rect 37696 9766 37726 9818
rect 37726 9766 37738 9818
rect 37738 9766 37752 9818
rect 37776 9766 37790 9818
rect 37790 9766 37802 9818
rect 37802 9766 37832 9818
rect 37856 9766 37866 9818
rect 37866 9766 37912 9818
rect 37616 9764 37672 9766
rect 37696 9764 37752 9766
rect 37776 9764 37832 9766
rect 37856 9764 37912 9766
rect 36956 9274 37012 9276
rect 37036 9274 37092 9276
rect 37116 9274 37172 9276
rect 37196 9274 37252 9276
rect 36956 9222 37002 9274
rect 37002 9222 37012 9274
rect 37036 9222 37066 9274
rect 37066 9222 37078 9274
rect 37078 9222 37092 9274
rect 37116 9222 37130 9274
rect 37130 9222 37142 9274
rect 37142 9222 37172 9274
rect 37196 9222 37206 9274
rect 37206 9222 37252 9274
rect 36956 9220 37012 9222
rect 37036 9220 37092 9222
rect 37116 9220 37172 9222
rect 37196 9220 37252 9222
rect 37616 8730 37672 8732
rect 37696 8730 37752 8732
rect 37776 8730 37832 8732
rect 37856 8730 37912 8732
rect 37616 8678 37662 8730
rect 37662 8678 37672 8730
rect 37696 8678 37726 8730
rect 37726 8678 37738 8730
rect 37738 8678 37752 8730
rect 37776 8678 37790 8730
rect 37790 8678 37802 8730
rect 37802 8678 37832 8730
rect 37856 8678 37866 8730
rect 37866 8678 37912 8730
rect 37616 8676 37672 8678
rect 37696 8676 37752 8678
rect 37776 8676 37832 8678
rect 37856 8676 37912 8678
rect 36956 8186 37012 8188
rect 37036 8186 37092 8188
rect 37116 8186 37172 8188
rect 37196 8186 37252 8188
rect 36956 8134 37002 8186
rect 37002 8134 37012 8186
rect 37036 8134 37066 8186
rect 37066 8134 37078 8186
rect 37078 8134 37092 8186
rect 37116 8134 37130 8186
rect 37130 8134 37142 8186
rect 37142 8134 37172 8186
rect 37196 8134 37206 8186
rect 37206 8134 37252 8186
rect 36956 8132 37012 8134
rect 37036 8132 37092 8134
rect 37116 8132 37172 8134
rect 37196 8132 37252 8134
rect 37616 7642 37672 7644
rect 37696 7642 37752 7644
rect 37776 7642 37832 7644
rect 37856 7642 37912 7644
rect 37616 7590 37662 7642
rect 37662 7590 37672 7642
rect 37696 7590 37726 7642
rect 37726 7590 37738 7642
rect 37738 7590 37752 7642
rect 37776 7590 37790 7642
rect 37790 7590 37802 7642
rect 37802 7590 37832 7642
rect 37856 7590 37866 7642
rect 37866 7590 37912 7642
rect 37616 7588 37672 7590
rect 37696 7588 37752 7590
rect 37776 7588 37832 7590
rect 37856 7588 37912 7590
rect 36956 7098 37012 7100
rect 37036 7098 37092 7100
rect 37116 7098 37172 7100
rect 37196 7098 37252 7100
rect 36956 7046 37002 7098
rect 37002 7046 37012 7098
rect 37036 7046 37066 7098
rect 37066 7046 37078 7098
rect 37078 7046 37092 7098
rect 37116 7046 37130 7098
rect 37130 7046 37142 7098
rect 37142 7046 37172 7098
rect 37196 7046 37206 7098
rect 37206 7046 37252 7098
rect 36956 7044 37012 7046
rect 37036 7044 37092 7046
rect 37116 7044 37172 7046
rect 37196 7044 37252 7046
rect 37616 6554 37672 6556
rect 37696 6554 37752 6556
rect 37776 6554 37832 6556
rect 37856 6554 37912 6556
rect 37616 6502 37662 6554
rect 37662 6502 37672 6554
rect 37696 6502 37726 6554
rect 37726 6502 37738 6554
rect 37738 6502 37752 6554
rect 37776 6502 37790 6554
rect 37790 6502 37802 6554
rect 37802 6502 37832 6554
rect 37856 6502 37866 6554
rect 37866 6502 37912 6554
rect 37616 6500 37672 6502
rect 37696 6500 37752 6502
rect 37776 6500 37832 6502
rect 37856 6500 37912 6502
rect 36956 6010 37012 6012
rect 37036 6010 37092 6012
rect 37116 6010 37172 6012
rect 37196 6010 37252 6012
rect 36956 5958 37002 6010
rect 37002 5958 37012 6010
rect 37036 5958 37066 6010
rect 37066 5958 37078 6010
rect 37078 5958 37092 6010
rect 37116 5958 37130 6010
rect 37130 5958 37142 6010
rect 37142 5958 37172 6010
rect 37196 5958 37206 6010
rect 37206 5958 37252 6010
rect 36956 5956 37012 5958
rect 37036 5956 37092 5958
rect 37116 5956 37172 5958
rect 37196 5956 37252 5958
rect 37616 5466 37672 5468
rect 37696 5466 37752 5468
rect 37776 5466 37832 5468
rect 37856 5466 37912 5468
rect 37616 5414 37662 5466
rect 37662 5414 37672 5466
rect 37696 5414 37726 5466
rect 37726 5414 37738 5466
rect 37738 5414 37752 5466
rect 37776 5414 37790 5466
rect 37790 5414 37802 5466
rect 37802 5414 37832 5466
rect 37856 5414 37866 5466
rect 37866 5414 37912 5466
rect 37616 5412 37672 5414
rect 37696 5412 37752 5414
rect 37776 5412 37832 5414
rect 37856 5412 37912 5414
rect 36956 4922 37012 4924
rect 37036 4922 37092 4924
rect 37116 4922 37172 4924
rect 37196 4922 37252 4924
rect 36956 4870 37002 4922
rect 37002 4870 37012 4922
rect 37036 4870 37066 4922
rect 37066 4870 37078 4922
rect 37078 4870 37092 4922
rect 37116 4870 37130 4922
rect 37130 4870 37142 4922
rect 37142 4870 37172 4922
rect 37196 4870 37206 4922
rect 37206 4870 37252 4922
rect 36956 4868 37012 4870
rect 37036 4868 37092 4870
rect 37116 4868 37172 4870
rect 37196 4868 37252 4870
rect 37616 4378 37672 4380
rect 37696 4378 37752 4380
rect 37776 4378 37832 4380
rect 37856 4378 37912 4380
rect 37616 4326 37662 4378
rect 37662 4326 37672 4378
rect 37696 4326 37726 4378
rect 37726 4326 37738 4378
rect 37738 4326 37752 4378
rect 37776 4326 37790 4378
rect 37790 4326 37802 4378
rect 37802 4326 37832 4378
rect 37856 4326 37866 4378
rect 37866 4326 37912 4378
rect 37616 4324 37672 4326
rect 37696 4324 37752 4326
rect 37776 4324 37832 4326
rect 37856 4324 37912 4326
rect 36956 3834 37012 3836
rect 37036 3834 37092 3836
rect 37116 3834 37172 3836
rect 37196 3834 37252 3836
rect 36956 3782 37002 3834
rect 37002 3782 37012 3834
rect 37036 3782 37066 3834
rect 37066 3782 37078 3834
rect 37078 3782 37092 3834
rect 37116 3782 37130 3834
rect 37130 3782 37142 3834
rect 37142 3782 37172 3834
rect 37196 3782 37206 3834
rect 37206 3782 37252 3834
rect 36956 3780 37012 3782
rect 37036 3780 37092 3782
rect 37116 3780 37172 3782
rect 37196 3780 37252 3782
rect 37616 3290 37672 3292
rect 37696 3290 37752 3292
rect 37776 3290 37832 3292
rect 37856 3290 37912 3292
rect 37616 3238 37662 3290
rect 37662 3238 37672 3290
rect 37696 3238 37726 3290
rect 37726 3238 37738 3290
rect 37738 3238 37752 3290
rect 37776 3238 37790 3290
rect 37790 3238 37802 3290
rect 37802 3238 37832 3290
rect 37856 3238 37866 3290
rect 37866 3238 37912 3290
rect 37616 3236 37672 3238
rect 37696 3236 37752 3238
rect 37776 3236 37832 3238
rect 37856 3236 37912 3238
rect 39118 30640 39174 30696
rect 38934 14356 38936 14376
rect 38936 14356 38988 14376
rect 38988 14356 38990 14376
rect 38934 14320 38990 14356
rect 40498 35944 40554 36000
rect 36956 2746 37012 2748
rect 37036 2746 37092 2748
rect 37116 2746 37172 2748
rect 37196 2746 37252 2748
rect 36956 2694 37002 2746
rect 37002 2694 37012 2746
rect 37036 2694 37066 2746
rect 37066 2694 37078 2746
rect 37078 2694 37092 2746
rect 37116 2694 37130 2746
rect 37130 2694 37142 2746
rect 37142 2694 37172 2746
rect 37196 2694 37206 2746
rect 37206 2694 37252 2746
rect 36956 2692 37012 2694
rect 37036 2692 37092 2694
rect 37116 2692 37172 2694
rect 37196 2692 37252 2694
rect 2616 2202 2672 2204
rect 2696 2202 2752 2204
rect 2776 2202 2832 2204
rect 2856 2202 2912 2204
rect 2616 2150 2662 2202
rect 2662 2150 2672 2202
rect 2696 2150 2726 2202
rect 2726 2150 2738 2202
rect 2738 2150 2752 2202
rect 2776 2150 2790 2202
rect 2790 2150 2802 2202
rect 2802 2150 2832 2202
rect 2856 2150 2866 2202
rect 2866 2150 2912 2202
rect 2616 2148 2672 2150
rect 2696 2148 2752 2150
rect 2776 2148 2832 2150
rect 2856 2148 2912 2150
rect 7616 2202 7672 2204
rect 7696 2202 7752 2204
rect 7776 2202 7832 2204
rect 7856 2202 7912 2204
rect 7616 2150 7662 2202
rect 7662 2150 7672 2202
rect 7696 2150 7726 2202
rect 7726 2150 7738 2202
rect 7738 2150 7752 2202
rect 7776 2150 7790 2202
rect 7790 2150 7802 2202
rect 7802 2150 7832 2202
rect 7856 2150 7866 2202
rect 7866 2150 7912 2202
rect 7616 2148 7672 2150
rect 7696 2148 7752 2150
rect 7776 2148 7832 2150
rect 7856 2148 7912 2150
rect 12616 2202 12672 2204
rect 12696 2202 12752 2204
rect 12776 2202 12832 2204
rect 12856 2202 12912 2204
rect 12616 2150 12662 2202
rect 12662 2150 12672 2202
rect 12696 2150 12726 2202
rect 12726 2150 12738 2202
rect 12738 2150 12752 2202
rect 12776 2150 12790 2202
rect 12790 2150 12802 2202
rect 12802 2150 12832 2202
rect 12856 2150 12866 2202
rect 12866 2150 12912 2202
rect 12616 2148 12672 2150
rect 12696 2148 12752 2150
rect 12776 2148 12832 2150
rect 12856 2148 12912 2150
rect 17616 2202 17672 2204
rect 17696 2202 17752 2204
rect 17776 2202 17832 2204
rect 17856 2202 17912 2204
rect 17616 2150 17662 2202
rect 17662 2150 17672 2202
rect 17696 2150 17726 2202
rect 17726 2150 17738 2202
rect 17738 2150 17752 2202
rect 17776 2150 17790 2202
rect 17790 2150 17802 2202
rect 17802 2150 17832 2202
rect 17856 2150 17866 2202
rect 17866 2150 17912 2202
rect 17616 2148 17672 2150
rect 17696 2148 17752 2150
rect 17776 2148 17832 2150
rect 17856 2148 17912 2150
rect 22616 2202 22672 2204
rect 22696 2202 22752 2204
rect 22776 2202 22832 2204
rect 22856 2202 22912 2204
rect 22616 2150 22662 2202
rect 22662 2150 22672 2202
rect 22696 2150 22726 2202
rect 22726 2150 22738 2202
rect 22738 2150 22752 2202
rect 22776 2150 22790 2202
rect 22790 2150 22802 2202
rect 22802 2150 22832 2202
rect 22856 2150 22866 2202
rect 22866 2150 22912 2202
rect 22616 2148 22672 2150
rect 22696 2148 22752 2150
rect 22776 2148 22832 2150
rect 22856 2148 22912 2150
rect 27616 2202 27672 2204
rect 27696 2202 27752 2204
rect 27776 2202 27832 2204
rect 27856 2202 27912 2204
rect 27616 2150 27662 2202
rect 27662 2150 27672 2202
rect 27696 2150 27726 2202
rect 27726 2150 27738 2202
rect 27738 2150 27752 2202
rect 27776 2150 27790 2202
rect 27790 2150 27802 2202
rect 27802 2150 27832 2202
rect 27856 2150 27866 2202
rect 27866 2150 27912 2202
rect 27616 2148 27672 2150
rect 27696 2148 27752 2150
rect 27776 2148 27832 2150
rect 27856 2148 27912 2150
rect 32616 2202 32672 2204
rect 32696 2202 32752 2204
rect 32776 2202 32832 2204
rect 32856 2202 32912 2204
rect 32616 2150 32662 2202
rect 32662 2150 32672 2202
rect 32696 2150 32726 2202
rect 32726 2150 32738 2202
rect 32738 2150 32752 2202
rect 32776 2150 32790 2202
rect 32790 2150 32802 2202
rect 32802 2150 32832 2202
rect 32856 2150 32866 2202
rect 32866 2150 32912 2202
rect 32616 2148 32672 2150
rect 32696 2148 32752 2150
rect 32776 2148 32832 2150
rect 32856 2148 32912 2150
rect 37616 2202 37672 2204
rect 37696 2202 37752 2204
rect 37776 2202 37832 2204
rect 37856 2202 37912 2204
rect 37616 2150 37662 2202
rect 37662 2150 37672 2202
rect 37696 2150 37726 2202
rect 37726 2150 37738 2202
rect 37738 2150 37752 2202
rect 37776 2150 37790 2202
rect 37790 2150 37802 2202
rect 37802 2150 37832 2202
rect 37856 2150 37866 2202
rect 37866 2150 37912 2202
rect 37616 2148 37672 2150
rect 37696 2148 37752 2150
rect 37776 2148 37832 2150
rect 37856 2148 37912 2150
<< metal3 >>
rect 2606 69664 2922 69665
rect 2606 69600 2612 69664
rect 2676 69600 2692 69664
rect 2756 69600 2772 69664
rect 2836 69600 2852 69664
rect 2916 69600 2922 69664
rect 2606 69599 2922 69600
rect 7606 69664 7922 69665
rect 7606 69600 7612 69664
rect 7676 69600 7692 69664
rect 7756 69600 7772 69664
rect 7836 69600 7852 69664
rect 7916 69600 7922 69664
rect 7606 69599 7922 69600
rect 12606 69664 12922 69665
rect 12606 69600 12612 69664
rect 12676 69600 12692 69664
rect 12756 69600 12772 69664
rect 12836 69600 12852 69664
rect 12916 69600 12922 69664
rect 12606 69599 12922 69600
rect 17606 69664 17922 69665
rect 17606 69600 17612 69664
rect 17676 69600 17692 69664
rect 17756 69600 17772 69664
rect 17836 69600 17852 69664
rect 17916 69600 17922 69664
rect 17606 69599 17922 69600
rect 22606 69664 22922 69665
rect 22606 69600 22612 69664
rect 22676 69600 22692 69664
rect 22756 69600 22772 69664
rect 22836 69600 22852 69664
rect 22916 69600 22922 69664
rect 22606 69599 22922 69600
rect 27606 69664 27922 69665
rect 27606 69600 27612 69664
rect 27676 69600 27692 69664
rect 27756 69600 27772 69664
rect 27836 69600 27852 69664
rect 27916 69600 27922 69664
rect 27606 69599 27922 69600
rect 32606 69664 32922 69665
rect 32606 69600 32612 69664
rect 32676 69600 32692 69664
rect 32756 69600 32772 69664
rect 32836 69600 32852 69664
rect 32916 69600 32922 69664
rect 32606 69599 32922 69600
rect 37606 69664 37922 69665
rect 37606 69600 37612 69664
rect 37676 69600 37692 69664
rect 37756 69600 37772 69664
rect 37836 69600 37852 69664
rect 37916 69600 37922 69664
rect 37606 69599 37922 69600
rect 1946 69120 2262 69121
rect 1946 69056 1952 69120
rect 2016 69056 2032 69120
rect 2096 69056 2112 69120
rect 2176 69056 2192 69120
rect 2256 69056 2262 69120
rect 1946 69055 2262 69056
rect 6946 69120 7262 69121
rect 6946 69056 6952 69120
rect 7016 69056 7032 69120
rect 7096 69056 7112 69120
rect 7176 69056 7192 69120
rect 7256 69056 7262 69120
rect 6946 69055 7262 69056
rect 11946 69120 12262 69121
rect 11946 69056 11952 69120
rect 12016 69056 12032 69120
rect 12096 69056 12112 69120
rect 12176 69056 12192 69120
rect 12256 69056 12262 69120
rect 11946 69055 12262 69056
rect 16946 69120 17262 69121
rect 16946 69056 16952 69120
rect 17016 69056 17032 69120
rect 17096 69056 17112 69120
rect 17176 69056 17192 69120
rect 17256 69056 17262 69120
rect 16946 69055 17262 69056
rect 21946 69120 22262 69121
rect 21946 69056 21952 69120
rect 22016 69056 22032 69120
rect 22096 69056 22112 69120
rect 22176 69056 22192 69120
rect 22256 69056 22262 69120
rect 21946 69055 22262 69056
rect 26946 69120 27262 69121
rect 26946 69056 26952 69120
rect 27016 69056 27032 69120
rect 27096 69056 27112 69120
rect 27176 69056 27192 69120
rect 27256 69056 27262 69120
rect 26946 69055 27262 69056
rect 31946 69120 32262 69121
rect 31946 69056 31952 69120
rect 32016 69056 32032 69120
rect 32096 69056 32112 69120
rect 32176 69056 32192 69120
rect 32256 69056 32262 69120
rect 31946 69055 32262 69056
rect 36946 69120 37262 69121
rect 36946 69056 36952 69120
rect 37016 69056 37032 69120
rect 37096 69056 37112 69120
rect 37176 69056 37192 69120
rect 37256 69056 37262 69120
rect 36946 69055 37262 69056
rect 2606 68576 2922 68577
rect 2606 68512 2612 68576
rect 2676 68512 2692 68576
rect 2756 68512 2772 68576
rect 2836 68512 2852 68576
rect 2916 68512 2922 68576
rect 2606 68511 2922 68512
rect 7606 68576 7922 68577
rect 7606 68512 7612 68576
rect 7676 68512 7692 68576
rect 7756 68512 7772 68576
rect 7836 68512 7852 68576
rect 7916 68512 7922 68576
rect 7606 68511 7922 68512
rect 12606 68576 12922 68577
rect 12606 68512 12612 68576
rect 12676 68512 12692 68576
rect 12756 68512 12772 68576
rect 12836 68512 12852 68576
rect 12916 68512 12922 68576
rect 12606 68511 12922 68512
rect 17606 68576 17922 68577
rect 17606 68512 17612 68576
rect 17676 68512 17692 68576
rect 17756 68512 17772 68576
rect 17836 68512 17852 68576
rect 17916 68512 17922 68576
rect 17606 68511 17922 68512
rect 22606 68576 22922 68577
rect 22606 68512 22612 68576
rect 22676 68512 22692 68576
rect 22756 68512 22772 68576
rect 22836 68512 22852 68576
rect 22916 68512 22922 68576
rect 22606 68511 22922 68512
rect 27606 68576 27922 68577
rect 27606 68512 27612 68576
rect 27676 68512 27692 68576
rect 27756 68512 27772 68576
rect 27836 68512 27852 68576
rect 27916 68512 27922 68576
rect 27606 68511 27922 68512
rect 32606 68576 32922 68577
rect 32606 68512 32612 68576
rect 32676 68512 32692 68576
rect 32756 68512 32772 68576
rect 32836 68512 32852 68576
rect 32916 68512 32922 68576
rect 32606 68511 32922 68512
rect 37606 68576 37922 68577
rect 37606 68512 37612 68576
rect 37676 68512 37692 68576
rect 37756 68512 37772 68576
rect 37836 68512 37852 68576
rect 37916 68512 37922 68576
rect 37606 68511 37922 68512
rect 1946 68032 2262 68033
rect 1946 67968 1952 68032
rect 2016 67968 2032 68032
rect 2096 67968 2112 68032
rect 2176 67968 2192 68032
rect 2256 67968 2262 68032
rect 1946 67967 2262 67968
rect 6946 68032 7262 68033
rect 6946 67968 6952 68032
rect 7016 67968 7032 68032
rect 7096 67968 7112 68032
rect 7176 67968 7192 68032
rect 7256 67968 7262 68032
rect 6946 67967 7262 67968
rect 11946 68032 12262 68033
rect 11946 67968 11952 68032
rect 12016 67968 12032 68032
rect 12096 67968 12112 68032
rect 12176 67968 12192 68032
rect 12256 67968 12262 68032
rect 11946 67967 12262 67968
rect 16946 68032 17262 68033
rect 16946 67968 16952 68032
rect 17016 67968 17032 68032
rect 17096 67968 17112 68032
rect 17176 67968 17192 68032
rect 17256 67968 17262 68032
rect 16946 67967 17262 67968
rect 21946 68032 22262 68033
rect 21946 67968 21952 68032
rect 22016 67968 22032 68032
rect 22096 67968 22112 68032
rect 22176 67968 22192 68032
rect 22256 67968 22262 68032
rect 21946 67967 22262 67968
rect 26946 68032 27262 68033
rect 26946 67968 26952 68032
rect 27016 67968 27032 68032
rect 27096 67968 27112 68032
rect 27176 67968 27192 68032
rect 27256 67968 27262 68032
rect 26946 67967 27262 67968
rect 31946 68032 32262 68033
rect 31946 67968 31952 68032
rect 32016 67968 32032 68032
rect 32096 67968 32112 68032
rect 32176 67968 32192 68032
rect 32256 67968 32262 68032
rect 31946 67967 32262 67968
rect 36946 68032 37262 68033
rect 36946 67968 36952 68032
rect 37016 67968 37032 68032
rect 37096 67968 37112 68032
rect 37176 67968 37192 68032
rect 37256 67968 37262 68032
rect 36946 67967 37262 67968
rect 31702 67628 31708 67692
rect 31772 67690 31778 67692
rect 32397 67690 32463 67693
rect 31772 67688 32463 67690
rect 31772 67632 32402 67688
rect 32458 67632 32463 67688
rect 31772 67630 32463 67632
rect 31772 67628 31778 67630
rect 32397 67627 32463 67630
rect 2606 67488 2922 67489
rect 2606 67424 2612 67488
rect 2676 67424 2692 67488
rect 2756 67424 2772 67488
rect 2836 67424 2852 67488
rect 2916 67424 2922 67488
rect 2606 67423 2922 67424
rect 7606 67488 7922 67489
rect 7606 67424 7612 67488
rect 7676 67424 7692 67488
rect 7756 67424 7772 67488
rect 7836 67424 7852 67488
rect 7916 67424 7922 67488
rect 7606 67423 7922 67424
rect 12606 67488 12922 67489
rect 12606 67424 12612 67488
rect 12676 67424 12692 67488
rect 12756 67424 12772 67488
rect 12836 67424 12852 67488
rect 12916 67424 12922 67488
rect 12606 67423 12922 67424
rect 17606 67488 17922 67489
rect 17606 67424 17612 67488
rect 17676 67424 17692 67488
rect 17756 67424 17772 67488
rect 17836 67424 17852 67488
rect 17916 67424 17922 67488
rect 17606 67423 17922 67424
rect 22606 67488 22922 67489
rect 22606 67424 22612 67488
rect 22676 67424 22692 67488
rect 22756 67424 22772 67488
rect 22836 67424 22852 67488
rect 22916 67424 22922 67488
rect 22606 67423 22922 67424
rect 27606 67488 27922 67489
rect 27606 67424 27612 67488
rect 27676 67424 27692 67488
rect 27756 67424 27772 67488
rect 27836 67424 27852 67488
rect 27916 67424 27922 67488
rect 27606 67423 27922 67424
rect 32606 67488 32922 67489
rect 32606 67424 32612 67488
rect 32676 67424 32692 67488
rect 32756 67424 32772 67488
rect 32836 67424 32852 67488
rect 32916 67424 32922 67488
rect 32606 67423 32922 67424
rect 37606 67488 37922 67489
rect 37606 67424 37612 67488
rect 37676 67424 37692 67488
rect 37756 67424 37772 67488
rect 37836 67424 37852 67488
rect 37916 67424 37922 67488
rect 37606 67423 37922 67424
rect 1946 66944 2262 66945
rect 1946 66880 1952 66944
rect 2016 66880 2032 66944
rect 2096 66880 2112 66944
rect 2176 66880 2192 66944
rect 2256 66880 2262 66944
rect 1946 66879 2262 66880
rect 6946 66944 7262 66945
rect 6946 66880 6952 66944
rect 7016 66880 7032 66944
rect 7096 66880 7112 66944
rect 7176 66880 7192 66944
rect 7256 66880 7262 66944
rect 6946 66879 7262 66880
rect 11946 66944 12262 66945
rect 11946 66880 11952 66944
rect 12016 66880 12032 66944
rect 12096 66880 12112 66944
rect 12176 66880 12192 66944
rect 12256 66880 12262 66944
rect 11946 66879 12262 66880
rect 16946 66944 17262 66945
rect 16946 66880 16952 66944
rect 17016 66880 17032 66944
rect 17096 66880 17112 66944
rect 17176 66880 17192 66944
rect 17256 66880 17262 66944
rect 16946 66879 17262 66880
rect 21946 66944 22262 66945
rect 21946 66880 21952 66944
rect 22016 66880 22032 66944
rect 22096 66880 22112 66944
rect 22176 66880 22192 66944
rect 22256 66880 22262 66944
rect 21946 66879 22262 66880
rect 26946 66944 27262 66945
rect 26946 66880 26952 66944
rect 27016 66880 27032 66944
rect 27096 66880 27112 66944
rect 27176 66880 27192 66944
rect 27256 66880 27262 66944
rect 26946 66879 27262 66880
rect 31946 66944 32262 66945
rect 31946 66880 31952 66944
rect 32016 66880 32032 66944
rect 32096 66880 32112 66944
rect 32176 66880 32192 66944
rect 32256 66880 32262 66944
rect 31946 66879 32262 66880
rect 36946 66944 37262 66945
rect 36946 66880 36952 66944
rect 37016 66880 37032 66944
rect 37096 66880 37112 66944
rect 37176 66880 37192 66944
rect 37256 66880 37262 66944
rect 36946 66879 37262 66880
rect 2606 66400 2922 66401
rect 2606 66336 2612 66400
rect 2676 66336 2692 66400
rect 2756 66336 2772 66400
rect 2836 66336 2852 66400
rect 2916 66336 2922 66400
rect 2606 66335 2922 66336
rect 7606 66400 7922 66401
rect 7606 66336 7612 66400
rect 7676 66336 7692 66400
rect 7756 66336 7772 66400
rect 7836 66336 7852 66400
rect 7916 66336 7922 66400
rect 7606 66335 7922 66336
rect 12606 66400 12922 66401
rect 12606 66336 12612 66400
rect 12676 66336 12692 66400
rect 12756 66336 12772 66400
rect 12836 66336 12852 66400
rect 12916 66336 12922 66400
rect 12606 66335 12922 66336
rect 17606 66400 17922 66401
rect 17606 66336 17612 66400
rect 17676 66336 17692 66400
rect 17756 66336 17772 66400
rect 17836 66336 17852 66400
rect 17916 66336 17922 66400
rect 17606 66335 17922 66336
rect 22606 66400 22922 66401
rect 22606 66336 22612 66400
rect 22676 66336 22692 66400
rect 22756 66336 22772 66400
rect 22836 66336 22852 66400
rect 22916 66336 22922 66400
rect 22606 66335 22922 66336
rect 27606 66400 27922 66401
rect 27606 66336 27612 66400
rect 27676 66336 27692 66400
rect 27756 66336 27772 66400
rect 27836 66336 27852 66400
rect 27916 66336 27922 66400
rect 27606 66335 27922 66336
rect 32606 66400 32922 66401
rect 32606 66336 32612 66400
rect 32676 66336 32692 66400
rect 32756 66336 32772 66400
rect 32836 66336 32852 66400
rect 32916 66336 32922 66400
rect 32606 66335 32922 66336
rect 37606 66400 37922 66401
rect 37606 66336 37612 66400
rect 37676 66336 37692 66400
rect 37756 66336 37772 66400
rect 37836 66336 37852 66400
rect 37916 66336 37922 66400
rect 37606 66335 37922 66336
rect 1946 65856 2262 65857
rect 1946 65792 1952 65856
rect 2016 65792 2032 65856
rect 2096 65792 2112 65856
rect 2176 65792 2192 65856
rect 2256 65792 2262 65856
rect 1946 65791 2262 65792
rect 6946 65856 7262 65857
rect 6946 65792 6952 65856
rect 7016 65792 7032 65856
rect 7096 65792 7112 65856
rect 7176 65792 7192 65856
rect 7256 65792 7262 65856
rect 6946 65791 7262 65792
rect 11946 65856 12262 65857
rect 11946 65792 11952 65856
rect 12016 65792 12032 65856
rect 12096 65792 12112 65856
rect 12176 65792 12192 65856
rect 12256 65792 12262 65856
rect 11946 65791 12262 65792
rect 16946 65856 17262 65857
rect 16946 65792 16952 65856
rect 17016 65792 17032 65856
rect 17096 65792 17112 65856
rect 17176 65792 17192 65856
rect 17256 65792 17262 65856
rect 16946 65791 17262 65792
rect 21946 65856 22262 65857
rect 21946 65792 21952 65856
rect 22016 65792 22032 65856
rect 22096 65792 22112 65856
rect 22176 65792 22192 65856
rect 22256 65792 22262 65856
rect 21946 65791 22262 65792
rect 26946 65856 27262 65857
rect 26946 65792 26952 65856
rect 27016 65792 27032 65856
rect 27096 65792 27112 65856
rect 27176 65792 27192 65856
rect 27256 65792 27262 65856
rect 26946 65791 27262 65792
rect 31946 65856 32262 65857
rect 31946 65792 31952 65856
rect 32016 65792 32032 65856
rect 32096 65792 32112 65856
rect 32176 65792 32192 65856
rect 32256 65792 32262 65856
rect 31946 65791 32262 65792
rect 36946 65856 37262 65857
rect 36946 65792 36952 65856
rect 37016 65792 37032 65856
rect 37096 65792 37112 65856
rect 37176 65792 37192 65856
rect 37256 65792 37262 65856
rect 36946 65791 37262 65792
rect 2606 65312 2922 65313
rect 2606 65248 2612 65312
rect 2676 65248 2692 65312
rect 2756 65248 2772 65312
rect 2836 65248 2852 65312
rect 2916 65248 2922 65312
rect 2606 65247 2922 65248
rect 7606 65312 7922 65313
rect 7606 65248 7612 65312
rect 7676 65248 7692 65312
rect 7756 65248 7772 65312
rect 7836 65248 7852 65312
rect 7916 65248 7922 65312
rect 7606 65247 7922 65248
rect 12606 65312 12922 65313
rect 12606 65248 12612 65312
rect 12676 65248 12692 65312
rect 12756 65248 12772 65312
rect 12836 65248 12852 65312
rect 12916 65248 12922 65312
rect 12606 65247 12922 65248
rect 17606 65312 17922 65313
rect 17606 65248 17612 65312
rect 17676 65248 17692 65312
rect 17756 65248 17772 65312
rect 17836 65248 17852 65312
rect 17916 65248 17922 65312
rect 17606 65247 17922 65248
rect 22606 65312 22922 65313
rect 22606 65248 22612 65312
rect 22676 65248 22692 65312
rect 22756 65248 22772 65312
rect 22836 65248 22852 65312
rect 22916 65248 22922 65312
rect 22606 65247 22922 65248
rect 27606 65312 27922 65313
rect 27606 65248 27612 65312
rect 27676 65248 27692 65312
rect 27756 65248 27772 65312
rect 27836 65248 27852 65312
rect 27916 65248 27922 65312
rect 27606 65247 27922 65248
rect 32606 65312 32922 65313
rect 32606 65248 32612 65312
rect 32676 65248 32692 65312
rect 32756 65248 32772 65312
rect 32836 65248 32852 65312
rect 32916 65248 32922 65312
rect 32606 65247 32922 65248
rect 37606 65312 37922 65313
rect 37606 65248 37612 65312
rect 37676 65248 37692 65312
rect 37756 65248 37772 65312
rect 37836 65248 37852 65312
rect 37916 65248 37922 65312
rect 37606 65247 37922 65248
rect 1946 64768 2262 64769
rect 1946 64704 1952 64768
rect 2016 64704 2032 64768
rect 2096 64704 2112 64768
rect 2176 64704 2192 64768
rect 2256 64704 2262 64768
rect 1946 64703 2262 64704
rect 6946 64768 7262 64769
rect 6946 64704 6952 64768
rect 7016 64704 7032 64768
rect 7096 64704 7112 64768
rect 7176 64704 7192 64768
rect 7256 64704 7262 64768
rect 6946 64703 7262 64704
rect 11946 64768 12262 64769
rect 11946 64704 11952 64768
rect 12016 64704 12032 64768
rect 12096 64704 12112 64768
rect 12176 64704 12192 64768
rect 12256 64704 12262 64768
rect 11946 64703 12262 64704
rect 16946 64768 17262 64769
rect 16946 64704 16952 64768
rect 17016 64704 17032 64768
rect 17096 64704 17112 64768
rect 17176 64704 17192 64768
rect 17256 64704 17262 64768
rect 16946 64703 17262 64704
rect 21946 64768 22262 64769
rect 21946 64704 21952 64768
rect 22016 64704 22032 64768
rect 22096 64704 22112 64768
rect 22176 64704 22192 64768
rect 22256 64704 22262 64768
rect 21946 64703 22262 64704
rect 26946 64768 27262 64769
rect 26946 64704 26952 64768
rect 27016 64704 27032 64768
rect 27096 64704 27112 64768
rect 27176 64704 27192 64768
rect 27256 64704 27262 64768
rect 26946 64703 27262 64704
rect 31946 64768 32262 64769
rect 31946 64704 31952 64768
rect 32016 64704 32032 64768
rect 32096 64704 32112 64768
rect 32176 64704 32192 64768
rect 32256 64704 32262 64768
rect 31946 64703 32262 64704
rect 36946 64768 37262 64769
rect 36946 64704 36952 64768
rect 37016 64704 37032 64768
rect 37096 64704 37112 64768
rect 37176 64704 37192 64768
rect 37256 64704 37262 64768
rect 36946 64703 37262 64704
rect 2606 64224 2922 64225
rect 2606 64160 2612 64224
rect 2676 64160 2692 64224
rect 2756 64160 2772 64224
rect 2836 64160 2852 64224
rect 2916 64160 2922 64224
rect 2606 64159 2922 64160
rect 7606 64224 7922 64225
rect 7606 64160 7612 64224
rect 7676 64160 7692 64224
rect 7756 64160 7772 64224
rect 7836 64160 7852 64224
rect 7916 64160 7922 64224
rect 7606 64159 7922 64160
rect 12606 64224 12922 64225
rect 12606 64160 12612 64224
rect 12676 64160 12692 64224
rect 12756 64160 12772 64224
rect 12836 64160 12852 64224
rect 12916 64160 12922 64224
rect 12606 64159 12922 64160
rect 17606 64224 17922 64225
rect 17606 64160 17612 64224
rect 17676 64160 17692 64224
rect 17756 64160 17772 64224
rect 17836 64160 17852 64224
rect 17916 64160 17922 64224
rect 17606 64159 17922 64160
rect 22606 64224 22922 64225
rect 22606 64160 22612 64224
rect 22676 64160 22692 64224
rect 22756 64160 22772 64224
rect 22836 64160 22852 64224
rect 22916 64160 22922 64224
rect 22606 64159 22922 64160
rect 27606 64224 27922 64225
rect 27606 64160 27612 64224
rect 27676 64160 27692 64224
rect 27756 64160 27772 64224
rect 27836 64160 27852 64224
rect 27916 64160 27922 64224
rect 27606 64159 27922 64160
rect 32606 64224 32922 64225
rect 32606 64160 32612 64224
rect 32676 64160 32692 64224
rect 32756 64160 32772 64224
rect 32836 64160 32852 64224
rect 32916 64160 32922 64224
rect 32606 64159 32922 64160
rect 37606 64224 37922 64225
rect 37606 64160 37612 64224
rect 37676 64160 37692 64224
rect 37756 64160 37772 64224
rect 37836 64160 37852 64224
rect 37916 64160 37922 64224
rect 37606 64159 37922 64160
rect 1946 63680 2262 63681
rect 1946 63616 1952 63680
rect 2016 63616 2032 63680
rect 2096 63616 2112 63680
rect 2176 63616 2192 63680
rect 2256 63616 2262 63680
rect 1946 63615 2262 63616
rect 6946 63680 7262 63681
rect 6946 63616 6952 63680
rect 7016 63616 7032 63680
rect 7096 63616 7112 63680
rect 7176 63616 7192 63680
rect 7256 63616 7262 63680
rect 6946 63615 7262 63616
rect 11946 63680 12262 63681
rect 11946 63616 11952 63680
rect 12016 63616 12032 63680
rect 12096 63616 12112 63680
rect 12176 63616 12192 63680
rect 12256 63616 12262 63680
rect 11946 63615 12262 63616
rect 16946 63680 17262 63681
rect 16946 63616 16952 63680
rect 17016 63616 17032 63680
rect 17096 63616 17112 63680
rect 17176 63616 17192 63680
rect 17256 63616 17262 63680
rect 16946 63615 17262 63616
rect 21946 63680 22262 63681
rect 21946 63616 21952 63680
rect 22016 63616 22032 63680
rect 22096 63616 22112 63680
rect 22176 63616 22192 63680
rect 22256 63616 22262 63680
rect 21946 63615 22262 63616
rect 26946 63680 27262 63681
rect 26946 63616 26952 63680
rect 27016 63616 27032 63680
rect 27096 63616 27112 63680
rect 27176 63616 27192 63680
rect 27256 63616 27262 63680
rect 26946 63615 27262 63616
rect 31946 63680 32262 63681
rect 31946 63616 31952 63680
rect 32016 63616 32032 63680
rect 32096 63616 32112 63680
rect 32176 63616 32192 63680
rect 32256 63616 32262 63680
rect 31946 63615 32262 63616
rect 36946 63680 37262 63681
rect 36946 63616 36952 63680
rect 37016 63616 37032 63680
rect 37096 63616 37112 63680
rect 37176 63616 37192 63680
rect 37256 63616 37262 63680
rect 36946 63615 37262 63616
rect 2606 63136 2922 63137
rect 2606 63072 2612 63136
rect 2676 63072 2692 63136
rect 2756 63072 2772 63136
rect 2836 63072 2852 63136
rect 2916 63072 2922 63136
rect 2606 63071 2922 63072
rect 7606 63136 7922 63137
rect 7606 63072 7612 63136
rect 7676 63072 7692 63136
rect 7756 63072 7772 63136
rect 7836 63072 7852 63136
rect 7916 63072 7922 63136
rect 7606 63071 7922 63072
rect 12606 63136 12922 63137
rect 12606 63072 12612 63136
rect 12676 63072 12692 63136
rect 12756 63072 12772 63136
rect 12836 63072 12852 63136
rect 12916 63072 12922 63136
rect 12606 63071 12922 63072
rect 17606 63136 17922 63137
rect 17606 63072 17612 63136
rect 17676 63072 17692 63136
rect 17756 63072 17772 63136
rect 17836 63072 17852 63136
rect 17916 63072 17922 63136
rect 17606 63071 17922 63072
rect 22606 63136 22922 63137
rect 22606 63072 22612 63136
rect 22676 63072 22692 63136
rect 22756 63072 22772 63136
rect 22836 63072 22852 63136
rect 22916 63072 22922 63136
rect 22606 63071 22922 63072
rect 27606 63136 27922 63137
rect 27606 63072 27612 63136
rect 27676 63072 27692 63136
rect 27756 63072 27772 63136
rect 27836 63072 27852 63136
rect 27916 63072 27922 63136
rect 27606 63071 27922 63072
rect 32606 63136 32922 63137
rect 32606 63072 32612 63136
rect 32676 63072 32692 63136
rect 32756 63072 32772 63136
rect 32836 63072 32852 63136
rect 32916 63072 32922 63136
rect 32606 63071 32922 63072
rect 37606 63136 37922 63137
rect 37606 63072 37612 63136
rect 37676 63072 37692 63136
rect 37756 63072 37772 63136
rect 37836 63072 37852 63136
rect 37916 63072 37922 63136
rect 37606 63071 37922 63072
rect 1946 62592 2262 62593
rect 1946 62528 1952 62592
rect 2016 62528 2032 62592
rect 2096 62528 2112 62592
rect 2176 62528 2192 62592
rect 2256 62528 2262 62592
rect 1946 62527 2262 62528
rect 6946 62592 7262 62593
rect 6946 62528 6952 62592
rect 7016 62528 7032 62592
rect 7096 62528 7112 62592
rect 7176 62528 7192 62592
rect 7256 62528 7262 62592
rect 6946 62527 7262 62528
rect 11946 62592 12262 62593
rect 11946 62528 11952 62592
rect 12016 62528 12032 62592
rect 12096 62528 12112 62592
rect 12176 62528 12192 62592
rect 12256 62528 12262 62592
rect 11946 62527 12262 62528
rect 16946 62592 17262 62593
rect 16946 62528 16952 62592
rect 17016 62528 17032 62592
rect 17096 62528 17112 62592
rect 17176 62528 17192 62592
rect 17256 62528 17262 62592
rect 16946 62527 17262 62528
rect 21946 62592 22262 62593
rect 21946 62528 21952 62592
rect 22016 62528 22032 62592
rect 22096 62528 22112 62592
rect 22176 62528 22192 62592
rect 22256 62528 22262 62592
rect 21946 62527 22262 62528
rect 26946 62592 27262 62593
rect 26946 62528 26952 62592
rect 27016 62528 27032 62592
rect 27096 62528 27112 62592
rect 27176 62528 27192 62592
rect 27256 62528 27262 62592
rect 26946 62527 27262 62528
rect 31946 62592 32262 62593
rect 31946 62528 31952 62592
rect 32016 62528 32032 62592
rect 32096 62528 32112 62592
rect 32176 62528 32192 62592
rect 32256 62528 32262 62592
rect 31946 62527 32262 62528
rect 36946 62592 37262 62593
rect 36946 62528 36952 62592
rect 37016 62528 37032 62592
rect 37096 62528 37112 62592
rect 37176 62528 37192 62592
rect 37256 62528 37262 62592
rect 36946 62527 37262 62528
rect 2606 62048 2922 62049
rect 2606 61984 2612 62048
rect 2676 61984 2692 62048
rect 2756 61984 2772 62048
rect 2836 61984 2852 62048
rect 2916 61984 2922 62048
rect 2606 61983 2922 61984
rect 7606 62048 7922 62049
rect 7606 61984 7612 62048
rect 7676 61984 7692 62048
rect 7756 61984 7772 62048
rect 7836 61984 7852 62048
rect 7916 61984 7922 62048
rect 7606 61983 7922 61984
rect 12606 62048 12922 62049
rect 12606 61984 12612 62048
rect 12676 61984 12692 62048
rect 12756 61984 12772 62048
rect 12836 61984 12852 62048
rect 12916 61984 12922 62048
rect 12606 61983 12922 61984
rect 17606 62048 17922 62049
rect 17606 61984 17612 62048
rect 17676 61984 17692 62048
rect 17756 61984 17772 62048
rect 17836 61984 17852 62048
rect 17916 61984 17922 62048
rect 17606 61983 17922 61984
rect 22606 62048 22922 62049
rect 22606 61984 22612 62048
rect 22676 61984 22692 62048
rect 22756 61984 22772 62048
rect 22836 61984 22852 62048
rect 22916 61984 22922 62048
rect 22606 61983 22922 61984
rect 27606 62048 27922 62049
rect 27606 61984 27612 62048
rect 27676 61984 27692 62048
rect 27756 61984 27772 62048
rect 27836 61984 27852 62048
rect 27916 61984 27922 62048
rect 27606 61983 27922 61984
rect 32606 62048 32922 62049
rect 32606 61984 32612 62048
rect 32676 61984 32692 62048
rect 32756 61984 32772 62048
rect 32836 61984 32852 62048
rect 32916 61984 32922 62048
rect 32606 61983 32922 61984
rect 37606 62048 37922 62049
rect 37606 61984 37612 62048
rect 37676 61984 37692 62048
rect 37756 61984 37772 62048
rect 37836 61984 37852 62048
rect 37916 61984 37922 62048
rect 37606 61983 37922 61984
rect 1946 61504 2262 61505
rect 1946 61440 1952 61504
rect 2016 61440 2032 61504
rect 2096 61440 2112 61504
rect 2176 61440 2192 61504
rect 2256 61440 2262 61504
rect 1946 61439 2262 61440
rect 6946 61504 7262 61505
rect 6946 61440 6952 61504
rect 7016 61440 7032 61504
rect 7096 61440 7112 61504
rect 7176 61440 7192 61504
rect 7256 61440 7262 61504
rect 6946 61439 7262 61440
rect 11946 61504 12262 61505
rect 11946 61440 11952 61504
rect 12016 61440 12032 61504
rect 12096 61440 12112 61504
rect 12176 61440 12192 61504
rect 12256 61440 12262 61504
rect 11946 61439 12262 61440
rect 16946 61504 17262 61505
rect 16946 61440 16952 61504
rect 17016 61440 17032 61504
rect 17096 61440 17112 61504
rect 17176 61440 17192 61504
rect 17256 61440 17262 61504
rect 16946 61439 17262 61440
rect 21946 61504 22262 61505
rect 21946 61440 21952 61504
rect 22016 61440 22032 61504
rect 22096 61440 22112 61504
rect 22176 61440 22192 61504
rect 22256 61440 22262 61504
rect 21946 61439 22262 61440
rect 26946 61504 27262 61505
rect 26946 61440 26952 61504
rect 27016 61440 27032 61504
rect 27096 61440 27112 61504
rect 27176 61440 27192 61504
rect 27256 61440 27262 61504
rect 26946 61439 27262 61440
rect 31946 61504 32262 61505
rect 31946 61440 31952 61504
rect 32016 61440 32032 61504
rect 32096 61440 32112 61504
rect 32176 61440 32192 61504
rect 32256 61440 32262 61504
rect 31946 61439 32262 61440
rect 36946 61504 37262 61505
rect 36946 61440 36952 61504
rect 37016 61440 37032 61504
rect 37096 61440 37112 61504
rect 37176 61440 37192 61504
rect 37256 61440 37262 61504
rect 36946 61439 37262 61440
rect 2606 60960 2922 60961
rect 2606 60896 2612 60960
rect 2676 60896 2692 60960
rect 2756 60896 2772 60960
rect 2836 60896 2852 60960
rect 2916 60896 2922 60960
rect 2606 60895 2922 60896
rect 7606 60960 7922 60961
rect 7606 60896 7612 60960
rect 7676 60896 7692 60960
rect 7756 60896 7772 60960
rect 7836 60896 7852 60960
rect 7916 60896 7922 60960
rect 7606 60895 7922 60896
rect 12606 60960 12922 60961
rect 12606 60896 12612 60960
rect 12676 60896 12692 60960
rect 12756 60896 12772 60960
rect 12836 60896 12852 60960
rect 12916 60896 12922 60960
rect 12606 60895 12922 60896
rect 17606 60960 17922 60961
rect 17606 60896 17612 60960
rect 17676 60896 17692 60960
rect 17756 60896 17772 60960
rect 17836 60896 17852 60960
rect 17916 60896 17922 60960
rect 17606 60895 17922 60896
rect 22606 60960 22922 60961
rect 22606 60896 22612 60960
rect 22676 60896 22692 60960
rect 22756 60896 22772 60960
rect 22836 60896 22852 60960
rect 22916 60896 22922 60960
rect 22606 60895 22922 60896
rect 27606 60960 27922 60961
rect 27606 60896 27612 60960
rect 27676 60896 27692 60960
rect 27756 60896 27772 60960
rect 27836 60896 27852 60960
rect 27916 60896 27922 60960
rect 27606 60895 27922 60896
rect 32606 60960 32922 60961
rect 32606 60896 32612 60960
rect 32676 60896 32692 60960
rect 32756 60896 32772 60960
rect 32836 60896 32852 60960
rect 32916 60896 32922 60960
rect 32606 60895 32922 60896
rect 37606 60960 37922 60961
rect 37606 60896 37612 60960
rect 37676 60896 37692 60960
rect 37756 60896 37772 60960
rect 37836 60896 37852 60960
rect 37916 60896 37922 60960
rect 37606 60895 37922 60896
rect 1946 60416 2262 60417
rect 1946 60352 1952 60416
rect 2016 60352 2032 60416
rect 2096 60352 2112 60416
rect 2176 60352 2192 60416
rect 2256 60352 2262 60416
rect 1946 60351 2262 60352
rect 6946 60416 7262 60417
rect 6946 60352 6952 60416
rect 7016 60352 7032 60416
rect 7096 60352 7112 60416
rect 7176 60352 7192 60416
rect 7256 60352 7262 60416
rect 6946 60351 7262 60352
rect 11946 60416 12262 60417
rect 11946 60352 11952 60416
rect 12016 60352 12032 60416
rect 12096 60352 12112 60416
rect 12176 60352 12192 60416
rect 12256 60352 12262 60416
rect 11946 60351 12262 60352
rect 16946 60416 17262 60417
rect 16946 60352 16952 60416
rect 17016 60352 17032 60416
rect 17096 60352 17112 60416
rect 17176 60352 17192 60416
rect 17256 60352 17262 60416
rect 16946 60351 17262 60352
rect 21946 60416 22262 60417
rect 21946 60352 21952 60416
rect 22016 60352 22032 60416
rect 22096 60352 22112 60416
rect 22176 60352 22192 60416
rect 22256 60352 22262 60416
rect 21946 60351 22262 60352
rect 26946 60416 27262 60417
rect 26946 60352 26952 60416
rect 27016 60352 27032 60416
rect 27096 60352 27112 60416
rect 27176 60352 27192 60416
rect 27256 60352 27262 60416
rect 26946 60351 27262 60352
rect 31946 60416 32262 60417
rect 31946 60352 31952 60416
rect 32016 60352 32032 60416
rect 32096 60352 32112 60416
rect 32176 60352 32192 60416
rect 32256 60352 32262 60416
rect 31946 60351 32262 60352
rect 36946 60416 37262 60417
rect 36946 60352 36952 60416
rect 37016 60352 37032 60416
rect 37096 60352 37112 60416
rect 37176 60352 37192 60416
rect 37256 60352 37262 60416
rect 36946 60351 37262 60352
rect 2606 59872 2922 59873
rect 2606 59808 2612 59872
rect 2676 59808 2692 59872
rect 2756 59808 2772 59872
rect 2836 59808 2852 59872
rect 2916 59808 2922 59872
rect 2606 59807 2922 59808
rect 7606 59872 7922 59873
rect 7606 59808 7612 59872
rect 7676 59808 7692 59872
rect 7756 59808 7772 59872
rect 7836 59808 7852 59872
rect 7916 59808 7922 59872
rect 7606 59807 7922 59808
rect 12606 59872 12922 59873
rect 12606 59808 12612 59872
rect 12676 59808 12692 59872
rect 12756 59808 12772 59872
rect 12836 59808 12852 59872
rect 12916 59808 12922 59872
rect 12606 59807 12922 59808
rect 17606 59872 17922 59873
rect 17606 59808 17612 59872
rect 17676 59808 17692 59872
rect 17756 59808 17772 59872
rect 17836 59808 17852 59872
rect 17916 59808 17922 59872
rect 17606 59807 17922 59808
rect 22606 59872 22922 59873
rect 22606 59808 22612 59872
rect 22676 59808 22692 59872
rect 22756 59808 22772 59872
rect 22836 59808 22852 59872
rect 22916 59808 22922 59872
rect 22606 59807 22922 59808
rect 27606 59872 27922 59873
rect 27606 59808 27612 59872
rect 27676 59808 27692 59872
rect 27756 59808 27772 59872
rect 27836 59808 27852 59872
rect 27916 59808 27922 59872
rect 27606 59807 27922 59808
rect 32606 59872 32922 59873
rect 32606 59808 32612 59872
rect 32676 59808 32692 59872
rect 32756 59808 32772 59872
rect 32836 59808 32852 59872
rect 32916 59808 32922 59872
rect 32606 59807 32922 59808
rect 37606 59872 37922 59873
rect 37606 59808 37612 59872
rect 37676 59808 37692 59872
rect 37756 59808 37772 59872
rect 37836 59808 37852 59872
rect 37916 59808 37922 59872
rect 37606 59807 37922 59808
rect 1946 59328 2262 59329
rect 1946 59264 1952 59328
rect 2016 59264 2032 59328
rect 2096 59264 2112 59328
rect 2176 59264 2192 59328
rect 2256 59264 2262 59328
rect 1946 59263 2262 59264
rect 6946 59328 7262 59329
rect 6946 59264 6952 59328
rect 7016 59264 7032 59328
rect 7096 59264 7112 59328
rect 7176 59264 7192 59328
rect 7256 59264 7262 59328
rect 6946 59263 7262 59264
rect 11946 59328 12262 59329
rect 11946 59264 11952 59328
rect 12016 59264 12032 59328
rect 12096 59264 12112 59328
rect 12176 59264 12192 59328
rect 12256 59264 12262 59328
rect 11946 59263 12262 59264
rect 16946 59328 17262 59329
rect 16946 59264 16952 59328
rect 17016 59264 17032 59328
rect 17096 59264 17112 59328
rect 17176 59264 17192 59328
rect 17256 59264 17262 59328
rect 16946 59263 17262 59264
rect 21946 59328 22262 59329
rect 21946 59264 21952 59328
rect 22016 59264 22032 59328
rect 22096 59264 22112 59328
rect 22176 59264 22192 59328
rect 22256 59264 22262 59328
rect 21946 59263 22262 59264
rect 26946 59328 27262 59329
rect 26946 59264 26952 59328
rect 27016 59264 27032 59328
rect 27096 59264 27112 59328
rect 27176 59264 27192 59328
rect 27256 59264 27262 59328
rect 26946 59263 27262 59264
rect 31946 59328 32262 59329
rect 31946 59264 31952 59328
rect 32016 59264 32032 59328
rect 32096 59264 32112 59328
rect 32176 59264 32192 59328
rect 32256 59264 32262 59328
rect 31946 59263 32262 59264
rect 36946 59328 37262 59329
rect 36946 59264 36952 59328
rect 37016 59264 37032 59328
rect 37096 59264 37112 59328
rect 37176 59264 37192 59328
rect 37256 59264 37262 59328
rect 36946 59263 37262 59264
rect 2606 58784 2922 58785
rect 2606 58720 2612 58784
rect 2676 58720 2692 58784
rect 2756 58720 2772 58784
rect 2836 58720 2852 58784
rect 2916 58720 2922 58784
rect 2606 58719 2922 58720
rect 7606 58784 7922 58785
rect 7606 58720 7612 58784
rect 7676 58720 7692 58784
rect 7756 58720 7772 58784
rect 7836 58720 7852 58784
rect 7916 58720 7922 58784
rect 7606 58719 7922 58720
rect 12606 58784 12922 58785
rect 12606 58720 12612 58784
rect 12676 58720 12692 58784
rect 12756 58720 12772 58784
rect 12836 58720 12852 58784
rect 12916 58720 12922 58784
rect 12606 58719 12922 58720
rect 17606 58784 17922 58785
rect 17606 58720 17612 58784
rect 17676 58720 17692 58784
rect 17756 58720 17772 58784
rect 17836 58720 17852 58784
rect 17916 58720 17922 58784
rect 17606 58719 17922 58720
rect 22606 58784 22922 58785
rect 22606 58720 22612 58784
rect 22676 58720 22692 58784
rect 22756 58720 22772 58784
rect 22836 58720 22852 58784
rect 22916 58720 22922 58784
rect 22606 58719 22922 58720
rect 27606 58784 27922 58785
rect 27606 58720 27612 58784
rect 27676 58720 27692 58784
rect 27756 58720 27772 58784
rect 27836 58720 27852 58784
rect 27916 58720 27922 58784
rect 27606 58719 27922 58720
rect 32606 58784 32922 58785
rect 32606 58720 32612 58784
rect 32676 58720 32692 58784
rect 32756 58720 32772 58784
rect 32836 58720 32852 58784
rect 32916 58720 32922 58784
rect 32606 58719 32922 58720
rect 37606 58784 37922 58785
rect 37606 58720 37612 58784
rect 37676 58720 37692 58784
rect 37756 58720 37772 58784
rect 37836 58720 37852 58784
rect 37916 58720 37922 58784
rect 37606 58719 37922 58720
rect 33225 58308 33291 58309
rect 33174 58306 33180 58308
rect 33134 58246 33180 58306
rect 33244 58304 33291 58308
rect 33286 58248 33291 58304
rect 33174 58244 33180 58246
rect 33244 58244 33291 58248
rect 33225 58243 33291 58244
rect 1946 58240 2262 58241
rect 1946 58176 1952 58240
rect 2016 58176 2032 58240
rect 2096 58176 2112 58240
rect 2176 58176 2192 58240
rect 2256 58176 2262 58240
rect 1946 58175 2262 58176
rect 6946 58240 7262 58241
rect 6946 58176 6952 58240
rect 7016 58176 7032 58240
rect 7096 58176 7112 58240
rect 7176 58176 7192 58240
rect 7256 58176 7262 58240
rect 6946 58175 7262 58176
rect 11946 58240 12262 58241
rect 11946 58176 11952 58240
rect 12016 58176 12032 58240
rect 12096 58176 12112 58240
rect 12176 58176 12192 58240
rect 12256 58176 12262 58240
rect 11946 58175 12262 58176
rect 16946 58240 17262 58241
rect 16946 58176 16952 58240
rect 17016 58176 17032 58240
rect 17096 58176 17112 58240
rect 17176 58176 17192 58240
rect 17256 58176 17262 58240
rect 16946 58175 17262 58176
rect 21946 58240 22262 58241
rect 21946 58176 21952 58240
rect 22016 58176 22032 58240
rect 22096 58176 22112 58240
rect 22176 58176 22192 58240
rect 22256 58176 22262 58240
rect 21946 58175 22262 58176
rect 26946 58240 27262 58241
rect 26946 58176 26952 58240
rect 27016 58176 27032 58240
rect 27096 58176 27112 58240
rect 27176 58176 27192 58240
rect 27256 58176 27262 58240
rect 26946 58175 27262 58176
rect 31946 58240 32262 58241
rect 31946 58176 31952 58240
rect 32016 58176 32032 58240
rect 32096 58176 32112 58240
rect 32176 58176 32192 58240
rect 32256 58176 32262 58240
rect 31946 58175 32262 58176
rect 36946 58240 37262 58241
rect 36946 58176 36952 58240
rect 37016 58176 37032 58240
rect 37096 58176 37112 58240
rect 37176 58176 37192 58240
rect 37256 58176 37262 58240
rect 36946 58175 37262 58176
rect 2606 57696 2922 57697
rect 2606 57632 2612 57696
rect 2676 57632 2692 57696
rect 2756 57632 2772 57696
rect 2836 57632 2852 57696
rect 2916 57632 2922 57696
rect 2606 57631 2922 57632
rect 7606 57696 7922 57697
rect 7606 57632 7612 57696
rect 7676 57632 7692 57696
rect 7756 57632 7772 57696
rect 7836 57632 7852 57696
rect 7916 57632 7922 57696
rect 7606 57631 7922 57632
rect 12606 57696 12922 57697
rect 12606 57632 12612 57696
rect 12676 57632 12692 57696
rect 12756 57632 12772 57696
rect 12836 57632 12852 57696
rect 12916 57632 12922 57696
rect 12606 57631 12922 57632
rect 17606 57696 17922 57697
rect 17606 57632 17612 57696
rect 17676 57632 17692 57696
rect 17756 57632 17772 57696
rect 17836 57632 17852 57696
rect 17916 57632 17922 57696
rect 17606 57631 17922 57632
rect 22606 57696 22922 57697
rect 22606 57632 22612 57696
rect 22676 57632 22692 57696
rect 22756 57632 22772 57696
rect 22836 57632 22852 57696
rect 22916 57632 22922 57696
rect 22606 57631 22922 57632
rect 27606 57696 27922 57697
rect 27606 57632 27612 57696
rect 27676 57632 27692 57696
rect 27756 57632 27772 57696
rect 27836 57632 27852 57696
rect 27916 57632 27922 57696
rect 27606 57631 27922 57632
rect 32606 57696 32922 57697
rect 32606 57632 32612 57696
rect 32676 57632 32692 57696
rect 32756 57632 32772 57696
rect 32836 57632 32852 57696
rect 32916 57632 32922 57696
rect 32606 57631 32922 57632
rect 37606 57696 37922 57697
rect 37606 57632 37612 57696
rect 37676 57632 37692 57696
rect 37756 57632 37772 57696
rect 37836 57632 37852 57696
rect 37916 57632 37922 57696
rect 37606 57631 37922 57632
rect 1946 57152 2262 57153
rect 1946 57088 1952 57152
rect 2016 57088 2032 57152
rect 2096 57088 2112 57152
rect 2176 57088 2192 57152
rect 2256 57088 2262 57152
rect 1946 57087 2262 57088
rect 6946 57152 7262 57153
rect 6946 57088 6952 57152
rect 7016 57088 7032 57152
rect 7096 57088 7112 57152
rect 7176 57088 7192 57152
rect 7256 57088 7262 57152
rect 6946 57087 7262 57088
rect 11946 57152 12262 57153
rect 11946 57088 11952 57152
rect 12016 57088 12032 57152
rect 12096 57088 12112 57152
rect 12176 57088 12192 57152
rect 12256 57088 12262 57152
rect 11946 57087 12262 57088
rect 16946 57152 17262 57153
rect 16946 57088 16952 57152
rect 17016 57088 17032 57152
rect 17096 57088 17112 57152
rect 17176 57088 17192 57152
rect 17256 57088 17262 57152
rect 16946 57087 17262 57088
rect 21946 57152 22262 57153
rect 21946 57088 21952 57152
rect 22016 57088 22032 57152
rect 22096 57088 22112 57152
rect 22176 57088 22192 57152
rect 22256 57088 22262 57152
rect 21946 57087 22262 57088
rect 26946 57152 27262 57153
rect 26946 57088 26952 57152
rect 27016 57088 27032 57152
rect 27096 57088 27112 57152
rect 27176 57088 27192 57152
rect 27256 57088 27262 57152
rect 26946 57087 27262 57088
rect 31946 57152 32262 57153
rect 31946 57088 31952 57152
rect 32016 57088 32032 57152
rect 32096 57088 32112 57152
rect 32176 57088 32192 57152
rect 32256 57088 32262 57152
rect 31946 57087 32262 57088
rect 36946 57152 37262 57153
rect 36946 57088 36952 57152
rect 37016 57088 37032 57152
rect 37096 57088 37112 57152
rect 37176 57088 37192 57152
rect 37256 57088 37262 57152
rect 36946 57087 37262 57088
rect 2606 56608 2922 56609
rect 2606 56544 2612 56608
rect 2676 56544 2692 56608
rect 2756 56544 2772 56608
rect 2836 56544 2852 56608
rect 2916 56544 2922 56608
rect 2606 56543 2922 56544
rect 7606 56608 7922 56609
rect 7606 56544 7612 56608
rect 7676 56544 7692 56608
rect 7756 56544 7772 56608
rect 7836 56544 7852 56608
rect 7916 56544 7922 56608
rect 7606 56543 7922 56544
rect 12606 56608 12922 56609
rect 12606 56544 12612 56608
rect 12676 56544 12692 56608
rect 12756 56544 12772 56608
rect 12836 56544 12852 56608
rect 12916 56544 12922 56608
rect 12606 56543 12922 56544
rect 17606 56608 17922 56609
rect 17606 56544 17612 56608
rect 17676 56544 17692 56608
rect 17756 56544 17772 56608
rect 17836 56544 17852 56608
rect 17916 56544 17922 56608
rect 17606 56543 17922 56544
rect 22606 56608 22922 56609
rect 22606 56544 22612 56608
rect 22676 56544 22692 56608
rect 22756 56544 22772 56608
rect 22836 56544 22852 56608
rect 22916 56544 22922 56608
rect 22606 56543 22922 56544
rect 27606 56608 27922 56609
rect 27606 56544 27612 56608
rect 27676 56544 27692 56608
rect 27756 56544 27772 56608
rect 27836 56544 27852 56608
rect 27916 56544 27922 56608
rect 27606 56543 27922 56544
rect 32606 56608 32922 56609
rect 32606 56544 32612 56608
rect 32676 56544 32692 56608
rect 32756 56544 32772 56608
rect 32836 56544 32852 56608
rect 32916 56544 32922 56608
rect 32606 56543 32922 56544
rect 37606 56608 37922 56609
rect 37606 56544 37612 56608
rect 37676 56544 37692 56608
rect 37756 56544 37772 56608
rect 37836 56544 37852 56608
rect 37916 56544 37922 56608
rect 37606 56543 37922 56544
rect 1946 56064 2262 56065
rect 1946 56000 1952 56064
rect 2016 56000 2032 56064
rect 2096 56000 2112 56064
rect 2176 56000 2192 56064
rect 2256 56000 2262 56064
rect 1946 55999 2262 56000
rect 6946 56064 7262 56065
rect 6946 56000 6952 56064
rect 7016 56000 7032 56064
rect 7096 56000 7112 56064
rect 7176 56000 7192 56064
rect 7256 56000 7262 56064
rect 6946 55999 7262 56000
rect 11946 56064 12262 56065
rect 11946 56000 11952 56064
rect 12016 56000 12032 56064
rect 12096 56000 12112 56064
rect 12176 56000 12192 56064
rect 12256 56000 12262 56064
rect 11946 55999 12262 56000
rect 16946 56064 17262 56065
rect 16946 56000 16952 56064
rect 17016 56000 17032 56064
rect 17096 56000 17112 56064
rect 17176 56000 17192 56064
rect 17256 56000 17262 56064
rect 16946 55999 17262 56000
rect 21946 56064 22262 56065
rect 21946 56000 21952 56064
rect 22016 56000 22032 56064
rect 22096 56000 22112 56064
rect 22176 56000 22192 56064
rect 22256 56000 22262 56064
rect 21946 55999 22262 56000
rect 26946 56064 27262 56065
rect 26946 56000 26952 56064
rect 27016 56000 27032 56064
rect 27096 56000 27112 56064
rect 27176 56000 27192 56064
rect 27256 56000 27262 56064
rect 26946 55999 27262 56000
rect 31946 56064 32262 56065
rect 31946 56000 31952 56064
rect 32016 56000 32032 56064
rect 32096 56000 32112 56064
rect 32176 56000 32192 56064
rect 32256 56000 32262 56064
rect 31946 55999 32262 56000
rect 36946 56064 37262 56065
rect 36946 56000 36952 56064
rect 37016 56000 37032 56064
rect 37096 56000 37112 56064
rect 37176 56000 37192 56064
rect 37256 56000 37262 56064
rect 36946 55999 37262 56000
rect 33869 55860 33935 55861
rect 33869 55856 33916 55860
rect 33980 55858 33986 55860
rect 33869 55800 33874 55856
rect 33869 55796 33916 55800
rect 33980 55798 34026 55858
rect 33980 55796 33986 55798
rect 33869 55795 33935 55796
rect 33501 55724 33567 55725
rect 33501 55720 33548 55724
rect 33612 55722 33618 55724
rect 33501 55664 33506 55720
rect 33501 55660 33548 55664
rect 33612 55662 33658 55722
rect 33612 55660 33618 55662
rect 33501 55659 33567 55660
rect 2606 55520 2922 55521
rect 2606 55456 2612 55520
rect 2676 55456 2692 55520
rect 2756 55456 2772 55520
rect 2836 55456 2852 55520
rect 2916 55456 2922 55520
rect 2606 55455 2922 55456
rect 7606 55520 7922 55521
rect 7606 55456 7612 55520
rect 7676 55456 7692 55520
rect 7756 55456 7772 55520
rect 7836 55456 7852 55520
rect 7916 55456 7922 55520
rect 7606 55455 7922 55456
rect 12606 55520 12922 55521
rect 12606 55456 12612 55520
rect 12676 55456 12692 55520
rect 12756 55456 12772 55520
rect 12836 55456 12852 55520
rect 12916 55456 12922 55520
rect 12606 55455 12922 55456
rect 17606 55520 17922 55521
rect 17606 55456 17612 55520
rect 17676 55456 17692 55520
rect 17756 55456 17772 55520
rect 17836 55456 17852 55520
rect 17916 55456 17922 55520
rect 17606 55455 17922 55456
rect 22606 55520 22922 55521
rect 22606 55456 22612 55520
rect 22676 55456 22692 55520
rect 22756 55456 22772 55520
rect 22836 55456 22852 55520
rect 22916 55456 22922 55520
rect 22606 55455 22922 55456
rect 27606 55520 27922 55521
rect 27606 55456 27612 55520
rect 27676 55456 27692 55520
rect 27756 55456 27772 55520
rect 27836 55456 27852 55520
rect 27916 55456 27922 55520
rect 27606 55455 27922 55456
rect 32606 55520 32922 55521
rect 32606 55456 32612 55520
rect 32676 55456 32692 55520
rect 32756 55456 32772 55520
rect 32836 55456 32852 55520
rect 32916 55456 32922 55520
rect 32606 55455 32922 55456
rect 37606 55520 37922 55521
rect 37606 55456 37612 55520
rect 37676 55456 37692 55520
rect 37756 55456 37772 55520
rect 37836 55456 37852 55520
rect 37916 55456 37922 55520
rect 37606 55455 37922 55456
rect 1946 54976 2262 54977
rect 1946 54912 1952 54976
rect 2016 54912 2032 54976
rect 2096 54912 2112 54976
rect 2176 54912 2192 54976
rect 2256 54912 2262 54976
rect 1946 54911 2262 54912
rect 6946 54976 7262 54977
rect 6946 54912 6952 54976
rect 7016 54912 7032 54976
rect 7096 54912 7112 54976
rect 7176 54912 7192 54976
rect 7256 54912 7262 54976
rect 6946 54911 7262 54912
rect 11946 54976 12262 54977
rect 11946 54912 11952 54976
rect 12016 54912 12032 54976
rect 12096 54912 12112 54976
rect 12176 54912 12192 54976
rect 12256 54912 12262 54976
rect 11946 54911 12262 54912
rect 16946 54976 17262 54977
rect 16946 54912 16952 54976
rect 17016 54912 17032 54976
rect 17096 54912 17112 54976
rect 17176 54912 17192 54976
rect 17256 54912 17262 54976
rect 16946 54911 17262 54912
rect 21946 54976 22262 54977
rect 21946 54912 21952 54976
rect 22016 54912 22032 54976
rect 22096 54912 22112 54976
rect 22176 54912 22192 54976
rect 22256 54912 22262 54976
rect 21946 54911 22262 54912
rect 26946 54976 27262 54977
rect 26946 54912 26952 54976
rect 27016 54912 27032 54976
rect 27096 54912 27112 54976
rect 27176 54912 27192 54976
rect 27256 54912 27262 54976
rect 26946 54911 27262 54912
rect 31946 54976 32262 54977
rect 31946 54912 31952 54976
rect 32016 54912 32032 54976
rect 32096 54912 32112 54976
rect 32176 54912 32192 54976
rect 32256 54912 32262 54976
rect 31946 54911 32262 54912
rect 36946 54976 37262 54977
rect 36946 54912 36952 54976
rect 37016 54912 37032 54976
rect 37096 54912 37112 54976
rect 37176 54912 37192 54976
rect 37256 54912 37262 54976
rect 36946 54911 37262 54912
rect 2606 54432 2922 54433
rect 2606 54368 2612 54432
rect 2676 54368 2692 54432
rect 2756 54368 2772 54432
rect 2836 54368 2852 54432
rect 2916 54368 2922 54432
rect 2606 54367 2922 54368
rect 7606 54432 7922 54433
rect 7606 54368 7612 54432
rect 7676 54368 7692 54432
rect 7756 54368 7772 54432
rect 7836 54368 7852 54432
rect 7916 54368 7922 54432
rect 7606 54367 7922 54368
rect 12606 54432 12922 54433
rect 12606 54368 12612 54432
rect 12676 54368 12692 54432
rect 12756 54368 12772 54432
rect 12836 54368 12852 54432
rect 12916 54368 12922 54432
rect 12606 54367 12922 54368
rect 17606 54432 17922 54433
rect 17606 54368 17612 54432
rect 17676 54368 17692 54432
rect 17756 54368 17772 54432
rect 17836 54368 17852 54432
rect 17916 54368 17922 54432
rect 17606 54367 17922 54368
rect 22606 54432 22922 54433
rect 22606 54368 22612 54432
rect 22676 54368 22692 54432
rect 22756 54368 22772 54432
rect 22836 54368 22852 54432
rect 22916 54368 22922 54432
rect 22606 54367 22922 54368
rect 27606 54432 27922 54433
rect 27606 54368 27612 54432
rect 27676 54368 27692 54432
rect 27756 54368 27772 54432
rect 27836 54368 27852 54432
rect 27916 54368 27922 54432
rect 27606 54367 27922 54368
rect 32606 54432 32922 54433
rect 32606 54368 32612 54432
rect 32676 54368 32692 54432
rect 32756 54368 32772 54432
rect 32836 54368 32852 54432
rect 32916 54368 32922 54432
rect 32606 54367 32922 54368
rect 37606 54432 37922 54433
rect 37606 54368 37612 54432
rect 37676 54368 37692 54432
rect 37756 54368 37772 54432
rect 37836 54368 37852 54432
rect 37916 54368 37922 54432
rect 37606 54367 37922 54368
rect 1946 53888 2262 53889
rect 1946 53824 1952 53888
rect 2016 53824 2032 53888
rect 2096 53824 2112 53888
rect 2176 53824 2192 53888
rect 2256 53824 2262 53888
rect 1946 53823 2262 53824
rect 6946 53888 7262 53889
rect 6946 53824 6952 53888
rect 7016 53824 7032 53888
rect 7096 53824 7112 53888
rect 7176 53824 7192 53888
rect 7256 53824 7262 53888
rect 6946 53823 7262 53824
rect 11946 53888 12262 53889
rect 11946 53824 11952 53888
rect 12016 53824 12032 53888
rect 12096 53824 12112 53888
rect 12176 53824 12192 53888
rect 12256 53824 12262 53888
rect 11946 53823 12262 53824
rect 16946 53888 17262 53889
rect 16946 53824 16952 53888
rect 17016 53824 17032 53888
rect 17096 53824 17112 53888
rect 17176 53824 17192 53888
rect 17256 53824 17262 53888
rect 16946 53823 17262 53824
rect 21946 53888 22262 53889
rect 21946 53824 21952 53888
rect 22016 53824 22032 53888
rect 22096 53824 22112 53888
rect 22176 53824 22192 53888
rect 22256 53824 22262 53888
rect 21946 53823 22262 53824
rect 26946 53888 27262 53889
rect 26946 53824 26952 53888
rect 27016 53824 27032 53888
rect 27096 53824 27112 53888
rect 27176 53824 27192 53888
rect 27256 53824 27262 53888
rect 26946 53823 27262 53824
rect 31946 53888 32262 53889
rect 31946 53824 31952 53888
rect 32016 53824 32032 53888
rect 32096 53824 32112 53888
rect 32176 53824 32192 53888
rect 32256 53824 32262 53888
rect 31946 53823 32262 53824
rect 36946 53888 37262 53889
rect 36946 53824 36952 53888
rect 37016 53824 37032 53888
rect 37096 53824 37112 53888
rect 37176 53824 37192 53888
rect 37256 53824 37262 53888
rect 36946 53823 37262 53824
rect 2606 53344 2922 53345
rect 2606 53280 2612 53344
rect 2676 53280 2692 53344
rect 2756 53280 2772 53344
rect 2836 53280 2852 53344
rect 2916 53280 2922 53344
rect 2606 53279 2922 53280
rect 7606 53344 7922 53345
rect 7606 53280 7612 53344
rect 7676 53280 7692 53344
rect 7756 53280 7772 53344
rect 7836 53280 7852 53344
rect 7916 53280 7922 53344
rect 7606 53279 7922 53280
rect 12606 53344 12922 53345
rect 12606 53280 12612 53344
rect 12676 53280 12692 53344
rect 12756 53280 12772 53344
rect 12836 53280 12852 53344
rect 12916 53280 12922 53344
rect 12606 53279 12922 53280
rect 17606 53344 17922 53345
rect 17606 53280 17612 53344
rect 17676 53280 17692 53344
rect 17756 53280 17772 53344
rect 17836 53280 17852 53344
rect 17916 53280 17922 53344
rect 17606 53279 17922 53280
rect 22606 53344 22922 53345
rect 22606 53280 22612 53344
rect 22676 53280 22692 53344
rect 22756 53280 22772 53344
rect 22836 53280 22852 53344
rect 22916 53280 22922 53344
rect 22606 53279 22922 53280
rect 27606 53344 27922 53345
rect 27606 53280 27612 53344
rect 27676 53280 27692 53344
rect 27756 53280 27772 53344
rect 27836 53280 27852 53344
rect 27916 53280 27922 53344
rect 27606 53279 27922 53280
rect 32606 53344 32922 53345
rect 32606 53280 32612 53344
rect 32676 53280 32692 53344
rect 32756 53280 32772 53344
rect 32836 53280 32852 53344
rect 32916 53280 32922 53344
rect 32606 53279 32922 53280
rect 37606 53344 37922 53345
rect 37606 53280 37612 53344
rect 37676 53280 37692 53344
rect 37756 53280 37772 53344
rect 37836 53280 37852 53344
rect 37916 53280 37922 53344
rect 37606 53279 37922 53280
rect 1946 52800 2262 52801
rect 1946 52736 1952 52800
rect 2016 52736 2032 52800
rect 2096 52736 2112 52800
rect 2176 52736 2192 52800
rect 2256 52736 2262 52800
rect 1946 52735 2262 52736
rect 6946 52800 7262 52801
rect 6946 52736 6952 52800
rect 7016 52736 7032 52800
rect 7096 52736 7112 52800
rect 7176 52736 7192 52800
rect 7256 52736 7262 52800
rect 6946 52735 7262 52736
rect 11946 52800 12262 52801
rect 11946 52736 11952 52800
rect 12016 52736 12032 52800
rect 12096 52736 12112 52800
rect 12176 52736 12192 52800
rect 12256 52736 12262 52800
rect 11946 52735 12262 52736
rect 16946 52800 17262 52801
rect 16946 52736 16952 52800
rect 17016 52736 17032 52800
rect 17096 52736 17112 52800
rect 17176 52736 17192 52800
rect 17256 52736 17262 52800
rect 16946 52735 17262 52736
rect 21946 52800 22262 52801
rect 21946 52736 21952 52800
rect 22016 52736 22032 52800
rect 22096 52736 22112 52800
rect 22176 52736 22192 52800
rect 22256 52736 22262 52800
rect 21946 52735 22262 52736
rect 26946 52800 27262 52801
rect 26946 52736 26952 52800
rect 27016 52736 27032 52800
rect 27096 52736 27112 52800
rect 27176 52736 27192 52800
rect 27256 52736 27262 52800
rect 26946 52735 27262 52736
rect 31946 52800 32262 52801
rect 31946 52736 31952 52800
rect 32016 52736 32032 52800
rect 32096 52736 32112 52800
rect 32176 52736 32192 52800
rect 32256 52736 32262 52800
rect 31946 52735 32262 52736
rect 36946 52800 37262 52801
rect 36946 52736 36952 52800
rect 37016 52736 37032 52800
rect 37096 52736 37112 52800
rect 37176 52736 37192 52800
rect 37256 52736 37262 52800
rect 36946 52735 37262 52736
rect 2606 52256 2922 52257
rect 2606 52192 2612 52256
rect 2676 52192 2692 52256
rect 2756 52192 2772 52256
rect 2836 52192 2852 52256
rect 2916 52192 2922 52256
rect 2606 52191 2922 52192
rect 7606 52256 7922 52257
rect 7606 52192 7612 52256
rect 7676 52192 7692 52256
rect 7756 52192 7772 52256
rect 7836 52192 7852 52256
rect 7916 52192 7922 52256
rect 7606 52191 7922 52192
rect 12606 52256 12922 52257
rect 12606 52192 12612 52256
rect 12676 52192 12692 52256
rect 12756 52192 12772 52256
rect 12836 52192 12852 52256
rect 12916 52192 12922 52256
rect 12606 52191 12922 52192
rect 17606 52256 17922 52257
rect 17606 52192 17612 52256
rect 17676 52192 17692 52256
rect 17756 52192 17772 52256
rect 17836 52192 17852 52256
rect 17916 52192 17922 52256
rect 17606 52191 17922 52192
rect 22606 52256 22922 52257
rect 22606 52192 22612 52256
rect 22676 52192 22692 52256
rect 22756 52192 22772 52256
rect 22836 52192 22852 52256
rect 22916 52192 22922 52256
rect 22606 52191 22922 52192
rect 27606 52256 27922 52257
rect 27606 52192 27612 52256
rect 27676 52192 27692 52256
rect 27756 52192 27772 52256
rect 27836 52192 27852 52256
rect 27916 52192 27922 52256
rect 27606 52191 27922 52192
rect 32606 52256 32922 52257
rect 32606 52192 32612 52256
rect 32676 52192 32692 52256
rect 32756 52192 32772 52256
rect 32836 52192 32852 52256
rect 32916 52192 32922 52256
rect 32606 52191 32922 52192
rect 37606 52256 37922 52257
rect 37606 52192 37612 52256
rect 37676 52192 37692 52256
rect 37756 52192 37772 52256
rect 37836 52192 37852 52256
rect 37916 52192 37922 52256
rect 37606 52191 37922 52192
rect 1946 51712 2262 51713
rect 1946 51648 1952 51712
rect 2016 51648 2032 51712
rect 2096 51648 2112 51712
rect 2176 51648 2192 51712
rect 2256 51648 2262 51712
rect 1946 51647 2262 51648
rect 6946 51712 7262 51713
rect 6946 51648 6952 51712
rect 7016 51648 7032 51712
rect 7096 51648 7112 51712
rect 7176 51648 7192 51712
rect 7256 51648 7262 51712
rect 6946 51647 7262 51648
rect 11946 51712 12262 51713
rect 11946 51648 11952 51712
rect 12016 51648 12032 51712
rect 12096 51648 12112 51712
rect 12176 51648 12192 51712
rect 12256 51648 12262 51712
rect 11946 51647 12262 51648
rect 16946 51712 17262 51713
rect 16946 51648 16952 51712
rect 17016 51648 17032 51712
rect 17096 51648 17112 51712
rect 17176 51648 17192 51712
rect 17256 51648 17262 51712
rect 16946 51647 17262 51648
rect 21946 51712 22262 51713
rect 21946 51648 21952 51712
rect 22016 51648 22032 51712
rect 22096 51648 22112 51712
rect 22176 51648 22192 51712
rect 22256 51648 22262 51712
rect 21946 51647 22262 51648
rect 26946 51712 27262 51713
rect 26946 51648 26952 51712
rect 27016 51648 27032 51712
rect 27096 51648 27112 51712
rect 27176 51648 27192 51712
rect 27256 51648 27262 51712
rect 26946 51647 27262 51648
rect 31946 51712 32262 51713
rect 31946 51648 31952 51712
rect 32016 51648 32032 51712
rect 32096 51648 32112 51712
rect 32176 51648 32192 51712
rect 32256 51648 32262 51712
rect 31946 51647 32262 51648
rect 36946 51712 37262 51713
rect 36946 51648 36952 51712
rect 37016 51648 37032 51712
rect 37096 51648 37112 51712
rect 37176 51648 37192 51712
rect 37256 51648 37262 51712
rect 36946 51647 37262 51648
rect 33133 51234 33199 51237
rect 33358 51234 33364 51236
rect 33133 51232 33364 51234
rect 33133 51176 33138 51232
rect 33194 51176 33364 51232
rect 33133 51174 33364 51176
rect 33133 51171 33199 51174
rect 33358 51172 33364 51174
rect 33428 51172 33434 51236
rect 2606 51168 2922 51169
rect 2606 51104 2612 51168
rect 2676 51104 2692 51168
rect 2756 51104 2772 51168
rect 2836 51104 2852 51168
rect 2916 51104 2922 51168
rect 2606 51103 2922 51104
rect 7606 51168 7922 51169
rect 7606 51104 7612 51168
rect 7676 51104 7692 51168
rect 7756 51104 7772 51168
rect 7836 51104 7852 51168
rect 7916 51104 7922 51168
rect 7606 51103 7922 51104
rect 12606 51168 12922 51169
rect 12606 51104 12612 51168
rect 12676 51104 12692 51168
rect 12756 51104 12772 51168
rect 12836 51104 12852 51168
rect 12916 51104 12922 51168
rect 12606 51103 12922 51104
rect 17606 51168 17922 51169
rect 17606 51104 17612 51168
rect 17676 51104 17692 51168
rect 17756 51104 17772 51168
rect 17836 51104 17852 51168
rect 17916 51104 17922 51168
rect 17606 51103 17922 51104
rect 22606 51168 22922 51169
rect 22606 51104 22612 51168
rect 22676 51104 22692 51168
rect 22756 51104 22772 51168
rect 22836 51104 22852 51168
rect 22916 51104 22922 51168
rect 22606 51103 22922 51104
rect 27606 51168 27922 51169
rect 27606 51104 27612 51168
rect 27676 51104 27692 51168
rect 27756 51104 27772 51168
rect 27836 51104 27852 51168
rect 27916 51104 27922 51168
rect 27606 51103 27922 51104
rect 32606 51168 32922 51169
rect 32606 51104 32612 51168
rect 32676 51104 32692 51168
rect 32756 51104 32772 51168
rect 32836 51104 32852 51168
rect 32916 51104 32922 51168
rect 32606 51103 32922 51104
rect 37606 51168 37922 51169
rect 37606 51104 37612 51168
rect 37676 51104 37692 51168
rect 37756 51104 37772 51168
rect 37836 51104 37852 51168
rect 37916 51104 37922 51168
rect 37606 51103 37922 51104
rect 31702 50900 31708 50964
rect 31772 50962 31778 50964
rect 32438 50962 32444 50964
rect 31772 50902 32444 50962
rect 31772 50900 31778 50902
rect 32438 50900 32444 50902
rect 32508 50900 32514 50964
rect 1946 50624 2262 50625
rect 1946 50560 1952 50624
rect 2016 50560 2032 50624
rect 2096 50560 2112 50624
rect 2176 50560 2192 50624
rect 2256 50560 2262 50624
rect 1946 50559 2262 50560
rect 6946 50624 7262 50625
rect 6946 50560 6952 50624
rect 7016 50560 7032 50624
rect 7096 50560 7112 50624
rect 7176 50560 7192 50624
rect 7256 50560 7262 50624
rect 6946 50559 7262 50560
rect 11946 50624 12262 50625
rect 11946 50560 11952 50624
rect 12016 50560 12032 50624
rect 12096 50560 12112 50624
rect 12176 50560 12192 50624
rect 12256 50560 12262 50624
rect 11946 50559 12262 50560
rect 16946 50624 17262 50625
rect 16946 50560 16952 50624
rect 17016 50560 17032 50624
rect 17096 50560 17112 50624
rect 17176 50560 17192 50624
rect 17256 50560 17262 50624
rect 16946 50559 17262 50560
rect 21946 50624 22262 50625
rect 21946 50560 21952 50624
rect 22016 50560 22032 50624
rect 22096 50560 22112 50624
rect 22176 50560 22192 50624
rect 22256 50560 22262 50624
rect 21946 50559 22262 50560
rect 26946 50624 27262 50625
rect 26946 50560 26952 50624
rect 27016 50560 27032 50624
rect 27096 50560 27112 50624
rect 27176 50560 27192 50624
rect 27256 50560 27262 50624
rect 26946 50559 27262 50560
rect 31946 50624 32262 50625
rect 31946 50560 31952 50624
rect 32016 50560 32032 50624
rect 32096 50560 32112 50624
rect 32176 50560 32192 50624
rect 32256 50560 32262 50624
rect 31946 50559 32262 50560
rect 36946 50624 37262 50625
rect 36946 50560 36952 50624
rect 37016 50560 37032 50624
rect 37096 50560 37112 50624
rect 37176 50560 37192 50624
rect 37256 50560 37262 50624
rect 36946 50559 37262 50560
rect 2606 50080 2922 50081
rect 2606 50016 2612 50080
rect 2676 50016 2692 50080
rect 2756 50016 2772 50080
rect 2836 50016 2852 50080
rect 2916 50016 2922 50080
rect 2606 50015 2922 50016
rect 7606 50080 7922 50081
rect 7606 50016 7612 50080
rect 7676 50016 7692 50080
rect 7756 50016 7772 50080
rect 7836 50016 7852 50080
rect 7916 50016 7922 50080
rect 7606 50015 7922 50016
rect 12606 50080 12922 50081
rect 12606 50016 12612 50080
rect 12676 50016 12692 50080
rect 12756 50016 12772 50080
rect 12836 50016 12852 50080
rect 12916 50016 12922 50080
rect 12606 50015 12922 50016
rect 17606 50080 17922 50081
rect 17606 50016 17612 50080
rect 17676 50016 17692 50080
rect 17756 50016 17772 50080
rect 17836 50016 17852 50080
rect 17916 50016 17922 50080
rect 17606 50015 17922 50016
rect 22606 50080 22922 50081
rect 22606 50016 22612 50080
rect 22676 50016 22692 50080
rect 22756 50016 22772 50080
rect 22836 50016 22852 50080
rect 22916 50016 22922 50080
rect 22606 50015 22922 50016
rect 27606 50080 27922 50081
rect 27606 50016 27612 50080
rect 27676 50016 27692 50080
rect 27756 50016 27772 50080
rect 27836 50016 27852 50080
rect 27916 50016 27922 50080
rect 27606 50015 27922 50016
rect 32606 50080 32922 50081
rect 32606 50016 32612 50080
rect 32676 50016 32692 50080
rect 32756 50016 32772 50080
rect 32836 50016 32852 50080
rect 32916 50016 32922 50080
rect 32606 50015 32922 50016
rect 37606 50080 37922 50081
rect 37606 50016 37612 50080
rect 37676 50016 37692 50080
rect 37756 50016 37772 50080
rect 37836 50016 37852 50080
rect 37916 50016 37922 50080
rect 37606 50015 37922 50016
rect 1946 49536 2262 49537
rect 1946 49472 1952 49536
rect 2016 49472 2032 49536
rect 2096 49472 2112 49536
rect 2176 49472 2192 49536
rect 2256 49472 2262 49536
rect 1946 49471 2262 49472
rect 6946 49536 7262 49537
rect 6946 49472 6952 49536
rect 7016 49472 7032 49536
rect 7096 49472 7112 49536
rect 7176 49472 7192 49536
rect 7256 49472 7262 49536
rect 6946 49471 7262 49472
rect 11946 49536 12262 49537
rect 11946 49472 11952 49536
rect 12016 49472 12032 49536
rect 12096 49472 12112 49536
rect 12176 49472 12192 49536
rect 12256 49472 12262 49536
rect 11946 49471 12262 49472
rect 16946 49536 17262 49537
rect 16946 49472 16952 49536
rect 17016 49472 17032 49536
rect 17096 49472 17112 49536
rect 17176 49472 17192 49536
rect 17256 49472 17262 49536
rect 16946 49471 17262 49472
rect 21946 49536 22262 49537
rect 21946 49472 21952 49536
rect 22016 49472 22032 49536
rect 22096 49472 22112 49536
rect 22176 49472 22192 49536
rect 22256 49472 22262 49536
rect 21946 49471 22262 49472
rect 26946 49536 27262 49537
rect 26946 49472 26952 49536
rect 27016 49472 27032 49536
rect 27096 49472 27112 49536
rect 27176 49472 27192 49536
rect 27256 49472 27262 49536
rect 26946 49471 27262 49472
rect 31946 49536 32262 49537
rect 31946 49472 31952 49536
rect 32016 49472 32032 49536
rect 32096 49472 32112 49536
rect 32176 49472 32192 49536
rect 32256 49472 32262 49536
rect 31946 49471 32262 49472
rect 36946 49536 37262 49537
rect 36946 49472 36952 49536
rect 37016 49472 37032 49536
rect 37096 49472 37112 49536
rect 37176 49472 37192 49536
rect 37256 49472 37262 49536
rect 36946 49471 37262 49472
rect 2606 48992 2922 48993
rect 2606 48928 2612 48992
rect 2676 48928 2692 48992
rect 2756 48928 2772 48992
rect 2836 48928 2852 48992
rect 2916 48928 2922 48992
rect 2606 48927 2922 48928
rect 7606 48992 7922 48993
rect 7606 48928 7612 48992
rect 7676 48928 7692 48992
rect 7756 48928 7772 48992
rect 7836 48928 7852 48992
rect 7916 48928 7922 48992
rect 7606 48927 7922 48928
rect 12606 48992 12922 48993
rect 12606 48928 12612 48992
rect 12676 48928 12692 48992
rect 12756 48928 12772 48992
rect 12836 48928 12852 48992
rect 12916 48928 12922 48992
rect 12606 48927 12922 48928
rect 17606 48992 17922 48993
rect 17606 48928 17612 48992
rect 17676 48928 17692 48992
rect 17756 48928 17772 48992
rect 17836 48928 17852 48992
rect 17916 48928 17922 48992
rect 17606 48927 17922 48928
rect 22606 48992 22922 48993
rect 22606 48928 22612 48992
rect 22676 48928 22692 48992
rect 22756 48928 22772 48992
rect 22836 48928 22852 48992
rect 22916 48928 22922 48992
rect 22606 48927 22922 48928
rect 27606 48992 27922 48993
rect 27606 48928 27612 48992
rect 27676 48928 27692 48992
rect 27756 48928 27772 48992
rect 27836 48928 27852 48992
rect 27916 48928 27922 48992
rect 27606 48927 27922 48928
rect 32606 48992 32922 48993
rect 32606 48928 32612 48992
rect 32676 48928 32692 48992
rect 32756 48928 32772 48992
rect 32836 48928 32852 48992
rect 32916 48928 32922 48992
rect 32606 48927 32922 48928
rect 37606 48992 37922 48993
rect 37606 48928 37612 48992
rect 37676 48928 37692 48992
rect 37756 48928 37772 48992
rect 37836 48928 37852 48992
rect 37916 48928 37922 48992
rect 37606 48927 37922 48928
rect 1946 48448 2262 48449
rect 1946 48384 1952 48448
rect 2016 48384 2032 48448
rect 2096 48384 2112 48448
rect 2176 48384 2192 48448
rect 2256 48384 2262 48448
rect 1946 48383 2262 48384
rect 6946 48448 7262 48449
rect 6946 48384 6952 48448
rect 7016 48384 7032 48448
rect 7096 48384 7112 48448
rect 7176 48384 7192 48448
rect 7256 48384 7262 48448
rect 6946 48383 7262 48384
rect 11946 48448 12262 48449
rect 11946 48384 11952 48448
rect 12016 48384 12032 48448
rect 12096 48384 12112 48448
rect 12176 48384 12192 48448
rect 12256 48384 12262 48448
rect 11946 48383 12262 48384
rect 16946 48448 17262 48449
rect 16946 48384 16952 48448
rect 17016 48384 17032 48448
rect 17096 48384 17112 48448
rect 17176 48384 17192 48448
rect 17256 48384 17262 48448
rect 16946 48383 17262 48384
rect 21946 48448 22262 48449
rect 21946 48384 21952 48448
rect 22016 48384 22032 48448
rect 22096 48384 22112 48448
rect 22176 48384 22192 48448
rect 22256 48384 22262 48448
rect 21946 48383 22262 48384
rect 26946 48448 27262 48449
rect 26946 48384 26952 48448
rect 27016 48384 27032 48448
rect 27096 48384 27112 48448
rect 27176 48384 27192 48448
rect 27256 48384 27262 48448
rect 26946 48383 27262 48384
rect 31946 48448 32262 48449
rect 31946 48384 31952 48448
rect 32016 48384 32032 48448
rect 32096 48384 32112 48448
rect 32176 48384 32192 48448
rect 32256 48384 32262 48448
rect 31946 48383 32262 48384
rect 36946 48448 37262 48449
rect 36946 48384 36952 48448
rect 37016 48384 37032 48448
rect 37096 48384 37112 48448
rect 37176 48384 37192 48448
rect 37256 48384 37262 48448
rect 36946 48383 37262 48384
rect 2606 47904 2922 47905
rect 2606 47840 2612 47904
rect 2676 47840 2692 47904
rect 2756 47840 2772 47904
rect 2836 47840 2852 47904
rect 2916 47840 2922 47904
rect 2606 47839 2922 47840
rect 7606 47904 7922 47905
rect 7606 47840 7612 47904
rect 7676 47840 7692 47904
rect 7756 47840 7772 47904
rect 7836 47840 7852 47904
rect 7916 47840 7922 47904
rect 7606 47839 7922 47840
rect 12606 47904 12922 47905
rect 12606 47840 12612 47904
rect 12676 47840 12692 47904
rect 12756 47840 12772 47904
rect 12836 47840 12852 47904
rect 12916 47840 12922 47904
rect 12606 47839 12922 47840
rect 17606 47904 17922 47905
rect 17606 47840 17612 47904
rect 17676 47840 17692 47904
rect 17756 47840 17772 47904
rect 17836 47840 17852 47904
rect 17916 47840 17922 47904
rect 17606 47839 17922 47840
rect 22606 47904 22922 47905
rect 22606 47840 22612 47904
rect 22676 47840 22692 47904
rect 22756 47840 22772 47904
rect 22836 47840 22852 47904
rect 22916 47840 22922 47904
rect 22606 47839 22922 47840
rect 27606 47904 27922 47905
rect 27606 47840 27612 47904
rect 27676 47840 27692 47904
rect 27756 47840 27772 47904
rect 27836 47840 27852 47904
rect 27916 47840 27922 47904
rect 27606 47839 27922 47840
rect 32606 47904 32922 47905
rect 32606 47840 32612 47904
rect 32676 47840 32692 47904
rect 32756 47840 32772 47904
rect 32836 47840 32852 47904
rect 32916 47840 32922 47904
rect 32606 47839 32922 47840
rect 37606 47904 37922 47905
rect 37606 47840 37612 47904
rect 37676 47840 37692 47904
rect 37756 47840 37772 47904
rect 37836 47840 37852 47904
rect 37916 47840 37922 47904
rect 37606 47839 37922 47840
rect 1946 47360 2262 47361
rect 1946 47296 1952 47360
rect 2016 47296 2032 47360
rect 2096 47296 2112 47360
rect 2176 47296 2192 47360
rect 2256 47296 2262 47360
rect 1946 47295 2262 47296
rect 6946 47360 7262 47361
rect 6946 47296 6952 47360
rect 7016 47296 7032 47360
rect 7096 47296 7112 47360
rect 7176 47296 7192 47360
rect 7256 47296 7262 47360
rect 6946 47295 7262 47296
rect 11946 47360 12262 47361
rect 11946 47296 11952 47360
rect 12016 47296 12032 47360
rect 12096 47296 12112 47360
rect 12176 47296 12192 47360
rect 12256 47296 12262 47360
rect 11946 47295 12262 47296
rect 16946 47360 17262 47361
rect 16946 47296 16952 47360
rect 17016 47296 17032 47360
rect 17096 47296 17112 47360
rect 17176 47296 17192 47360
rect 17256 47296 17262 47360
rect 16946 47295 17262 47296
rect 21946 47360 22262 47361
rect 21946 47296 21952 47360
rect 22016 47296 22032 47360
rect 22096 47296 22112 47360
rect 22176 47296 22192 47360
rect 22256 47296 22262 47360
rect 21946 47295 22262 47296
rect 26946 47360 27262 47361
rect 26946 47296 26952 47360
rect 27016 47296 27032 47360
rect 27096 47296 27112 47360
rect 27176 47296 27192 47360
rect 27256 47296 27262 47360
rect 26946 47295 27262 47296
rect 31946 47360 32262 47361
rect 31946 47296 31952 47360
rect 32016 47296 32032 47360
rect 32096 47296 32112 47360
rect 32176 47296 32192 47360
rect 32256 47296 32262 47360
rect 31946 47295 32262 47296
rect 36946 47360 37262 47361
rect 36946 47296 36952 47360
rect 37016 47296 37032 47360
rect 37096 47296 37112 47360
rect 37176 47296 37192 47360
rect 37256 47296 37262 47360
rect 36946 47295 37262 47296
rect 2606 46816 2922 46817
rect 2606 46752 2612 46816
rect 2676 46752 2692 46816
rect 2756 46752 2772 46816
rect 2836 46752 2852 46816
rect 2916 46752 2922 46816
rect 2606 46751 2922 46752
rect 7606 46816 7922 46817
rect 7606 46752 7612 46816
rect 7676 46752 7692 46816
rect 7756 46752 7772 46816
rect 7836 46752 7852 46816
rect 7916 46752 7922 46816
rect 7606 46751 7922 46752
rect 12606 46816 12922 46817
rect 12606 46752 12612 46816
rect 12676 46752 12692 46816
rect 12756 46752 12772 46816
rect 12836 46752 12852 46816
rect 12916 46752 12922 46816
rect 12606 46751 12922 46752
rect 17606 46816 17922 46817
rect 17606 46752 17612 46816
rect 17676 46752 17692 46816
rect 17756 46752 17772 46816
rect 17836 46752 17852 46816
rect 17916 46752 17922 46816
rect 17606 46751 17922 46752
rect 22606 46816 22922 46817
rect 22606 46752 22612 46816
rect 22676 46752 22692 46816
rect 22756 46752 22772 46816
rect 22836 46752 22852 46816
rect 22916 46752 22922 46816
rect 22606 46751 22922 46752
rect 27606 46816 27922 46817
rect 27606 46752 27612 46816
rect 27676 46752 27692 46816
rect 27756 46752 27772 46816
rect 27836 46752 27852 46816
rect 27916 46752 27922 46816
rect 27606 46751 27922 46752
rect 32606 46816 32922 46817
rect 32606 46752 32612 46816
rect 32676 46752 32692 46816
rect 32756 46752 32772 46816
rect 32836 46752 32852 46816
rect 32916 46752 32922 46816
rect 32606 46751 32922 46752
rect 37606 46816 37922 46817
rect 37606 46752 37612 46816
rect 37676 46752 37692 46816
rect 37756 46752 37772 46816
rect 37836 46752 37852 46816
rect 37916 46752 37922 46816
rect 37606 46751 37922 46752
rect 1946 46272 2262 46273
rect 1946 46208 1952 46272
rect 2016 46208 2032 46272
rect 2096 46208 2112 46272
rect 2176 46208 2192 46272
rect 2256 46208 2262 46272
rect 1946 46207 2262 46208
rect 6946 46272 7262 46273
rect 6946 46208 6952 46272
rect 7016 46208 7032 46272
rect 7096 46208 7112 46272
rect 7176 46208 7192 46272
rect 7256 46208 7262 46272
rect 6946 46207 7262 46208
rect 11946 46272 12262 46273
rect 11946 46208 11952 46272
rect 12016 46208 12032 46272
rect 12096 46208 12112 46272
rect 12176 46208 12192 46272
rect 12256 46208 12262 46272
rect 11946 46207 12262 46208
rect 16946 46272 17262 46273
rect 16946 46208 16952 46272
rect 17016 46208 17032 46272
rect 17096 46208 17112 46272
rect 17176 46208 17192 46272
rect 17256 46208 17262 46272
rect 16946 46207 17262 46208
rect 21946 46272 22262 46273
rect 21946 46208 21952 46272
rect 22016 46208 22032 46272
rect 22096 46208 22112 46272
rect 22176 46208 22192 46272
rect 22256 46208 22262 46272
rect 21946 46207 22262 46208
rect 26946 46272 27262 46273
rect 26946 46208 26952 46272
rect 27016 46208 27032 46272
rect 27096 46208 27112 46272
rect 27176 46208 27192 46272
rect 27256 46208 27262 46272
rect 26946 46207 27262 46208
rect 31946 46272 32262 46273
rect 31946 46208 31952 46272
rect 32016 46208 32032 46272
rect 32096 46208 32112 46272
rect 32176 46208 32192 46272
rect 32256 46208 32262 46272
rect 31946 46207 32262 46208
rect 36946 46272 37262 46273
rect 36946 46208 36952 46272
rect 37016 46208 37032 46272
rect 37096 46208 37112 46272
rect 37176 46208 37192 46272
rect 37256 46208 37262 46272
rect 36946 46207 37262 46208
rect 14549 45930 14615 45933
rect 21030 45930 21036 45932
rect 14549 45928 21036 45930
rect 14549 45872 14554 45928
rect 14610 45872 21036 45928
rect 14549 45870 21036 45872
rect 14549 45867 14615 45870
rect 21030 45868 21036 45870
rect 21100 45930 21106 45932
rect 28809 45930 28875 45933
rect 21100 45928 28875 45930
rect 21100 45872 28814 45928
rect 28870 45872 28875 45928
rect 21100 45870 28875 45872
rect 21100 45868 21106 45870
rect 28809 45867 28875 45870
rect 2606 45728 2922 45729
rect 2606 45664 2612 45728
rect 2676 45664 2692 45728
rect 2756 45664 2772 45728
rect 2836 45664 2852 45728
rect 2916 45664 2922 45728
rect 2606 45663 2922 45664
rect 7606 45728 7922 45729
rect 7606 45664 7612 45728
rect 7676 45664 7692 45728
rect 7756 45664 7772 45728
rect 7836 45664 7852 45728
rect 7916 45664 7922 45728
rect 7606 45663 7922 45664
rect 12606 45728 12922 45729
rect 12606 45664 12612 45728
rect 12676 45664 12692 45728
rect 12756 45664 12772 45728
rect 12836 45664 12852 45728
rect 12916 45664 12922 45728
rect 12606 45663 12922 45664
rect 17606 45728 17922 45729
rect 17606 45664 17612 45728
rect 17676 45664 17692 45728
rect 17756 45664 17772 45728
rect 17836 45664 17852 45728
rect 17916 45664 17922 45728
rect 17606 45663 17922 45664
rect 22606 45728 22922 45729
rect 22606 45664 22612 45728
rect 22676 45664 22692 45728
rect 22756 45664 22772 45728
rect 22836 45664 22852 45728
rect 22916 45664 22922 45728
rect 22606 45663 22922 45664
rect 27606 45728 27922 45729
rect 27606 45664 27612 45728
rect 27676 45664 27692 45728
rect 27756 45664 27772 45728
rect 27836 45664 27852 45728
rect 27916 45664 27922 45728
rect 27606 45663 27922 45664
rect 32606 45728 32922 45729
rect 32606 45664 32612 45728
rect 32676 45664 32692 45728
rect 32756 45664 32772 45728
rect 32836 45664 32852 45728
rect 32916 45664 32922 45728
rect 32606 45663 32922 45664
rect 37606 45728 37922 45729
rect 37606 45664 37612 45728
rect 37676 45664 37692 45728
rect 37756 45664 37772 45728
rect 37836 45664 37852 45728
rect 37916 45664 37922 45728
rect 37606 45663 37922 45664
rect 1946 45184 2262 45185
rect 1946 45120 1952 45184
rect 2016 45120 2032 45184
rect 2096 45120 2112 45184
rect 2176 45120 2192 45184
rect 2256 45120 2262 45184
rect 1946 45119 2262 45120
rect 6946 45184 7262 45185
rect 6946 45120 6952 45184
rect 7016 45120 7032 45184
rect 7096 45120 7112 45184
rect 7176 45120 7192 45184
rect 7256 45120 7262 45184
rect 6946 45119 7262 45120
rect 11946 45184 12262 45185
rect 11946 45120 11952 45184
rect 12016 45120 12032 45184
rect 12096 45120 12112 45184
rect 12176 45120 12192 45184
rect 12256 45120 12262 45184
rect 11946 45119 12262 45120
rect 16946 45184 17262 45185
rect 16946 45120 16952 45184
rect 17016 45120 17032 45184
rect 17096 45120 17112 45184
rect 17176 45120 17192 45184
rect 17256 45120 17262 45184
rect 16946 45119 17262 45120
rect 21946 45184 22262 45185
rect 21946 45120 21952 45184
rect 22016 45120 22032 45184
rect 22096 45120 22112 45184
rect 22176 45120 22192 45184
rect 22256 45120 22262 45184
rect 21946 45119 22262 45120
rect 26946 45184 27262 45185
rect 26946 45120 26952 45184
rect 27016 45120 27032 45184
rect 27096 45120 27112 45184
rect 27176 45120 27192 45184
rect 27256 45120 27262 45184
rect 26946 45119 27262 45120
rect 31946 45184 32262 45185
rect 31946 45120 31952 45184
rect 32016 45120 32032 45184
rect 32096 45120 32112 45184
rect 32176 45120 32192 45184
rect 32256 45120 32262 45184
rect 31946 45119 32262 45120
rect 36946 45184 37262 45185
rect 36946 45120 36952 45184
rect 37016 45120 37032 45184
rect 37096 45120 37112 45184
rect 37176 45120 37192 45184
rect 37256 45120 37262 45184
rect 36946 45119 37262 45120
rect 2606 44640 2922 44641
rect 2606 44576 2612 44640
rect 2676 44576 2692 44640
rect 2756 44576 2772 44640
rect 2836 44576 2852 44640
rect 2916 44576 2922 44640
rect 2606 44575 2922 44576
rect 7606 44640 7922 44641
rect 7606 44576 7612 44640
rect 7676 44576 7692 44640
rect 7756 44576 7772 44640
rect 7836 44576 7852 44640
rect 7916 44576 7922 44640
rect 7606 44575 7922 44576
rect 12606 44640 12922 44641
rect 12606 44576 12612 44640
rect 12676 44576 12692 44640
rect 12756 44576 12772 44640
rect 12836 44576 12852 44640
rect 12916 44576 12922 44640
rect 12606 44575 12922 44576
rect 17606 44640 17922 44641
rect 17606 44576 17612 44640
rect 17676 44576 17692 44640
rect 17756 44576 17772 44640
rect 17836 44576 17852 44640
rect 17916 44576 17922 44640
rect 17606 44575 17922 44576
rect 22606 44640 22922 44641
rect 22606 44576 22612 44640
rect 22676 44576 22692 44640
rect 22756 44576 22772 44640
rect 22836 44576 22852 44640
rect 22916 44576 22922 44640
rect 22606 44575 22922 44576
rect 27606 44640 27922 44641
rect 27606 44576 27612 44640
rect 27676 44576 27692 44640
rect 27756 44576 27772 44640
rect 27836 44576 27852 44640
rect 27916 44576 27922 44640
rect 27606 44575 27922 44576
rect 32606 44640 32922 44641
rect 32606 44576 32612 44640
rect 32676 44576 32692 44640
rect 32756 44576 32772 44640
rect 32836 44576 32852 44640
rect 32916 44576 32922 44640
rect 32606 44575 32922 44576
rect 37606 44640 37922 44641
rect 37606 44576 37612 44640
rect 37676 44576 37692 44640
rect 37756 44576 37772 44640
rect 37836 44576 37852 44640
rect 37916 44576 37922 44640
rect 37606 44575 37922 44576
rect 1946 44096 2262 44097
rect 1946 44032 1952 44096
rect 2016 44032 2032 44096
rect 2096 44032 2112 44096
rect 2176 44032 2192 44096
rect 2256 44032 2262 44096
rect 1946 44031 2262 44032
rect 6946 44096 7262 44097
rect 6946 44032 6952 44096
rect 7016 44032 7032 44096
rect 7096 44032 7112 44096
rect 7176 44032 7192 44096
rect 7256 44032 7262 44096
rect 6946 44031 7262 44032
rect 11946 44096 12262 44097
rect 11946 44032 11952 44096
rect 12016 44032 12032 44096
rect 12096 44032 12112 44096
rect 12176 44032 12192 44096
rect 12256 44032 12262 44096
rect 11946 44031 12262 44032
rect 16946 44096 17262 44097
rect 16946 44032 16952 44096
rect 17016 44032 17032 44096
rect 17096 44032 17112 44096
rect 17176 44032 17192 44096
rect 17256 44032 17262 44096
rect 16946 44031 17262 44032
rect 21946 44096 22262 44097
rect 21946 44032 21952 44096
rect 22016 44032 22032 44096
rect 22096 44032 22112 44096
rect 22176 44032 22192 44096
rect 22256 44032 22262 44096
rect 21946 44031 22262 44032
rect 26946 44096 27262 44097
rect 26946 44032 26952 44096
rect 27016 44032 27032 44096
rect 27096 44032 27112 44096
rect 27176 44032 27192 44096
rect 27256 44032 27262 44096
rect 26946 44031 27262 44032
rect 31946 44096 32262 44097
rect 31946 44032 31952 44096
rect 32016 44032 32032 44096
rect 32096 44032 32112 44096
rect 32176 44032 32192 44096
rect 32256 44032 32262 44096
rect 31946 44031 32262 44032
rect 36946 44096 37262 44097
rect 36946 44032 36952 44096
rect 37016 44032 37032 44096
rect 37096 44032 37112 44096
rect 37176 44032 37192 44096
rect 37256 44032 37262 44096
rect 36946 44031 37262 44032
rect 2606 43552 2922 43553
rect 2606 43488 2612 43552
rect 2676 43488 2692 43552
rect 2756 43488 2772 43552
rect 2836 43488 2852 43552
rect 2916 43488 2922 43552
rect 2606 43487 2922 43488
rect 7606 43552 7922 43553
rect 7606 43488 7612 43552
rect 7676 43488 7692 43552
rect 7756 43488 7772 43552
rect 7836 43488 7852 43552
rect 7916 43488 7922 43552
rect 7606 43487 7922 43488
rect 12606 43552 12922 43553
rect 12606 43488 12612 43552
rect 12676 43488 12692 43552
rect 12756 43488 12772 43552
rect 12836 43488 12852 43552
rect 12916 43488 12922 43552
rect 12606 43487 12922 43488
rect 17606 43552 17922 43553
rect 17606 43488 17612 43552
rect 17676 43488 17692 43552
rect 17756 43488 17772 43552
rect 17836 43488 17852 43552
rect 17916 43488 17922 43552
rect 17606 43487 17922 43488
rect 22606 43552 22922 43553
rect 22606 43488 22612 43552
rect 22676 43488 22692 43552
rect 22756 43488 22772 43552
rect 22836 43488 22852 43552
rect 22916 43488 22922 43552
rect 22606 43487 22922 43488
rect 27606 43552 27922 43553
rect 27606 43488 27612 43552
rect 27676 43488 27692 43552
rect 27756 43488 27772 43552
rect 27836 43488 27852 43552
rect 27916 43488 27922 43552
rect 27606 43487 27922 43488
rect 32606 43552 32922 43553
rect 32606 43488 32612 43552
rect 32676 43488 32692 43552
rect 32756 43488 32772 43552
rect 32836 43488 32852 43552
rect 32916 43488 32922 43552
rect 32606 43487 32922 43488
rect 37606 43552 37922 43553
rect 37606 43488 37612 43552
rect 37676 43488 37692 43552
rect 37756 43488 37772 43552
rect 37836 43488 37852 43552
rect 37916 43488 37922 43552
rect 37606 43487 37922 43488
rect 1946 43008 2262 43009
rect 1946 42944 1952 43008
rect 2016 42944 2032 43008
rect 2096 42944 2112 43008
rect 2176 42944 2192 43008
rect 2256 42944 2262 43008
rect 1946 42943 2262 42944
rect 6946 43008 7262 43009
rect 6946 42944 6952 43008
rect 7016 42944 7032 43008
rect 7096 42944 7112 43008
rect 7176 42944 7192 43008
rect 7256 42944 7262 43008
rect 6946 42943 7262 42944
rect 11946 43008 12262 43009
rect 11946 42944 11952 43008
rect 12016 42944 12032 43008
rect 12096 42944 12112 43008
rect 12176 42944 12192 43008
rect 12256 42944 12262 43008
rect 11946 42943 12262 42944
rect 16946 43008 17262 43009
rect 16946 42944 16952 43008
rect 17016 42944 17032 43008
rect 17096 42944 17112 43008
rect 17176 42944 17192 43008
rect 17256 42944 17262 43008
rect 16946 42943 17262 42944
rect 21946 43008 22262 43009
rect 21946 42944 21952 43008
rect 22016 42944 22032 43008
rect 22096 42944 22112 43008
rect 22176 42944 22192 43008
rect 22256 42944 22262 43008
rect 21946 42943 22262 42944
rect 26946 43008 27262 43009
rect 26946 42944 26952 43008
rect 27016 42944 27032 43008
rect 27096 42944 27112 43008
rect 27176 42944 27192 43008
rect 27256 42944 27262 43008
rect 26946 42943 27262 42944
rect 31946 43008 32262 43009
rect 31946 42944 31952 43008
rect 32016 42944 32032 43008
rect 32096 42944 32112 43008
rect 32176 42944 32192 43008
rect 32256 42944 32262 43008
rect 31946 42943 32262 42944
rect 36946 43008 37262 43009
rect 36946 42944 36952 43008
rect 37016 42944 37032 43008
rect 37096 42944 37112 43008
rect 37176 42944 37192 43008
rect 37256 42944 37262 43008
rect 36946 42943 37262 42944
rect 2606 42464 2922 42465
rect 2606 42400 2612 42464
rect 2676 42400 2692 42464
rect 2756 42400 2772 42464
rect 2836 42400 2852 42464
rect 2916 42400 2922 42464
rect 2606 42399 2922 42400
rect 7606 42464 7922 42465
rect 7606 42400 7612 42464
rect 7676 42400 7692 42464
rect 7756 42400 7772 42464
rect 7836 42400 7852 42464
rect 7916 42400 7922 42464
rect 7606 42399 7922 42400
rect 12606 42464 12922 42465
rect 12606 42400 12612 42464
rect 12676 42400 12692 42464
rect 12756 42400 12772 42464
rect 12836 42400 12852 42464
rect 12916 42400 12922 42464
rect 12606 42399 12922 42400
rect 17606 42464 17922 42465
rect 17606 42400 17612 42464
rect 17676 42400 17692 42464
rect 17756 42400 17772 42464
rect 17836 42400 17852 42464
rect 17916 42400 17922 42464
rect 17606 42399 17922 42400
rect 22606 42464 22922 42465
rect 22606 42400 22612 42464
rect 22676 42400 22692 42464
rect 22756 42400 22772 42464
rect 22836 42400 22852 42464
rect 22916 42400 22922 42464
rect 22606 42399 22922 42400
rect 27606 42464 27922 42465
rect 27606 42400 27612 42464
rect 27676 42400 27692 42464
rect 27756 42400 27772 42464
rect 27836 42400 27852 42464
rect 27916 42400 27922 42464
rect 27606 42399 27922 42400
rect 32606 42464 32922 42465
rect 32606 42400 32612 42464
rect 32676 42400 32692 42464
rect 32756 42400 32772 42464
rect 32836 42400 32852 42464
rect 32916 42400 32922 42464
rect 32606 42399 32922 42400
rect 37606 42464 37922 42465
rect 37606 42400 37612 42464
rect 37676 42400 37692 42464
rect 37756 42400 37772 42464
rect 37836 42400 37852 42464
rect 37916 42400 37922 42464
rect 37606 42399 37922 42400
rect 1946 41920 2262 41921
rect 1946 41856 1952 41920
rect 2016 41856 2032 41920
rect 2096 41856 2112 41920
rect 2176 41856 2192 41920
rect 2256 41856 2262 41920
rect 1946 41855 2262 41856
rect 6946 41920 7262 41921
rect 6946 41856 6952 41920
rect 7016 41856 7032 41920
rect 7096 41856 7112 41920
rect 7176 41856 7192 41920
rect 7256 41856 7262 41920
rect 6946 41855 7262 41856
rect 11946 41920 12262 41921
rect 11946 41856 11952 41920
rect 12016 41856 12032 41920
rect 12096 41856 12112 41920
rect 12176 41856 12192 41920
rect 12256 41856 12262 41920
rect 11946 41855 12262 41856
rect 16946 41920 17262 41921
rect 16946 41856 16952 41920
rect 17016 41856 17032 41920
rect 17096 41856 17112 41920
rect 17176 41856 17192 41920
rect 17256 41856 17262 41920
rect 16946 41855 17262 41856
rect 21946 41920 22262 41921
rect 21946 41856 21952 41920
rect 22016 41856 22032 41920
rect 22096 41856 22112 41920
rect 22176 41856 22192 41920
rect 22256 41856 22262 41920
rect 21946 41855 22262 41856
rect 26946 41920 27262 41921
rect 26946 41856 26952 41920
rect 27016 41856 27032 41920
rect 27096 41856 27112 41920
rect 27176 41856 27192 41920
rect 27256 41856 27262 41920
rect 26946 41855 27262 41856
rect 31946 41920 32262 41921
rect 31946 41856 31952 41920
rect 32016 41856 32032 41920
rect 32096 41856 32112 41920
rect 32176 41856 32192 41920
rect 32256 41856 32262 41920
rect 31946 41855 32262 41856
rect 36946 41920 37262 41921
rect 36946 41856 36952 41920
rect 37016 41856 37032 41920
rect 37096 41856 37112 41920
rect 37176 41856 37192 41920
rect 37256 41856 37262 41920
rect 36946 41855 37262 41856
rect 31702 41380 31708 41444
rect 31772 41442 31778 41444
rect 32438 41442 32444 41444
rect 31772 41382 32444 41442
rect 31772 41380 31778 41382
rect 32438 41380 32444 41382
rect 32508 41380 32514 41444
rect 2606 41376 2922 41377
rect 2606 41312 2612 41376
rect 2676 41312 2692 41376
rect 2756 41312 2772 41376
rect 2836 41312 2852 41376
rect 2916 41312 2922 41376
rect 2606 41311 2922 41312
rect 7606 41376 7922 41377
rect 7606 41312 7612 41376
rect 7676 41312 7692 41376
rect 7756 41312 7772 41376
rect 7836 41312 7852 41376
rect 7916 41312 7922 41376
rect 7606 41311 7922 41312
rect 12606 41376 12922 41377
rect 12606 41312 12612 41376
rect 12676 41312 12692 41376
rect 12756 41312 12772 41376
rect 12836 41312 12852 41376
rect 12916 41312 12922 41376
rect 12606 41311 12922 41312
rect 17606 41376 17922 41377
rect 17606 41312 17612 41376
rect 17676 41312 17692 41376
rect 17756 41312 17772 41376
rect 17836 41312 17852 41376
rect 17916 41312 17922 41376
rect 17606 41311 17922 41312
rect 22606 41376 22922 41377
rect 22606 41312 22612 41376
rect 22676 41312 22692 41376
rect 22756 41312 22772 41376
rect 22836 41312 22852 41376
rect 22916 41312 22922 41376
rect 22606 41311 22922 41312
rect 27606 41376 27922 41377
rect 27606 41312 27612 41376
rect 27676 41312 27692 41376
rect 27756 41312 27772 41376
rect 27836 41312 27852 41376
rect 27916 41312 27922 41376
rect 27606 41311 27922 41312
rect 32606 41376 32922 41377
rect 32606 41312 32612 41376
rect 32676 41312 32692 41376
rect 32756 41312 32772 41376
rect 32836 41312 32852 41376
rect 32916 41312 32922 41376
rect 32606 41311 32922 41312
rect 37606 41376 37922 41377
rect 37606 41312 37612 41376
rect 37676 41312 37692 41376
rect 37756 41312 37772 41376
rect 37836 41312 37852 41376
rect 37916 41312 37922 41376
rect 37606 41311 37922 41312
rect 1946 40832 2262 40833
rect 1946 40768 1952 40832
rect 2016 40768 2032 40832
rect 2096 40768 2112 40832
rect 2176 40768 2192 40832
rect 2256 40768 2262 40832
rect 1946 40767 2262 40768
rect 6946 40832 7262 40833
rect 6946 40768 6952 40832
rect 7016 40768 7032 40832
rect 7096 40768 7112 40832
rect 7176 40768 7192 40832
rect 7256 40768 7262 40832
rect 6946 40767 7262 40768
rect 11946 40832 12262 40833
rect 11946 40768 11952 40832
rect 12016 40768 12032 40832
rect 12096 40768 12112 40832
rect 12176 40768 12192 40832
rect 12256 40768 12262 40832
rect 11946 40767 12262 40768
rect 16946 40832 17262 40833
rect 16946 40768 16952 40832
rect 17016 40768 17032 40832
rect 17096 40768 17112 40832
rect 17176 40768 17192 40832
rect 17256 40768 17262 40832
rect 16946 40767 17262 40768
rect 21946 40832 22262 40833
rect 21946 40768 21952 40832
rect 22016 40768 22032 40832
rect 22096 40768 22112 40832
rect 22176 40768 22192 40832
rect 22256 40768 22262 40832
rect 21946 40767 22262 40768
rect 26946 40832 27262 40833
rect 26946 40768 26952 40832
rect 27016 40768 27032 40832
rect 27096 40768 27112 40832
rect 27176 40768 27192 40832
rect 27256 40768 27262 40832
rect 26946 40767 27262 40768
rect 31946 40832 32262 40833
rect 31946 40768 31952 40832
rect 32016 40768 32032 40832
rect 32096 40768 32112 40832
rect 32176 40768 32192 40832
rect 32256 40768 32262 40832
rect 31946 40767 32262 40768
rect 36946 40832 37262 40833
rect 36946 40768 36952 40832
rect 37016 40768 37032 40832
rect 37096 40768 37112 40832
rect 37176 40768 37192 40832
rect 37256 40768 37262 40832
rect 36946 40767 37262 40768
rect 2606 40288 2922 40289
rect 2606 40224 2612 40288
rect 2676 40224 2692 40288
rect 2756 40224 2772 40288
rect 2836 40224 2852 40288
rect 2916 40224 2922 40288
rect 2606 40223 2922 40224
rect 7606 40288 7922 40289
rect 7606 40224 7612 40288
rect 7676 40224 7692 40288
rect 7756 40224 7772 40288
rect 7836 40224 7852 40288
rect 7916 40224 7922 40288
rect 7606 40223 7922 40224
rect 12606 40288 12922 40289
rect 12606 40224 12612 40288
rect 12676 40224 12692 40288
rect 12756 40224 12772 40288
rect 12836 40224 12852 40288
rect 12916 40224 12922 40288
rect 12606 40223 12922 40224
rect 17606 40288 17922 40289
rect 17606 40224 17612 40288
rect 17676 40224 17692 40288
rect 17756 40224 17772 40288
rect 17836 40224 17852 40288
rect 17916 40224 17922 40288
rect 17606 40223 17922 40224
rect 22606 40288 22922 40289
rect 22606 40224 22612 40288
rect 22676 40224 22692 40288
rect 22756 40224 22772 40288
rect 22836 40224 22852 40288
rect 22916 40224 22922 40288
rect 22606 40223 22922 40224
rect 27606 40288 27922 40289
rect 27606 40224 27612 40288
rect 27676 40224 27692 40288
rect 27756 40224 27772 40288
rect 27836 40224 27852 40288
rect 27916 40224 27922 40288
rect 27606 40223 27922 40224
rect 32606 40288 32922 40289
rect 32606 40224 32612 40288
rect 32676 40224 32692 40288
rect 32756 40224 32772 40288
rect 32836 40224 32852 40288
rect 32916 40224 32922 40288
rect 32606 40223 32922 40224
rect 37606 40288 37922 40289
rect 37606 40224 37612 40288
rect 37676 40224 37692 40288
rect 37756 40224 37772 40288
rect 37836 40224 37852 40288
rect 37916 40224 37922 40288
rect 37606 40223 37922 40224
rect 1946 39744 2262 39745
rect 1946 39680 1952 39744
rect 2016 39680 2032 39744
rect 2096 39680 2112 39744
rect 2176 39680 2192 39744
rect 2256 39680 2262 39744
rect 1946 39679 2262 39680
rect 6946 39744 7262 39745
rect 6946 39680 6952 39744
rect 7016 39680 7032 39744
rect 7096 39680 7112 39744
rect 7176 39680 7192 39744
rect 7256 39680 7262 39744
rect 6946 39679 7262 39680
rect 11946 39744 12262 39745
rect 11946 39680 11952 39744
rect 12016 39680 12032 39744
rect 12096 39680 12112 39744
rect 12176 39680 12192 39744
rect 12256 39680 12262 39744
rect 11946 39679 12262 39680
rect 16946 39744 17262 39745
rect 16946 39680 16952 39744
rect 17016 39680 17032 39744
rect 17096 39680 17112 39744
rect 17176 39680 17192 39744
rect 17256 39680 17262 39744
rect 16946 39679 17262 39680
rect 21946 39744 22262 39745
rect 21946 39680 21952 39744
rect 22016 39680 22032 39744
rect 22096 39680 22112 39744
rect 22176 39680 22192 39744
rect 22256 39680 22262 39744
rect 21946 39679 22262 39680
rect 26946 39744 27262 39745
rect 26946 39680 26952 39744
rect 27016 39680 27032 39744
rect 27096 39680 27112 39744
rect 27176 39680 27192 39744
rect 27256 39680 27262 39744
rect 26946 39679 27262 39680
rect 31946 39744 32262 39745
rect 31946 39680 31952 39744
rect 32016 39680 32032 39744
rect 32096 39680 32112 39744
rect 32176 39680 32192 39744
rect 32256 39680 32262 39744
rect 31946 39679 32262 39680
rect 36946 39744 37262 39745
rect 36946 39680 36952 39744
rect 37016 39680 37032 39744
rect 37096 39680 37112 39744
rect 37176 39680 37192 39744
rect 37256 39680 37262 39744
rect 36946 39679 37262 39680
rect 2606 39200 2922 39201
rect 2606 39136 2612 39200
rect 2676 39136 2692 39200
rect 2756 39136 2772 39200
rect 2836 39136 2852 39200
rect 2916 39136 2922 39200
rect 2606 39135 2922 39136
rect 7606 39200 7922 39201
rect 7606 39136 7612 39200
rect 7676 39136 7692 39200
rect 7756 39136 7772 39200
rect 7836 39136 7852 39200
rect 7916 39136 7922 39200
rect 7606 39135 7922 39136
rect 12606 39200 12922 39201
rect 12606 39136 12612 39200
rect 12676 39136 12692 39200
rect 12756 39136 12772 39200
rect 12836 39136 12852 39200
rect 12916 39136 12922 39200
rect 12606 39135 12922 39136
rect 17606 39200 17922 39201
rect 17606 39136 17612 39200
rect 17676 39136 17692 39200
rect 17756 39136 17772 39200
rect 17836 39136 17852 39200
rect 17916 39136 17922 39200
rect 17606 39135 17922 39136
rect 22606 39200 22922 39201
rect 22606 39136 22612 39200
rect 22676 39136 22692 39200
rect 22756 39136 22772 39200
rect 22836 39136 22852 39200
rect 22916 39136 22922 39200
rect 22606 39135 22922 39136
rect 27606 39200 27922 39201
rect 27606 39136 27612 39200
rect 27676 39136 27692 39200
rect 27756 39136 27772 39200
rect 27836 39136 27852 39200
rect 27916 39136 27922 39200
rect 27606 39135 27922 39136
rect 32606 39200 32922 39201
rect 32606 39136 32612 39200
rect 32676 39136 32692 39200
rect 32756 39136 32772 39200
rect 32836 39136 32852 39200
rect 32916 39136 32922 39200
rect 32606 39135 32922 39136
rect 37606 39200 37922 39201
rect 37606 39136 37612 39200
rect 37676 39136 37692 39200
rect 37756 39136 37772 39200
rect 37836 39136 37852 39200
rect 37916 39136 37922 39200
rect 37606 39135 37922 39136
rect 1946 38656 2262 38657
rect 1946 38592 1952 38656
rect 2016 38592 2032 38656
rect 2096 38592 2112 38656
rect 2176 38592 2192 38656
rect 2256 38592 2262 38656
rect 1946 38591 2262 38592
rect 6946 38656 7262 38657
rect 6946 38592 6952 38656
rect 7016 38592 7032 38656
rect 7096 38592 7112 38656
rect 7176 38592 7192 38656
rect 7256 38592 7262 38656
rect 6946 38591 7262 38592
rect 11946 38656 12262 38657
rect 11946 38592 11952 38656
rect 12016 38592 12032 38656
rect 12096 38592 12112 38656
rect 12176 38592 12192 38656
rect 12256 38592 12262 38656
rect 11946 38591 12262 38592
rect 16946 38656 17262 38657
rect 16946 38592 16952 38656
rect 17016 38592 17032 38656
rect 17096 38592 17112 38656
rect 17176 38592 17192 38656
rect 17256 38592 17262 38656
rect 16946 38591 17262 38592
rect 21946 38656 22262 38657
rect 21946 38592 21952 38656
rect 22016 38592 22032 38656
rect 22096 38592 22112 38656
rect 22176 38592 22192 38656
rect 22256 38592 22262 38656
rect 21946 38591 22262 38592
rect 26946 38656 27262 38657
rect 26946 38592 26952 38656
rect 27016 38592 27032 38656
rect 27096 38592 27112 38656
rect 27176 38592 27192 38656
rect 27256 38592 27262 38656
rect 26946 38591 27262 38592
rect 31946 38656 32262 38657
rect 31946 38592 31952 38656
rect 32016 38592 32032 38656
rect 32096 38592 32112 38656
rect 32176 38592 32192 38656
rect 32256 38592 32262 38656
rect 31946 38591 32262 38592
rect 36946 38656 37262 38657
rect 36946 38592 36952 38656
rect 37016 38592 37032 38656
rect 37096 38592 37112 38656
rect 37176 38592 37192 38656
rect 37256 38592 37262 38656
rect 36946 38591 37262 38592
rect 2606 38112 2922 38113
rect 2606 38048 2612 38112
rect 2676 38048 2692 38112
rect 2756 38048 2772 38112
rect 2836 38048 2852 38112
rect 2916 38048 2922 38112
rect 2606 38047 2922 38048
rect 7606 38112 7922 38113
rect 7606 38048 7612 38112
rect 7676 38048 7692 38112
rect 7756 38048 7772 38112
rect 7836 38048 7852 38112
rect 7916 38048 7922 38112
rect 7606 38047 7922 38048
rect 12606 38112 12922 38113
rect 12606 38048 12612 38112
rect 12676 38048 12692 38112
rect 12756 38048 12772 38112
rect 12836 38048 12852 38112
rect 12916 38048 12922 38112
rect 12606 38047 12922 38048
rect 17606 38112 17922 38113
rect 17606 38048 17612 38112
rect 17676 38048 17692 38112
rect 17756 38048 17772 38112
rect 17836 38048 17852 38112
rect 17916 38048 17922 38112
rect 17606 38047 17922 38048
rect 22606 38112 22922 38113
rect 22606 38048 22612 38112
rect 22676 38048 22692 38112
rect 22756 38048 22772 38112
rect 22836 38048 22852 38112
rect 22916 38048 22922 38112
rect 22606 38047 22922 38048
rect 27606 38112 27922 38113
rect 27606 38048 27612 38112
rect 27676 38048 27692 38112
rect 27756 38048 27772 38112
rect 27836 38048 27852 38112
rect 27916 38048 27922 38112
rect 27606 38047 27922 38048
rect 32606 38112 32922 38113
rect 32606 38048 32612 38112
rect 32676 38048 32692 38112
rect 32756 38048 32772 38112
rect 32836 38048 32852 38112
rect 32916 38048 32922 38112
rect 32606 38047 32922 38048
rect 37606 38112 37922 38113
rect 37606 38048 37612 38112
rect 37676 38048 37692 38112
rect 37756 38048 37772 38112
rect 37836 38048 37852 38112
rect 37916 38048 37922 38112
rect 37606 38047 37922 38048
rect 1946 37568 2262 37569
rect 1946 37504 1952 37568
rect 2016 37504 2032 37568
rect 2096 37504 2112 37568
rect 2176 37504 2192 37568
rect 2256 37504 2262 37568
rect 1946 37503 2262 37504
rect 6946 37568 7262 37569
rect 6946 37504 6952 37568
rect 7016 37504 7032 37568
rect 7096 37504 7112 37568
rect 7176 37504 7192 37568
rect 7256 37504 7262 37568
rect 6946 37503 7262 37504
rect 11946 37568 12262 37569
rect 11946 37504 11952 37568
rect 12016 37504 12032 37568
rect 12096 37504 12112 37568
rect 12176 37504 12192 37568
rect 12256 37504 12262 37568
rect 11946 37503 12262 37504
rect 16946 37568 17262 37569
rect 16946 37504 16952 37568
rect 17016 37504 17032 37568
rect 17096 37504 17112 37568
rect 17176 37504 17192 37568
rect 17256 37504 17262 37568
rect 16946 37503 17262 37504
rect 21946 37568 22262 37569
rect 21946 37504 21952 37568
rect 22016 37504 22032 37568
rect 22096 37504 22112 37568
rect 22176 37504 22192 37568
rect 22256 37504 22262 37568
rect 21946 37503 22262 37504
rect 26946 37568 27262 37569
rect 26946 37504 26952 37568
rect 27016 37504 27032 37568
rect 27096 37504 27112 37568
rect 27176 37504 27192 37568
rect 27256 37504 27262 37568
rect 26946 37503 27262 37504
rect 31946 37568 32262 37569
rect 31946 37504 31952 37568
rect 32016 37504 32032 37568
rect 32096 37504 32112 37568
rect 32176 37504 32192 37568
rect 32256 37504 32262 37568
rect 31946 37503 32262 37504
rect 36946 37568 37262 37569
rect 36946 37504 36952 37568
rect 37016 37504 37032 37568
rect 37096 37504 37112 37568
rect 37176 37504 37192 37568
rect 37256 37504 37262 37568
rect 36946 37503 37262 37504
rect 2606 37024 2922 37025
rect 2606 36960 2612 37024
rect 2676 36960 2692 37024
rect 2756 36960 2772 37024
rect 2836 36960 2852 37024
rect 2916 36960 2922 37024
rect 2606 36959 2922 36960
rect 7606 37024 7922 37025
rect 7606 36960 7612 37024
rect 7676 36960 7692 37024
rect 7756 36960 7772 37024
rect 7836 36960 7852 37024
rect 7916 36960 7922 37024
rect 7606 36959 7922 36960
rect 12606 37024 12922 37025
rect 12606 36960 12612 37024
rect 12676 36960 12692 37024
rect 12756 36960 12772 37024
rect 12836 36960 12852 37024
rect 12916 36960 12922 37024
rect 12606 36959 12922 36960
rect 17606 37024 17922 37025
rect 17606 36960 17612 37024
rect 17676 36960 17692 37024
rect 17756 36960 17772 37024
rect 17836 36960 17852 37024
rect 17916 36960 17922 37024
rect 17606 36959 17922 36960
rect 22606 37024 22922 37025
rect 22606 36960 22612 37024
rect 22676 36960 22692 37024
rect 22756 36960 22772 37024
rect 22836 36960 22852 37024
rect 22916 36960 22922 37024
rect 22606 36959 22922 36960
rect 27606 37024 27922 37025
rect 27606 36960 27612 37024
rect 27676 36960 27692 37024
rect 27756 36960 27772 37024
rect 27836 36960 27852 37024
rect 27916 36960 27922 37024
rect 27606 36959 27922 36960
rect 32606 37024 32922 37025
rect 32606 36960 32612 37024
rect 32676 36960 32692 37024
rect 32756 36960 32772 37024
rect 32836 36960 32852 37024
rect 32916 36960 32922 37024
rect 32606 36959 32922 36960
rect 37606 37024 37922 37025
rect 37606 36960 37612 37024
rect 37676 36960 37692 37024
rect 37756 36960 37772 37024
rect 37836 36960 37852 37024
rect 37916 36960 37922 37024
rect 37606 36959 37922 36960
rect 1946 36480 2262 36481
rect 1946 36416 1952 36480
rect 2016 36416 2032 36480
rect 2096 36416 2112 36480
rect 2176 36416 2192 36480
rect 2256 36416 2262 36480
rect 1946 36415 2262 36416
rect 6946 36480 7262 36481
rect 6946 36416 6952 36480
rect 7016 36416 7032 36480
rect 7096 36416 7112 36480
rect 7176 36416 7192 36480
rect 7256 36416 7262 36480
rect 6946 36415 7262 36416
rect 11946 36480 12262 36481
rect 11946 36416 11952 36480
rect 12016 36416 12032 36480
rect 12096 36416 12112 36480
rect 12176 36416 12192 36480
rect 12256 36416 12262 36480
rect 11946 36415 12262 36416
rect 16946 36480 17262 36481
rect 16946 36416 16952 36480
rect 17016 36416 17032 36480
rect 17096 36416 17112 36480
rect 17176 36416 17192 36480
rect 17256 36416 17262 36480
rect 16946 36415 17262 36416
rect 21946 36480 22262 36481
rect 21946 36416 21952 36480
rect 22016 36416 22032 36480
rect 22096 36416 22112 36480
rect 22176 36416 22192 36480
rect 22256 36416 22262 36480
rect 21946 36415 22262 36416
rect 26946 36480 27262 36481
rect 26946 36416 26952 36480
rect 27016 36416 27032 36480
rect 27096 36416 27112 36480
rect 27176 36416 27192 36480
rect 27256 36416 27262 36480
rect 26946 36415 27262 36416
rect 31946 36480 32262 36481
rect 31946 36416 31952 36480
rect 32016 36416 32032 36480
rect 32096 36416 32112 36480
rect 32176 36416 32192 36480
rect 32256 36416 32262 36480
rect 31946 36415 32262 36416
rect 36946 36480 37262 36481
rect 36946 36416 36952 36480
rect 37016 36416 37032 36480
rect 37096 36416 37112 36480
rect 37176 36416 37192 36480
rect 37256 36416 37262 36480
rect 36946 36415 37262 36416
rect 18086 36138 18092 36140
rect 2454 36078 18092 36138
rect 0 36002 800 36032
rect 2454 36002 2514 36078
rect 18086 36076 18092 36078
rect 18156 36076 18162 36140
rect 0 35942 2514 36002
rect 40493 36002 40559 36005
rect 41200 36002 42000 36032
rect 40493 36000 42000 36002
rect 40493 35944 40498 36000
rect 40554 35944 42000 36000
rect 40493 35942 42000 35944
rect 0 35912 800 35942
rect 40493 35939 40559 35942
rect 2606 35936 2922 35937
rect 2606 35872 2612 35936
rect 2676 35872 2692 35936
rect 2756 35872 2772 35936
rect 2836 35872 2852 35936
rect 2916 35872 2922 35936
rect 2606 35871 2922 35872
rect 7606 35936 7922 35937
rect 7606 35872 7612 35936
rect 7676 35872 7692 35936
rect 7756 35872 7772 35936
rect 7836 35872 7852 35936
rect 7916 35872 7922 35936
rect 7606 35871 7922 35872
rect 12606 35936 12922 35937
rect 12606 35872 12612 35936
rect 12676 35872 12692 35936
rect 12756 35872 12772 35936
rect 12836 35872 12852 35936
rect 12916 35872 12922 35936
rect 12606 35871 12922 35872
rect 17606 35936 17922 35937
rect 17606 35872 17612 35936
rect 17676 35872 17692 35936
rect 17756 35872 17772 35936
rect 17836 35872 17852 35936
rect 17916 35872 17922 35936
rect 17606 35871 17922 35872
rect 22606 35936 22922 35937
rect 22606 35872 22612 35936
rect 22676 35872 22692 35936
rect 22756 35872 22772 35936
rect 22836 35872 22852 35936
rect 22916 35872 22922 35936
rect 22606 35871 22922 35872
rect 27606 35936 27922 35937
rect 27606 35872 27612 35936
rect 27676 35872 27692 35936
rect 27756 35872 27772 35936
rect 27836 35872 27852 35936
rect 27916 35872 27922 35936
rect 27606 35871 27922 35872
rect 32606 35936 32922 35937
rect 32606 35872 32612 35936
rect 32676 35872 32692 35936
rect 32756 35872 32772 35936
rect 32836 35872 32852 35936
rect 32916 35872 32922 35936
rect 32606 35871 32922 35872
rect 37606 35936 37922 35937
rect 37606 35872 37612 35936
rect 37676 35872 37692 35936
rect 37756 35872 37772 35936
rect 37836 35872 37852 35936
rect 37916 35872 37922 35936
rect 41200 35912 42000 35942
rect 37606 35871 37922 35872
rect 1946 35392 2262 35393
rect 1946 35328 1952 35392
rect 2016 35328 2032 35392
rect 2096 35328 2112 35392
rect 2176 35328 2192 35392
rect 2256 35328 2262 35392
rect 1946 35327 2262 35328
rect 6946 35392 7262 35393
rect 6946 35328 6952 35392
rect 7016 35328 7032 35392
rect 7096 35328 7112 35392
rect 7176 35328 7192 35392
rect 7256 35328 7262 35392
rect 6946 35327 7262 35328
rect 11946 35392 12262 35393
rect 11946 35328 11952 35392
rect 12016 35328 12032 35392
rect 12096 35328 12112 35392
rect 12176 35328 12192 35392
rect 12256 35328 12262 35392
rect 11946 35327 12262 35328
rect 16946 35392 17262 35393
rect 16946 35328 16952 35392
rect 17016 35328 17032 35392
rect 17096 35328 17112 35392
rect 17176 35328 17192 35392
rect 17256 35328 17262 35392
rect 16946 35327 17262 35328
rect 21946 35392 22262 35393
rect 21946 35328 21952 35392
rect 22016 35328 22032 35392
rect 22096 35328 22112 35392
rect 22176 35328 22192 35392
rect 22256 35328 22262 35392
rect 21946 35327 22262 35328
rect 26946 35392 27262 35393
rect 26946 35328 26952 35392
rect 27016 35328 27032 35392
rect 27096 35328 27112 35392
rect 27176 35328 27192 35392
rect 27256 35328 27262 35392
rect 26946 35327 27262 35328
rect 31946 35392 32262 35393
rect 31946 35328 31952 35392
rect 32016 35328 32032 35392
rect 32096 35328 32112 35392
rect 32176 35328 32192 35392
rect 32256 35328 32262 35392
rect 31946 35327 32262 35328
rect 36946 35392 37262 35393
rect 36946 35328 36952 35392
rect 37016 35328 37032 35392
rect 37096 35328 37112 35392
rect 37176 35328 37192 35392
rect 37256 35328 37262 35392
rect 36946 35327 37262 35328
rect 2606 34848 2922 34849
rect 2606 34784 2612 34848
rect 2676 34784 2692 34848
rect 2756 34784 2772 34848
rect 2836 34784 2852 34848
rect 2916 34784 2922 34848
rect 2606 34783 2922 34784
rect 7606 34848 7922 34849
rect 7606 34784 7612 34848
rect 7676 34784 7692 34848
rect 7756 34784 7772 34848
rect 7836 34784 7852 34848
rect 7916 34784 7922 34848
rect 7606 34783 7922 34784
rect 12606 34848 12922 34849
rect 12606 34784 12612 34848
rect 12676 34784 12692 34848
rect 12756 34784 12772 34848
rect 12836 34784 12852 34848
rect 12916 34784 12922 34848
rect 12606 34783 12922 34784
rect 17606 34848 17922 34849
rect 17606 34784 17612 34848
rect 17676 34784 17692 34848
rect 17756 34784 17772 34848
rect 17836 34784 17852 34848
rect 17916 34784 17922 34848
rect 17606 34783 17922 34784
rect 22606 34848 22922 34849
rect 22606 34784 22612 34848
rect 22676 34784 22692 34848
rect 22756 34784 22772 34848
rect 22836 34784 22852 34848
rect 22916 34784 22922 34848
rect 22606 34783 22922 34784
rect 27606 34848 27922 34849
rect 27606 34784 27612 34848
rect 27676 34784 27692 34848
rect 27756 34784 27772 34848
rect 27836 34784 27852 34848
rect 27916 34784 27922 34848
rect 27606 34783 27922 34784
rect 32606 34848 32922 34849
rect 32606 34784 32612 34848
rect 32676 34784 32692 34848
rect 32756 34784 32772 34848
rect 32836 34784 32852 34848
rect 32916 34784 32922 34848
rect 32606 34783 32922 34784
rect 37606 34848 37922 34849
rect 37606 34784 37612 34848
rect 37676 34784 37692 34848
rect 37756 34784 37772 34848
rect 37836 34784 37852 34848
rect 37916 34784 37922 34848
rect 37606 34783 37922 34784
rect 18086 34444 18092 34508
rect 18156 34506 18162 34508
rect 19609 34506 19675 34509
rect 18156 34504 19675 34506
rect 18156 34448 19614 34504
rect 19670 34448 19675 34504
rect 18156 34446 19675 34448
rect 18156 34444 18162 34446
rect 19609 34443 19675 34446
rect 1946 34304 2262 34305
rect 1946 34240 1952 34304
rect 2016 34240 2032 34304
rect 2096 34240 2112 34304
rect 2176 34240 2192 34304
rect 2256 34240 2262 34304
rect 1946 34239 2262 34240
rect 6946 34304 7262 34305
rect 6946 34240 6952 34304
rect 7016 34240 7032 34304
rect 7096 34240 7112 34304
rect 7176 34240 7192 34304
rect 7256 34240 7262 34304
rect 6946 34239 7262 34240
rect 11946 34304 12262 34305
rect 11946 34240 11952 34304
rect 12016 34240 12032 34304
rect 12096 34240 12112 34304
rect 12176 34240 12192 34304
rect 12256 34240 12262 34304
rect 11946 34239 12262 34240
rect 16946 34304 17262 34305
rect 16946 34240 16952 34304
rect 17016 34240 17032 34304
rect 17096 34240 17112 34304
rect 17176 34240 17192 34304
rect 17256 34240 17262 34304
rect 16946 34239 17262 34240
rect 21946 34304 22262 34305
rect 21946 34240 21952 34304
rect 22016 34240 22032 34304
rect 22096 34240 22112 34304
rect 22176 34240 22192 34304
rect 22256 34240 22262 34304
rect 21946 34239 22262 34240
rect 26946 34304 27262 34305
rect 26946 34240 26952 34304
rect 27016 34240 27032 34304
rect 27096 34240 27112 34304
rect 27176 34240 27192 34304
rect 27256 34240 27262 34304
rect 26946 34239 27262 34240
rect 31946 34304 32262 34305
rect 31946 34240 31952 34304
rect 32016 34240 32032 34304
rect 32096 34240 32112 34304
rect 32176 34240 32192 34304
rect 32256 34240 32262 34304
rect 31946 34239 32262 34240
rect 36946 34304 37262 34305
rect 36946 34240 36952 34304
rect 37016 34240 37032 34304
rect 37096 34240 37112 34304
rect 37176 34240 37192 34304
rect 37256 34240 37262 34304
rect 36946 34239 37262 34240
rect 21081 33828 21147 33829
rect 21030 33764 21036 33828
rect 21100 33826 21147 33828
rect 21100 33824 21192 33826
rect 21142 33768 21192 33824
rect 21100 33766 21192 33768
rect 21100 33764 21147 33766
rect 21081 33763 21147 33764
rect 2606 33760 2922 33761
rect 2606 33696 2612 33760
rect 2676 33696 2692 33760
rect 2756 33696 2772 33760
rect 2836 33696 2852 33760
rect 2916 33696 2922 33760
rect 2606 33695 2922 33696
rect 7606 33760 7922 33761
rect 7606 33696 7612 33760
rect 7676 33696 7692 33760
rect 7756 33696 7772 33760
rect 7836 33696 7852 33760
rect 7916 33696 7922 33760
rect 7606 33695 7922 33696
rect 12606 33760 12922 33761
rect 12606 33696 12612 33760
rect 12676 33696 12692 33760
rect 12756 33696 12772 33760
rect 12836 33696 12852 33760
rect 12916 33696 12922 33760
rect 12606 33695 12922 33696
rect 17606 33760 17922 33761
rect 17606 33696 17612 33760
rect 17676 33696 17692 33760
rect 17756 33696 17772 33760
rect 17836 33696 17852 33760
rect 17916 33696 17922 33760
rect 17606 33695 17922 33696
rect 22606 33760 22922 33761
rect 22606 33696 22612 33760
rect 22676 33696 22692 33760
rect 22756 33696 22772 33760
rect 22836 33696 22852 33760
rect 22916 33696 22922 33760
rect 22606 33695 22922 33696
rect 27606 33760 27922 33761
rect 27606 33696 27612 33760
rect 27676 33696 27692 33760
rect 27756 33696 27772 33760
rect 27836 33696 27852 33760
rect 27916 33696 27922 33760
rect 27606 33695 27922 33696
rect 32606 33760 32922 33761
rect 32606 33696 32612 33760
rect 32676 33696 32692 33760
rect 32756 33696 32772 33760
rect 32836 33696 32852 33760
rect 32916 33696 32922 33760
rect 32606 33695 32922 33696
rect 37606 33760 37922 33761
rect 37606 33696 37612 33760
rect 37676 33696 37692 33760
rect 37756 33696 37772 33760
rect 37836 33696 37852 33760
rect 37916 33696 37922 33760
rect 37606 33695 37922 33696
rect 1946 33216 2262 33217
rect 1946 33152 1952 33216
rect 2016 33152 2032 33216
rect 2096 33152 2112 33216
rect 2176 33152 2192 33216
rect 2256 33152 2262 33216
rect 1946 33151 2262 33152
rect 6946 33216 7262 33217
rect 6946 33152 6952 33216
rect 7016 33152 7032 33216
rect 7096 33152 7112 33216
rect 7176 33152 7192 33216
rect 7256 33152 7262 33216
rect 6946 33151 7262 33152
rect 11946 33216 12262 33217
rect 11946 33152 11952 33216
rect 12016 33152 12032 33216
rect 12096 33152 12112 33216
rect 12176 33152 12192 33216
rect 12256 33152 12262 33216
rect 11946 33151 12262 33152
rect 16946 33216 17262 33217
rect 16946 33152 16952 33216
rect 17016 33152 17032 33216
rect 17096 33152 17112 33216
rect 17176 33152 17192 33216
rect 17256 33152 17262 33216
rect 16946 33151 17262 33152
rect 21946 33216 22262 33217
rect 21946 33152 21952 33216
rect 22016 33152 22032 33216
rect 22096 33152 22112 33216
rect 22176 33152 22192 33216
rect 22256 33152 22262 33216
rect 21946 33151 22262 33152
rect 26946 33216 27262 33217
rect 26946 33152 26952 33216
rect 27016 33152 27032 33216
rect 27096 33152 27112 33216
rect 27176 33152 27192 33216
rect 27256 33152 27262 33216
rect 26946 33151 27262 33152
rect 31946 33216 32262 33217
rect 31946 33152 31952 33216
rect 32016 33152 32032 33216
rect 32096 33152 32112 33216
rect 32176 33152 32192 33216
rect 32256 33152 32262 33216
rect 31946 33151 32262 33152
rect 36946 33216 37262 33217
rect 36946 33152 36952 33216
rect 37016 33152 37032 33216
rect 37096 33152 37112 33216
rect 37176 33152 37192 33216
rect 37256 33152 37262 33216
rect 36946 33151 37262 33152
rect 2606 32672 2922 32673
rect 2606 32608 2612 32672
rect 2676 32608 2692 32672
rect 2756 32608 2772 32672
rect 2836 32608 2852 32672
rect 2916 32608 2922 32672
rect 2606 32607 2922 32608
rect 7606 32672 7922 32673
rect 7606 32608 7612 32672
rect 7676 32608 7692 32672
rect 7756 32608 7772 32672
rect 7836 32608 7852 32672
rect 7916 32608 7922 32672
rect 7606 32607 7922 32608
rect 12606 32672 12922 32673
rect 12606 32608 12612 32672
rect 12676 32608 12692 32672
rect 12756 32608 12772 32672
rect 12836 32608 12852 32672
rect 12916 32608 12922 32672
rect 12606 32607 12922 32608
rect 17606 32672 17922 32673
rect 17606 32608 17612 32672
rect 17676 32608 17692 32672
rect 17756 32608 17772 32672
rect 17836 32608 17852 32672
rect 17916 32608 17922 32672
rect 17606 32607 17922 32608
rect 22606 32672 22922 32673
rect 22606 32608 22612 32672
rect 22676 32608 22692 32672
rect 22756 32608 22772 32672
rect 22836 32608 22852 32672
rect 22916 32608 22922 32672
rect 22606 32607 22922 32608
rect 27606 32672 27922 32673
rect 27606 32608 27612 32672
rect 27676 32608 27692 32672
rect 27756 32608 27772 32672
rect 27836 32608 27852 32672
rect 27916 32608 27922 32672
rect 27606 32607 27922 32608
rect 32606 32672 32922 32673
rect 32606 32608 32612 32672
rect 32676 32608 32692 32672
rect 32756 32608 32772 32672
rect 32836 32608 32852 32672
rect 32916 32608 32922 32672
rect 32606 32607 32922 32608
rect 37606 32672 37922 32673
rect 37606 32608 37612 32672
rect 37676 32608 37692 32672
rect 37756 32608 37772 32672
rect 37836 32608 37852 32672
rect 37916 32608 37922 32672
rect 37606 32607 37922 32608
rect 1946 32128 2262 32129
rect 1946 32064 1952 32128
rect 2016 32064 2032 32128
rect 2096 32064 2112 32128
rect 2176 32064 2192 32128
rect 2256 32064 2262 32128
rect 1946 32063 2262 32064
rect 6946 32128 7262 32129
rect 6946 32064 6952 32128
rect 7016 32064 7032 32128
rect 7096 32064 7112 32128
rect 7176 32064 7192 32128
rect 7256 32064 7262 32128
rect 6946 32063 7262 32064
rect 11946 32128 12262 32129
rect 11946 32064 11952 32128
rect 12016 32064 12032 32128
rect 12096 32064 12112 32128
rect 12176 32064 12192 32128
rect 12256 32064 12262 32128
rect 11946 32063 12262 32064
rect 16946 32128 17262 32129
rect 16946 32064 16952 32128
rect 17016 32064 17032 32128
rect 17096 32064 17112 32128
rect 17176 32064 17192 32128
rect 17256 32064 17262 32128
rect 16946 32063 17262 32064
rect 21946 32128 22262 32129
rect 21946 32064 21952 32128
rect 22016 32064 22032 32128
rect 22096 32064 22112 32128
rect 22176 32064 22192 32128
rect 22256 32064 22262 32128
rect 21946 32063 22262 32064
rect 26946 32128 27262 32129
rect 26946 32064 26952 32128
rect 27016 32064 27032 32128
rect 27096 32064 27112 32128
rect 27176 32064 27192 32128
rect 27256 32064 27262 32128
rect 26946 32063 27262 32064
rect 31946 32128 32262 32129
rect 31946 32064 31952 32128
rect 32016 32064 32032 32128
rect 32096 32064 32112 32128
rect 32176 32064 32192 32128
rect 32256 32064 32262 32128
rect 31946 32063 32262 32064
rect 36946 32128 37262 32129
rect 36946 32064 36952 32128
rect 37016 32064 37032 32128
rect 37096 32064 37112 32128
rect 37176 32064 37192 32128
rect 37256 32064 37262 32128
rect 36946 32063 37262 32064
rect 2606 31584 2922 31585
rect 2606 31520 2612 31584
rect 2676 31520 2692 31584
rect 2756 31520 2772 31584
rect 2836 31520 2852 31584
rect 2916 31520 2922 31584
rect 2606 31519 2922 31520
rect 7606 31584 7922 31585
rect 7606 31520 7612 31584
rect 7676 31520 7692 31584
rect 7756 31520 7772 31584
rect 7836 31520 7852 31584
rect 7916 31520 7922 31584
rect 7606 31519 7922 31520
rect 12606 31584 12922 31585
rect 12606 31520 12612 31584
rect 12676 31520 12692 31584
rect 12756 31520 12772 31584
rect 12836 31520 12852 31584
rect 12916 31520 12922 31584
rect 12606 31519 12922 31520
rect 17606 31584 17922 31585
rect 17606 31520 17612 31584
rect 17676 31520 17692 31584
rect 17756 31520 17772 31584
rect 17836 31520 17852 31584
rect 17916 31520 17922 31584
rect 17606 31519 17922 31520
rect 22606 31584 22922 31585
rect 22606 31520 22612 31584
rect 22676 31520 22692 31584
rect 22756 31520 22772 31584
rect 22836 31520 22852 31584
rect 22916 31520 22922 31584
rect 22606 31519 22922 31520
rect 27606 31584 27922 31585
rect 27606 31520 27612 31584
rect 27676 31520 27692 31584
rect 27756 31520 27772 31584
rect 27836 31520 27852 31584
rect 27916 31520 27922 31584
rect 27606 31519 27922 31520
rect 32606 31584 32922 31585
rect 32606 31520 32612 31584
rect 32676 31520 32692 31584
rect 32756 31520 32772 31584
rect 32836 31520 32852 31584
rect 32916 31520 32922 31584
rect 32606 31519 32922 31520
rect 37606 31584 37922 31585
rect 37606 31520 37612 31584
rect 37676 31520 37692 31584
rect 37756 31520 37772 31584
rect 37836 31520 37852 31584
rect 37916 31520 37922 31584
rect 37606 31519 37922 31520
rect 1946 31040 2262 31041
rect 1946 30976 1952 31040
rect 2016 30976 2032 31040
rect 2096 30976 2112 31040
rect 2176 30976 2192 31040
rect 2256 30976 2262 31040
rect 1946 30975 2262 30976
rect 6946 31040 7262 31041
rect 6946 30976 6952 31040
rect 7016 30976 7032 31040
rect 7096 30976 7112 31040
rect 7176 30976 7192 31040
rect 7256 30976 7262 31040
rect 6946 30975 7262 30976
rect 11946 31040 12262 31041
rect 11946 30976 11952 31040
rect 12016 30976 12032 31040
rect 12096 30976 12112 31040
rect 12176 30976 12192 31040
rect 12256 30976 12262 31040
rect 11946 30975 12262 30976
rect 16946 31040 17262 31041
rect 16946 30976 16952 31040
rect 17016 30976 17032 31040
rect 17096 30976 17112 31040
rect 17176 30976 17192 31040
rect 17256 30976 17262 31040
rect 16946 30975 17262 30976
rect 21946 31040 22262 31041
rect 21946 30976 21952 31040
rect 22016 30976 22032 31040
rect 22096 30976 22112 31040
rect 22176 30976 22192 31040
rect 22256 30976 22262 31040
rect 21946 30975 22262 30976
rect 26946 31040 27262 31041
rect 26946 30976 26952 31040
rect 27016 30976 27032 31040
rect 27096 30976 27112 31040
rect 27176 30976 27192 31040
rect 27256 30976 27262 31040
rect 26946 30975 27262 30976
rect 31946 31040 32262 31041
rect 31946 30976 31952 31040
rect 32016 30976 32032 31040
rect 32096 30976 32112 31040
rect 32176 30976 32192 31040
rect 32256 30976 32262 31040
rect 31946 30975 32262 30976
rect 36946 31040 37262 31041
rect 36946 30976 36952 31040
rect 37016 30976 37032 31040
rect 37096 30976 37112 31040
rect 37176 30976 37192 31040
rect 37256 30976 37262 31040
rect 36946 30975 37262 30976
rect 9029 30698 9095 30701
rect 39113 30698 39179 30701
rect 9029 30696 39179 30698
rect 9029 30640 9034 30696
rect 9090 30640 39118 30696
rect 39174 30640 39179 30696
rect 9029 30638 39179 30640
rect 9029 30635 9095 30638
rect 39113 30635 39179 30638
rect 2606 30496 2922 30497
rect 2606 30432 2612 30496
rect 2676 30432 2692 30496
rect 2756 30432 2772 30496
rect 2836 30432 2852 30496
rect 2916 30432 2922 30496
rect 2606 30431 2922 30432
rect 7606 30496 7922 30497
rect 7606 30432 7612 30496
rect 7676 30432 7692 30496
rect 7756 30432 7772 30496
rect 7836 30432 7852 30496
rect 7916 30432 7922 30496
rect 7606 30431 7922 30432
rect 12606 30496 12922 30497
rect 12606 30432 12612 30496
rect 12676 30432 12692 30496
rect 12756 30432 12772 30496
rect 12836 30432 12852 30496
rect 12916 30432 12922 30496
rect 12606 30431 12922 30432
rect 17606 30496 17922 30497
rect 17606 30432 17612 30496
rect 17676 30432 17692 30496
rect 17756 30432 17772 30496
rect 17836 30432 17852 30496
rect 17916 30432 17922 30496
rect 17606 30431 17922 30432
rect 22606 30496 22922 30497
rect 22606 30432 22612 30496
rect 22676 30432 22692 30496
rect 22756 30432 22772 30496
rect 22836 30432 22852 30496
rect 22916 30432 22922 30496
rect 22606 30431 22922 30432
rect 27606 30496 27922 30497
rect 27606 30432 27612 30496
rect 27676 30432 27692 30496
rect 27756 30432 27772 30496
rect 27836 30432 27852 30496
rect 27916 30432 27922 30496
rect 27606 30431 27922 30432
rect 32606 30496 32922 30497
rect 32606 30432 32612 30496
rect 32676 30432 32692 30496
rect 32756 30432 32772 30496
rect 32836 30432 32852 30496
rect 32916 30432 32922 30496
rect 32606 30431 32922 30432
rect 37606 30496 37922 30497
rect 37606 30432 37612 30496
rect 37676 30432 37692 30496
rect 37756 30432 37772 30496
rect 37836 30432 37852 30496
rect 37916 30432 37922 30496
rect 37606 30431 37922 30432
rect 1946 29952 2262 29953
rect 1946 29888 1952 29952
rect 2016 29888 2032 29952
rect 2096 29888 2112 29952
rect 2176 29888 2192 29952
rect 2256 29888 2262 29952
rect 1946 29887 2262 29888
rect 6946 29952 7262 29953
rect 6946 29888 6952 29952
rect 7016 29888 7032 29952
rect 7096 29888 7112 29952
rect 7176 29888 7192 29952
rect 7256 29888 7262 29952
rect 6946 29887 7262 29888
rect 11946 29952 12262 29953
rect 11946 29888 11952 29952
rect 12016 29888 12032 29952
rect 12096 29888 12112 29952
rect 12176 29888 12192 29952
rect 12256 29888 12262 29952
rect 11946 29887 12262 29888
rect 16946 29952 17262 29953
rect 16946 29888 16952 29952
rect 17016 29888 17032 29952
rect 17096 29888 17112 29952
rect 17176 29888 17192 29952
rect 17256 29888 17262 29952
rect 16946 29887 17262 29888
rect 21946 29952 22262 29953
rect 21946 29888 21952 29952
rect 22016 29888 22032 29952
rect 22096 29888 22112 29952
rect 22176 29888 22192 29952
rect 22256 29888 22262 29952
rect 21946 29887 22262 29888
rect 26946 29952 27262 29953
rect 26946 29888 26952 29952
rect 27016 29888 27032 29952
rect 27096 29888 27112 29952
rect 27176 29888 27192 29952
rect 27256 29888 27262 29952
rect 26946 29887 27262 29888
rect 31946 29952 32262 29953
rect 31946 29888 31952 29952
rect 32016 29888 32032 29952
rect 32096 29888 32112 29952
rect 32176 29888 32192 29952
rect 32256 29888 32262 29952
rect 31946 29887 32262 29888
rect 36946 29952 37262 29953
rect 36946 29888 36952 29952
rect 37016 29888 37032 29952
rect 37096 29888 37112 29952
rect 37176 29888 37192 29952
rect 37256 29888 37262 29952
rect 36946 29887 37262 29888
rect 2606 29408 2922 29409
rect 2606 29344 2612 29408
rect 2676 29344 2692 29408
rect 2756 29344 2772 29408
rect 2836 29344 2852 29408
rect 2916 29344 2922 29408
rect 2606 29343 2922 29344
rect 7606 29408 7922 29409
rect 7606 29344 7612 29408
rect 7676 29344 7692 29408
rect 7756 29344 7772 29408
rect 7836 29344 7852 29408
rect 7916 29344 7922 29408
rect 7606 29343 7922 29344
rect 12606 29408 12922 29409
rect 12606 29344 12612 29408
rect 12676 29344 12692 29408
rect 12756 29344 12772 29408
rect 12836 29344 12852 29408
rect 12916 29344 12922 29408
rect 12606 29343 12922 29344
rect 17606 29408 17922 29409
rect 17606 29344 17612 29408
rect 17676 29344 17692 29408
rect 17756 29344 17772 29408
rect 17836 29344 17852 29408
rect 17916 29344 17922 29408
rect 17606 29343 17922 29344
rect 22606 29408 22922 29409
rect 22606 29344 22612 29408
rect 22676 29344 22692 29408
rect 22756 29344 22772 29408
rect 22836 29344 22852 29408
rect 22916 29344 22922 29408
rect 22606 29343 22922 29344
rect 27606 29408 27922 29409
rect 27606 29344 27612 29408
rect 27676 29344 27692 29408
rect 27756 29344 27772 29408
rect 27836 29344 27852 29408
rect 27916 29344 27922 29408
rect 27606 29343 27922 29344
rect 32606 29408 32922 29409
rect 32606 29344 32612 29408
rect 32676 29344 32692 29408
rect 32756 29344 32772 29408
rect 32836 29344 32852 29408
rect 32916 29344 32922 29408
rect 32606 29343 32922 29344
rect 37606 29408 37922 29409
rect 37606 29344 37612 29408
rect 37676 29344 37692 29408
rect 37756 29344 37772 29408
rect 37836 29344 37852 29408
rect 37916 29344 37922 29408
rect 37606 29343 37922 29344
rect 1946 28864 2262 28865
rect 1946 28800 1952 28864
rect 2016 28800 2032 28864
rect 2096 28800 2112 28864
rect 2176 28800 2192 28864
rect 2256 28800 2262 28864
rect 1946 28799 2262 28800
rect 6946 28864 7262 28865
rect 6946 28800 6952 28864
rect 7016 28800 7032 28864
rect 7096 28800 7112 28864
rect 7176 28800 7192 28864
rect 7256 28800 7262 28864
rect 6946 28799 7262 28800
rect 11946 28864 12262 28865
rect 11946 28800 11952 28864
rect 12016 28800 12032 28864
rect 12096 28800 12112 28864
rect 12176 28800 12192 28864
rect 12256 28800 12262 28864
rect 11946 28799 12262 28800
rect 16946 28864 17262 28865
rect 16946 28800 16952 28864
rect 17016 28800 17032 28864
rect 17096 28800 17112 28864
rect 17176 28800 17192 28864
rect 17256 28800 17262 28864
rect 16946 28799 17262 28800
rect 21946 28864 22262 28865
rect 21946 28800 21952 28864
rect 22016 28800 22032 28864
rect 22096 28800 22112 28864
rect 22176 28800 22192 28864
rect 22256 28800 22262 28864
rect 21946 28799 22262 28800
rect 26946 28864 27262 28865
rect 26946 28800 26952 28864
rect 27016 28800 27032 28864
rect 27096 28800 27112 28864
rect 27176 28800 27192 28864
rect 27256 28800 27262 28864
rect 26946 28799 27262 28800
rect 31946 28864 32262 28865
rect 31946 28800 31952 28864
rect 32016 28800 32032 28864
rect 32096 28800 32112 28864
rect 32176 28800 32192 28864
rect 32256 28800 32262 28864
rect 31946 28799 32262 28800
rect 36946 28864 37262 28865
rect 36946 28800 36952 28864
rect 37016 28800 37032 28864
rect 37096 28800 37112 28864
rect 37176 28800 37192 28864
rect 37256 28800 37262 28864
rect 36946 28799 37262 28800
rect 30557 28794 30623 28797
rect 31702 28794 31708 28796
rect 30557 28792 31708 28794
rect 30557 28736 30562 28792
rect 30618 28736 31708 28792
rect 30557 28734 31708 28736
rect 30557 28731 30623 28734
rect 31702 28732 31708 28734
rect 31772 28732 31778 28796
rect 2606 28320 2922 28321
rect 2606 28256 2612 28320
rect 2676 28256 2692 28320
rect 2756 28256 2772 28320
rect 2836 28256 2852 28320
rect 2916 28256 2922 28320
rect 2606 28255 2922 28256
rect 7606 28320 7922 28321
rect 7606 28256 7612 28320
rect 7676 28256 7692 28320
rect 7756 28256 7772 28320
rect 7836 28256 7852 28320
rect 7916 28256 7922 28320
rect 7606 28255 7922 28256
rect 12606 28320 12922 28321
rect 12606 28256 12612 28320
rect 12676 28256 12692 28320
rect 12756 28256 12772 28320
rect 12836 28256 12852 28320
rect 12916 28256 12922 28320
rect 12606 28255 12922 28256
rect 17606 28320 17922 28321
rect 17606 28256 17612 28320
rect 17676 28256 17692 28320
rect 17756 28256 17772 28320
rect 17836 28256 17852 28320
rect 17916 28256 17922 28320
rect 17606 28255 17922 28256
rect 22606 28320 22922 28321
rect 22606 28256 22612 28320
rect 22676 28256 22692 28320
rect 22756 28256 22772 28320
rect 22836 28256 22852 28320
rect 22916 28256 22922 28320
rect 22606 28255 22922 28256
rect 27606 28320 27922 28321
rect 27606 28256 27612 28320
rect 27676 28256 27692 28320
rect 27756 28256 27772 28320
rect 27836 28256 27852 28320
rect 27916 28256 27922 28320
rect 27606 28255 27922 28256
rect 32606 28320 32922 28321
rect 32606 28256 32612 28320
rect 32676 28256 32692 28320
rect 32756 28256 32772 28320
rect 32836 28256 32852 28320
rect 32916 28256 32922 28320
rect 32606 28255 32922 28256
rect 37606 28320 37922 28321
rect 37606 28256 37612 28320
rect 37676 28256 37692 28320
rect 37756 28256 37772 28320
rect 37836 28256 37852 28320
rect 37916 28256 37922 28320
rect 37606 28255 37922 28256
rect 1946 27776 2262 27777
rect 1946 27712 1952 27776
rect 2016 27712 2032 27776
rect 2096 27712 2112 27776
rect 2176 27712 2192 27776
rect 2256 27712 2262 27776
rect 1946 27711 2262 27712
rect 6946 27776 7262 27777
rect 6946 27712 6952 27776
rect 7016 27712 7032 27776
rect 7096 27712 7112 27776
rect 7176 27712 7192 27776
rect 7256 27712 7262 27776
rect 6946 27711 7262 27712
rect 11946 27776 12262 27777
rect 11946 27712 11952 27776
rect 12016 27712 12032 27776
rect 12096 27712 12112 27776
rect 12176 27712 12192 27776
rect 12256 27712 12262 27776
rect 11946 27711 12262 27712
rect 16946 27776 17262 27777
rect 16946 27712 16952 27776
rect 17016 27712 17032 27776
rect 17096 27712 17112 27776
rect 17176 27712 17192 27776
rect 17256 27712 17262 27776
rect 16946 27711 17262 27712
rect 21946 27776 22262 27777
rect 21946 27712 21952 27776
rect 22016 27712 22032 27776
rect 22096 27712 22112 27776
rect 22176 27712 22192 27776
rect 22256 27712 22262 27776
rect 21946 27711 22262 27712
rect 26946 27776 27262 27777
rect 26946 27712 26952 27776
rect 27016 27712 27032 27776
rect 27096 27712 27112 27776
rect 27176 27712 27192 27776
rect 27256 27712 27262 27776
rect 26946 27711 27262 27712
rect 31946 27776 32262 27777
rect 31946 27712 31952 27776
rect 32016 27712 32032 27776
rect 32096 27712 32112 27776
rect 32176 27712 32192 27776
rect 32256 27712 32262 27776
rect 31946 27711 32262 27712
rect 36946 27776 37262 27777
rect 36946 27712 36952 27776
rect 37016 27712 37032 27776
rect 37096 27712 37112 27776
rect 37176 27712 37192 27776
rect 37256 27712 37262 27776
rect 36946 27711 37262 27712
rect 2606 27232 2922 27233
rect 2606 27168 2612 27232
rect 2676 27168 2692 27232
rect 2756 27168 2772 27232
rect 2836 27168 2852 27232
rect 2916 27168 2922 27232
rect 2606 27167 2922 27168
rect 7606 27232 7922 27233
rect 7606 27168 7612 27232
rect 7676 27168 7692 27232
rect 7756 27168 7772 27232
rect 7836 27168 7852 27232
rect 7916 27168 7922 27232
rect 7606 27167 7922 27168
rect 12606 27232 12922 27233
rect 12606 27168 12612 27232
rect 12676 27168 12692 27232
rect 12756 27168 12772 27232
rect 12836 27168 12852 27232
rect 12916 27168 12922 27232
rect 12606 27167 12922 27168
rect 17606 27232 17922 27233
rect 17606 27168 17612 27232
rect 17676 27168 17692 27232
rect 17756 27168 17772 27232
rect 17836 27168 17852 27232
rect 17916 27168 17922 27232
rect 17606 27167 17922 27168
rect 22606 27232 22922 27233
rect 22606 27168 22612 27232
rect 22676 27168 22692 27232
rect 22756 27168 22772 27232
rect 22836 27168 22852 27232
rect 22916 27168 22922 27232
rect 22606 27167 22922 27168
rect 27606 27232 27922 27233
rect 27606 27168 27612 27232
rect 27676 27168 27692 27232
rect 27756 27168 27772 27232
rect 27836 27168 27852 27232
rect 27916 27168 27922 27232
rect 27606 27167 27922 27168
rect 32606 27232 32922 27233
rect 32606 27168 32612 27232
rect 32676 27168 32692 27232
rect 32756 27168 32772 27232
rect 32836 27168 32852 27232
rect 32916 27168 32922 27232
rect 32606 27167 32922 27168
rect 37606 27232 37922 27233
rect 37606 27168 37612 27232
rect 37676 27168 37692 27232
rect 37756 27168 37772 27232
rect 37836 27168 37852 27232
rect 37916 27168 37922 27232
rect 37606 27167 37922 27168
rect 1946 26688 2262 26689
rect 1946 26624 1952 26688
rect 2016 26624 2032 26688
rect 2096 26624 2112 26688
rect 2176 26624 2192 26688
rect 2256 26624 2262 26688
rect 1946 26623 2262 26624
rect 6946 26688 7262 26689
rect 6946 26624 6952 26688
rect 7016 26624 7032 26688
rect 7096 26624 7112 26688
rect 7176 26624 7192 26688
rect 7256 26624 7262 26688
rect 6946 26623 7262 26624
rect 11946 26688 12262 26689
rect 11946 26624 11952 26688
rect 12016 26624 12032 26688
rect 12096 26624 12112 26688
rect 12176 26624 12192 26688
rect 12256 26624 12262 26688
rect 11946 26623 12262 26624
rect 16946 26688 17262 26689
rect 16946 26624 16952 26688
rect 17016 26624 17032 26688
rect 17096 26624 17112 26688
rect 17176 26624 17192 26688
rect 17256 26624 17262 26688
rect 16946 26623 17262 26624
rect 21946 26688 22262 26689
rect 21946 26624 21952 26688
rect 22016 26624 22032 26688
rect 22096 26624 22112 26688
rect 22176 26624 22192 26688
rect 22256 26624 22262 26688
rect 21946 26623 22262 26624
rect 26946 26688 27262 26689
rect 26946 26624 26952 26688
rect 27016 26624 27032 26688
rect 27096 26624 27112 26688
rect 27176 26624 27192 26688
rect 27256 26624 27262 26688
rect 26946 26623 27262 26624
rect 31946 26688 32262 26689
rect 31946 26624 31952 26688
rect 32016 26624 32032 26688
rect 32096 26624 32112 26688
rect 32176 26624 32192 26688
rect 32256 26624 32262 26688
rect 31946 26623 32262 26624
rect 36946 26688 37262 26689
rect 36946 26624 36952 26688
rect 37016 26624 37032 26688
rect 37096 26624 37112 26688
rect 37176 26624 37192 26688
rect 37256 26624 37262 26688
rect 36946 26623 37262 26624
rect 2606 26144 2922 26145
rect 2606 26080 2612 26144
rect 2676 26080 2692 26144
rect 2756 26080 2772 26144
rect 2836 26080 2852 26144
rect 2916 26080 2922 26144
rect 2606 26079 2922 26080
rect 7606 26144 7922 26145
rect 7606 26080 7612 26144
rect 7676 26080 7692 26144
rect 7756 26080 7772 26144
rect 7836 26080 7852 26144
rect 7916 26080 7922 26144
rect 7606 26079 7922 26080
rect 12606 26144 12922 26145
rect 12606 26080 12612 26144
rect 12676 26080 12692 26144
rect 12756 26080 12772 26144
rect 12836 26080 12852 26144
rect 12916 26080 12922 26144
rect 12606 26079 12922 26080
rect 17606 26144 17922 26145
rect 17606 26080 17612 26144
rect 17676 26080 17692 26144
rect 17756 26080 17772 26144
rect 17836 26080 17852 26144
rect 17916 26080 17922 26144
rect 17606 26079 17922 26080
rect 22606 26144 22922 26145
rect 22606 26080 22612 26144
rect 22676 26080 22692 26144
rect 22756 26080 22772 26144
rect 22836 26080 22852 26144
rect 22916 26080 22922 26144
rect 22606 26079 22922 26080
rect 27606 26144 27922 26145
rect 27606 26080 27612 26144
rect 27676 26080 27692 26144
rect 27756 26080 27772 26144
rect 27836 26080 27852 26144
rect 27916 26080 27922 26144
rect 27606 26079 27922 26080
rect 32606 26144 32922 26145
rect 32606 26080 32612 26144
rect 32676 26080 32692 26144
rect 32756 26080 32772 26144
rect 32836 26080 32852 26144
rect 32916 26080 32922 26144
rect 32606 26079 32922 26080
rect 37606 26144 37922 26145
rect 37606 26080 37612 26144
rect 37676 26080 37692 26144
rect 37756 26080 37772 26144
rect 37836 26080 37852 26144
rect 37916 26080 37922 26144
rect 37606 26079 37922 26080
rect 1946 25600 2262 25601
rect 1946 25536 1952 25600
rect 2016 25536 2032 25600
rect 2096 25536 2112 25600
rect 2176 25536 2192 25600
rect 2256 25536 2262 25600
rect 1946 25535 2262 25536
rect 6946 25600 7262 25601
rect 6946 25536 6952 25600
rect 7016 25536 7032 25600
rect 7096 25536 7112 25600
rect 7176 25536 7192 25600
rect 7256 25536 7262 25600
rect 6946 25535 7262 25536
rect 11946 25600 12262 25601
rect 11946 25536 11952 25600
rect 12016 25536 12032 25600
rect 12096 25536 12112 25600
rect 12176 25536 12192 25600
rect 12256 25536 12262 25600
rect 11946 25535 12262 25536
rect 16946 25600 17262 25601
rect 16946 25536 16952 25600
rect 17016 25536 17032 25600
rect 17096 25536 17112 25600
rect 17176 25536 17192 25600
rect 17256 25536 17262 25600
rect 16946 25535 17262 25536
rect 21946 25600 22262 25601
rect 21946 25536 21952 25600
rect 22016 25536 22032 25600
rect 22096 25536 22112 25600
rect 22176 25536 22192 25600
rect 22256 25536 22262 25600
rect 21946 25535 22262 25536
rect 26946 25600 27262 25601
rect 26946 25536 26952 25600
rect 27016 25536 27032 25600
rect 27096 25536 27112 25600
rect 27176 25536 27192 25600
rect 27256 25536 27262 25600
rect 26946 25535 27262 25536
rect 31946 25600 32262 25601
rect 31946 25536 31952 25600
rect 32016 25536 32032 25600
rect 32096 25536 32112 25600
rect 32176 25536 32192 25600
rect 32256 25536 32262 25600
rect 31946 25535 32262 25536
rect 36946 25600 37262 25601
rect 36946 25536 36952 25600
rect 37016 25536 37032 25600
rect 37096 25536 37112 25600
rect 37176 25536 37192 25600
rect 37256 25536 37262 25600
rect 36946 25535 37262 25536
rect 2606 25056 2922 25057
rect 2606 24992 2612 25056
rect 2676 24992 2692 25056
rect 2756 24992 2772 25056
rect 2836 24992 2852 25056
rect 2916 24992 2922 25056
rect 2606 24991 2922 24992
rect 7606 25056 7922 25057
rect 7606 24992 7612 25056
rect 7676 24992 7692 25056
rect 7756 24992 7772 25056
rect 7836 24992 7852 25056
rect 7916 24992 7922 25056
rect 7606 24991 7922 24992
rect 12606 25056 12922 25057
rect 12606 24992 12612 25056
rect 12676 24992 12692 25056
rect 12756 24992 12772 25056
rect 12836 24992 12852 25056
rect 12916 24992 12922 25056
rect 12606 24991 12922 24992
rect 17606 25056 17922 25057
rect 17606 24992 17612 25056
rect 17676 24992 17692 25056
rect 17756 24992 17772 25056
rect 17836 24992 17852 25056
rect 17916 24992 17922 25056
rect 17606 24991 17922 24992
rect 22606 25056 22922 25057
rect 22606 24992 22612 25056
rect 22676 24992 22692 25056
rect 22756 24992 22772 25056
rect 22836 24992 22852 25056
rect 22916 24992 22922 25056
rect 22606 24991 22922 24992
rect 27606 25056 27922 25057
rect 27606 24992 27612 25056
rect 27676 24992 27692 25056
rect 27756 24992 27772 25056
rect 27836 24992 27852 25056
rect 27916 24992 27922 25056
rect 27606 24991 27922 24992
rect 32606 25056 32922 25057
rect 32606 24992 32612 25056
rect 32676 24992 32692 25056
rect 32756 24992 32772 25056
rect 32836 24992 32852 25056
rect 32916 24992 32922 25056
rect 32606 24991 32922 24992
rect 37606 25056 37922 25057
rect 37606 24992 37612 25056
rect 37676 24992 37692 25056
rect 37756 24992 37772 25056
rect 37836 24992 37852 25056
rect 37916 24992 37922 25056
rect 37606 24991 37922 24992
rect 1946 24512 2262 24513
rect 1946 24448 1952 24512
rect 2016 24448 2032 24512
rect 2096 24448 2112 24512
rect 2176 24448 2192 24512
rect 2256 24448 2262 24512
rect 1946 24447 2262 24448
rect 6946 24512 7262 24513
rect 6946 24448 6952 24512
rect 7016 24448 7032 24512
rect 7096 24448 7112 24512
rect 7176 24448 7192 24512
rect 7256 24448 7262 24512
rect 6946 24447 7262 24448
rect 11946 24512 12262 24513
rect 11946 24448 11952 24512
rect 12016 24448 12032 24512
rect 12096 24448 12112 24512
rect 12176 24448 12192 24512
rect 12256 24448 12262 24512
rect 11946 24447 12262 24448
rect 16946 24512 17262 24513
rect 16946 24448 16952 24512
rect 17016 24448 17032 24512
rect 17096 24448 17112 24512
rect 17176 24448 17192 24512
rect 17256 24448 17262 24512
rect 16946 24447 17262 24448
rect 21946 24512 22262 24513
rect 21946 24448 21952 24512
rect 22016 24448 22032 24512
rect 22096 24448 22112 24512
rect 22176 24448 22192 24512
rect 22256 24448 22262 24512
rect 21946 24447 22262 24448
rect 26946 24512 27262 24513
rect 26946 24448 26952 24512
rect 27016 24448 27032 24512
rect 27096 24448 27112 24512
rect 27176 24448 27192 24512
rect 27256 24448 27262 24512
rect 26946 24447 27262 24448
rect 31946 24512 32262 24513
rect 31946 24448 31952 24512
rect 32016 24448 32032 24512
rect 32096 24448 32112 24512
rect 32176 24448 32192 24512
rect 32256 24448 32262 24512
rect 31946 24447 32262 24448
rect 36946 24512 37262 24513
rect 36946 24448 36952 24512
rect 37016 24448 37032 24512
rect 37096 24448 37112 24512
rect 37176 24448 37192 24512
rect 37256 24448 37262 24512
rect 36946 24447 37262 24448
rect 2606 23968 2922 23969
rect 2606 23904 2612 23968
rect 2676 23904 2692 23968
rect 2756 23904 2772 23968
rect 2836 23904 2852 23968
rect 2916 23904 2922 23968
rect 2606 23903 2922 23904
rect 7606 23968 7922 23969
rect 7606 23904 7612 23968
rect 7676 23904 7692 23968
rect 7756 23904 7772 23968
rect 7836 23904 7852 23968
rect 7916 23904 7922 23968
rect 7606 23903 7922 23904
rect 12606 23968 12922 23969
rect 12606 23904 12612 23968
rect 12676 23904 12692 23968
rect 12756 23904 12772 23968
rect 12836 23904 12852 23968
rect 12916 23904 12922 23968
rect 12606 23903 12922 23904
rect 17606 23968 17922 23969
rect 17606 23904 17612 23968
rect 17676 23904 17692 23968
rect 17756 23904 17772 23968
rect 17836 23904 17852 23968
rect 17916 23904 17922 23968
rect 17606 23903 17922 23904
rect 22606 23968 22922 23969
rect 22606 23904 22612 23968
rect 22676 23904 22692 23968
rect 22756 23904 22772 23968
rect 22836 23904 22852 23968
rect 22916 23904 22922 23968
rect 22606 23903 22922 23904
rect 27606 23968 27922 23969
rect 27606 23904 27612 23968
rect 27676 23904 27692 23968
rect 27756 23904 27772 23968
rect 27836 23904 27852 23968
rect 27916 23904 27922 23968
rect 27606 23903 27922 23904
rect 32606 23968 32922 23969
rect 32606 23904 32612 23968
rect 32676 23904 32692 23968
rect 32756 23904 32772 23968
rect 32836 23904 32852 23968
rect 32916 23904 32922 23968
rect 32606 23903 32922 23904
rect 37606 23968 37922 23969
rect 37606 23904 37612 23968
rect 37676 23904 37692 23968
rect 37756 23904 37772 23968
rect 37836 23904 37852 23968
rect 37916 23904 37922 23968
rect 37606 23903 37922 23904
rect 1946 23424 2262 23425
rect 1946 23360 1952 23424
rect 2016 23360 2032 23424
rect 2096 23360 2112 23424
rect 2176 23360 2192 23424
rect 2256 23360 2262 23424
rect 1946 23359 2262 23360
rect 6946 23424 7262 23425
rect 6946 23360 6952 23424
rect 7016 23360 7032 23424
rect 7096 23360 7112 23424
rect 7176 23360 7192 23424
rect 7256 23360 7262 23424
rect 6946 23359 7262 23360
rect 11946 23424 12262 23425
rect 11946 23360 11952 23424
rect 12016 23360 12032 23424
rect 12096 23360 12112 23424
rect 12176 23360 12192 23424
rect 12256 23360 12262 23424
rect 11946 23359 12262 23360
rect 16946 23424 17262 23425
rect 16946 23360 16952 23424
rect 17016 23360 17032 23424
rect 17096 23360 17112 23424
rect 17176 23360 17192 23424
rect 17256 23360 17262 23424
rect 16946 23359 17262 23360
rect 21946 23424 22262 23425
rect 21946 23360 21952 23424
rect 22016 23360 22032 23424
rect 22096 23360 22112 23424
rect 22176 23360 22192 23424
rect 22256 23360 22262 23424
rect 21946 23359 22262 23360
rect 26946 23424 27262 23425
rect 26946 23360 26952 23424
rect 27016 23360 27032 23424
rect 27096 23360 27112 23424
rect 27176 23360 27192 23424
rect 27256 23360 27262 23424
rect 26946 23359 27262 23360
rect 31946 23424 32262 23425
rect 31946 23360 31952 23424
rect 32016 23360 32032 23424
rect 32096 23360 32112 23424
rect 32176 23360 32192 23424
rect 32256 23360 32262 23424
rect 31946 23359 32262 23360
rect 36946 23424 37262 23425
rect 36946 23360 36952 23424
rect 37016 23360 37032 23424
rect 37096 23360 37112 23424
rect 37176 23360 37192 23424
rect 37256 23360 37262 23424
rect 36946 23359 37262 23360
rect 2606 22880 2922 22881
rect 2606 22816 2612 22880
rect 2676 22816 2692 22880
rect 2756 22816 2772 22880
rect 2836 22816 2852 22880
rect 2916 22816 2922 22880
rect 2606 22815 2922 22816
rect 7606 22880 7922 22881
rect 7606 22816 7612 22880
rect 7676 22816 7692 22880
rect 7756 22816 7772 22880
rect 7836 22816 7852 22880
rect 7916 22816 7922 22880
rect 7606 22815 7922 22816
rect 12606 22880 12922 22881
rect 12606 22816 12612 22880
rect 12676 22816 12692 22880
rect 12756 22816 12772 22880
rect 12836 22816 12852 22880
rect 12916 22816 12922 22880
rect 12606 22815 12922 22816
rect 17606 22880 17922 22881
rect 17606 22816 17612 22880
rect 17676 22816 17692 22880
rect 17756 22816 17772 22880
rect 17836 22816 17852 22880
rect 17916 22816 17922 22880
rect 17606 22815 17922 22816
rect 22606 22880 22922 22881
rect 22606 22816 22612 22880
rect 22676 22816 22692 22880
rect 22756 22816 22772 22880
rect 22836 22816 22852 22880
rect 22916 22816 22922 22880
rect 22606 22815 22922 22816
rect 27606 22880 27922 22881
rect 27606 22816 27612 22880
rect 27676 22816 27692 22880
rect 27756 22816 27772 22880
rect 27836 22816 27852 22880
rect 27916 22816 27922 22880
rect 27606 22815 27922 22816
rect 32606 22880 32922 22881
rect 32606 22816 32612 22880
rect 32676 22816 32692 22880
rect 32756 22816 32772 22880
rect 32836 22816 32852 22880
rect 32916 22816 32922 22880
rect 32606 22815 32922 22816
rect 37606 22880 37922 22881
rect 37606 22816 37612 22880
rect 37676 22816 37692 22880
rect 37756 22816 37772 22880
rect 37836 22816 37852 22880
rect 37916 22816 37922 22880
rect 37606 22815 37922 22816
rect 3233 22674 3299 22677
rect 6913 22674 6979 22677
rect 3233 22672 6979 22674
rect 3233 22616 3238 22672
rect 3294 22616 6918 22672
rect 6974 22616 6979 22672
rect 3233 22614 6979 22616
rect 3233 22611 3299 22614
rect 6913 22611 6979 22614
rect 21030 22612 21036 22676
rect 21100 22674 21106 22676
rect 24577 22674 24643 22677
rect 21100 22672 24643 22674
rect 21100 22616 24582 22672
rect 24638 22616 24643 22672
rect 21100 22614 24643 22616
rect 21100 22612 21106 22614
rect 24577 22611 24643 22614
rect 1946 22336 2262 22337
rect 1946 22272 1952 22336
rect 2016 22272 2032 22336
rect 2096 22272 2112 22336
rect 2176 22272 2192 22336
rect 2256 22272 2262 22336
rect 1946 22271 2262 22272
rect 6946 22336 7262 22337
rect 6946 22272 6952 22336
rect 7016 22272 7032 22336
rect 7096 22272 7112 22336
rect 7176 22272 7192 22336
rect 7256 22272 7262 22336
rect 6946 22271 7262 22272
rect 11946 22336 12262 22337
rect 11946 22272 11952 22336
rect 12016 22272 12032 22336
rect 12096 22272 12112 22336
rect 12176 22272 12192 22336
rect 12256 22272 12262 22336
rect 11946 22271 12262 22272
rect 16946 22336 17262 22337
rect 16946 22272 16952 22336
rect 17016 22272 17032 22336
rect 17096 22272 17112 22336
rect 17176 22272 17192 22336
rect 17256 22272 17262 22336
rect 16946 22271 17262 22272
rect 21946 22336 22262 22337
rect 21946 22272 21952 22336
rect 22016 22272 22032 22336
rect 22096 22272 22112 22336
rect 22176 22272 22192 22336
rect 22256 22272 22262 22336
rect 21946 22271 22262 22272
rect 26946 22336 27262 22337
rect 26946 22272 26952 22336
rect 27016 22272 27032 22336
rect 27096 22272 27112 22336
rect 27176 22272 27192 22336
rect 27256 22272 27262 22336
rect 26946 22271 27262 22272
rect 31946 22336 32262 22337
rect 31946 22272 31952 22336
rect 32016 22272 32032 22336
rect 32096 22272 32112 22336
rect 32176 22272 32192 22336
rect 32256 22272 32262 22336
rect 31946 22271 32262 22272
rect 36946 22336 37262 22337
rect 36946 22272 36952 22336
rect 37016 22272 37032 22336
rect 37096 22272 37112 22336
rect 37176 22272 37192 22336
rect 37256 22272 37262 22336
rect 36946 22271 37262 22272
rect 11053 21994 11119 21997
rect 21030 21994 21036 21996
rect 11053 21992 21036 21994
rect 11053 21936 11058 21992
rect 11114 21936 21036 21992
rect 11053 21934 21036 21936
rect 11053 21931 11119 21934
rect 21030 21932 21036 21934
rect 21100 21932 21106 21996
rect 2606 21792 2922 21793
rect 2606 21728 2612 21792
rect 2676 21728 2692 21792
rect 2756 21728 2772 21792
rect 2836 21728 2852 21792
rect 2916 21728 2922 21792
rect 2606 21727 2922 21728
rect 7606 21792 7922 21793
rect 7606 21728 7612 21792
rect 7676 21728 7692 21792
rect 7756 21728 7772 21792
rect 7836 21728 7852 21792
rect 7916 21728 7922 21792
rect 7606 21727 7922 21728
rect 12606 21792 12922 21793
rect 12606 21728 12612 21792
rect 12676 21728 12692 21792
rect 12756 21728 12772 21792
rect 12836 21728 12852 21792
rect 12916 21728 12922 21792
rect 12606 21727 12922 21728
rect 17606 21792 17922 21793
rect 17606 21728 17612 21792
rect 17676 21728 17692 21792
rect 17756 21728 17772 21792
rect 17836 21728 17852 21792
rect 17916 21728 17922 21792
rect 17606 21727 17922 21728
rect 22606 21792 22922 21793
rect 22606 21728 22612 21792
rect 22676 21728 22692 21792
rect 22756 21728 22772 21792
rect 22836 21728 22852 21792
rect 22916 21728 22922 21792
rect 22606 21727 22922 21728
rect 27606 21792 27922 21793
rect 27606 21728 27612 21792
rect 27676 21728 27692 21792
rect 27756 21728 27772 21792
rect 27836 21728 27852 21792
rect 27916 21728 27922 21792
rect 27606 21727 27922 21728
rect 32606 21792 32922 21793
rect 32606 21728 32612 21792
rect 32676 21728 32692 21792
rect 32756 21728 32772 21792
rect 32836 21728 32852 21792
rect 32916 21728 32922 21792
rect 32606 21727 32922 21728
rect 37606 21792 37922 21793
rect 37606 21728 37612 21792
rect 37676 21728 37692 21792
rect 37756 21728 37772 21792
rect 37836 21728 37852 21792
rect 37916 21728 37922 21792
rect 37606 21727 37922 21728
rect 1946 21248 2262 21249
rect 1946 21184 1952 21248
rect 2016 21184 2032 21248
rect 2096 21184 2112 21248
rect 2176 21184 2192 21248
rect 2256 21184 2262 21248
rect 1946 21183 2262 21184
rect 6946 21248 7262 21249
rect 6946 21184 6952 21248
rect 7016 21184 7032 21248
rect 7096 21184 7112 21248
rect 7176 21184 7192 21248
rect 7256 21184 7262 21248
rect 6946 21183 7262 21184
rect 11946 21248 12262 21249
rect 11946 21184 11952 21248
rect 12016 21184 12032 21248
rect 12096 21184 12112 21248
rect 12176 21184 12192 21248
rect 12256 21184 12262 21248
rect 11946 21183 12262 21184
rect 16946 21248 17262 21249
rect 16946 21184 16952 21248
rect 17016 21184 17032 21248
rect 17096 21184 17112 21248
rect 17176 21184 17192 21248
rect 17256 21184 17262 21248
rect 16946 21183 17262 21184
rect 21946 21248 22262 21249
rect 21946 21184 21952 21248
rect 22016 21184 22032 21248
rect 22096 21184 22112 21248
rect 22176 21184 22192 21248
rect 22256 21184 22262 21248
rect 21946 21183 22262 21184
rect 26946 21248 27262 21249
rect 26946 21184 26952 21248
rect 27016 21184 27032 21248
rect 27096 21184 27112 21248
rect 27176 21184 27192 21248
rect 27256 21184 27262 21248
rect 26946 21183 27262 21184
rect 31946 21248 32262 21249
rect 31946 21184 31952 21248
rect 32016 21184 32032 21248
rect 32096 21184 32112 21248
rect 32176 21184 32192 21248
rect 32256 21184 32262 21248
rect 31946 21183 32262 21184
rect 36946 21248 37262 21249
rect 36946 21184 36952 21248
rect 37016 21184 37032 21248
rect 37096 21184 37112 21248
rect 37176 21184 37192 21248
rect 37256 21184 37262 21248
rect 36946 21183 37262 21184
rect 2606 20704 2922 20705
rect 2606 20640 2612 20704
rect 2676 20640 2692 20704
rect 2756 20640 2772 20704
rect 2836 20640 2852 20704
rect 2916 20640 2922 20704
rect 2606 20639 2922 20640
rect 7606 20704 7922 20705
rect 7606 20640 7612 20704
rect 7676 20640 7692 20704
rect 7756 20640 7772 20704
rect 7836 20640 7852 20704
rect 7916 20640 7922 20704
rect 7606 20639 7922 20640
rect 12606 20704 12922 20705
rect 12606 20640 12612 20704
rect 12676 20640 12692 20704
rect 12756 20640 12772 20704
rect 12836 20640 12852 20704
rect 12916 20640 12922 20704
rect 12606 20639 12922 20640
rect 17606 20704 17922 20705
rect 17606 20640 17612 20704
rect 17676 20640 17692 20704
rect 17756 20640 17772 20704
rect 17836 20640 17852 20704
rect 17916 20640 17922 20704
rect 17606 20639 17922 20640
rect 22606 20704 22922 20705
rect 22606 20640 22612 20704
rect 22676 20640 22692 20704
rect 22756 20640 22772 20704
rect 22836 20640 22852 20704
rect 22916 20640 22922 20704
rect 22606 20639 22922 20640
rect 27606 20704 27922 20705
rect 27606 20640 27612 20704
rect 27676 20640 27692 20704
rect 27756 20640 27772 20704
rect 27836 20640 27852 20704
rect 27916 20640 27922 20704
rect 27606 20639 27922 20640
rect 32606 20704 32922 20705
rect 32606 20640 32612 20704
rect 32676 20640 32692 20704
rect 32756 20640 32772 20704
rect 32836 20640 32852 20704
rect 32916 20640 32922 20704
rect 32606 20639 32922 20640
rect 37606 20704 37922 20705
rect 37606 20640 37612 20704
rect 37676 20640 37692 20704
rect 37756 20640 37772 20704
rect 37836 20640 37852 20704
rect 37916 20640 37922 20704
rect 37606 20639 37922 20640
rect 1946 20160 2262 20161
rect 1946 20096 1952 20160
rect 2016 20096 2032 20160
rect 2096 20096 2112 20160
rect 2176 20096 2192 20160
rect 2256 20096 2262 20160
rect 1946 20095 2262 20096
rect 6946 20160 7262 20161
rect 6946 20096 6952 20160
rect 7016 20096 7032 20160
rect 7096 20096 7112 20160
rect 7176 20096 7192 20160
rect 7256 20096 7262 20160
rect 6946 20095 7262 20096
rect 11946 20160 12262 20161
rect 11946 20096 11952 20160
rect 12016 20096 12032 20160
rect 12096 20096 12112 20160
rect 12176 20096 12192 20160
rect 12256 20096 12262 20160
rect 11946 20095 12262 20096
rect 16946 20160 17262 20161
rect 16946 20096 16952 20160
rect 17016 20096 17032 20160
rect 17096 20096 17112 20160
rect 17176 20096 17192 20160
rect 17256 20096 17262 20160
rect 16946 20095 17262 20096
rect 21946 20160 22262 20161
rect 21946 20096 21952 20160
rect 22016 20096 22032 20160
rect 22096 20096 22112 20160
rect 22176 20096 22192 20160
rect 22256 20096 22262 20160
rect 21946 20095 22262 20096
rect 26946 20160 27262 20161
rect 26946 20096 26952 20160
rect 27016 20096 27032 20160
rect 27096 20096 27112 20160
rect 27176 20096 27192 20160
rect 27256 20096 27262 20160
rect 26946 20095 27262 20096
rect 31946 20160 32262 20161
rect 31946 20096 31952 20160
rect 32016 20096 32032 20160
rect 32096 20096 32112 20160
rect 32176 20096 32192 20160
rect 32256 20096 32262 20160
rect 31946 20095 32262 20096
rect 36946 20160 37262 20161
rect 36946 20096 36952 20160
rect 37016 20096 37032 20160
rect 37096 20096 37112 20160
rect 37176 20096 37192 20160
rect 37256 20096 37262 20160
rect 36946 20095 37262 20096
rect 2606 19616 2922 19617
rect 2606 19552 2612 19616
rect 2676 19552 2692 19616
rect 2756 19552 2772 19616
rect 2836 19552 2852 19616
rect 2916 19552 2922 19616
rect 2606 19551 2922 19552
rect 7606 19616 7922 19617
rect 7606 19552 7612 19616
rect 7676 19552 7692 19616
rect 7756 19552 7772 19616
rect 7836 19552 7852 19616
rect 7916 19552 7922 19616
rect 7606 19551 7922 19552
rect 12606 19616 12922 19617
rect 12606 19552 12612 19616
rect 12676 19552 12692 19616
rect 12756 19552 12772 19616
rect 12836 19552 12852 19616
rect 12916 19552 12922 19616
rect 12606 19551 12922 19552
rect 17606 19616 17922 19617
rect 17606 19552 17612 19616
rect 17676 19552 17692 19616
rect 17756 19552 17772 19616
rect 17836 19552 17852 19616
rect 17916 19552 17922 19616
rect 17606 19551 17922 19552
rect 22606 19616 22922 19617
rect 22606 19552 22612 19616
rect 22676 19552 22692 19616
rect 22756 19552 22772 19616
rect 22836 19552 22852 19616
rect 22916 19552 22922 19616
rect 22606 19551 22922 19552
rect 27606 19616 27922 19617
rect 27606 19552 27612 19616
rect 27676 19552 27692 19616
rect 27756 19552 27772 19616
rect 27836 19552 27852 19616
rect 27916 19552 27922 19616
rect 27606 19551 27922 19552
rect 32606 19616 32922 19617
rect 32606 19552 32612 19616
rect 32676 19552 32692 19616
rect 32756 19552 32772 19616
rect 32836 19552 32852 19616
rect 32916 19552 32922 19616
rect 32606 19551 32922 19552
rect 37606 19616 37922 19617
rect 37606 19552 37612 19616
rect 37676 19552 37692 19616
rect 37756 19552 37772 19616
rect 37836 19552 37852 19616
rect 37916 19552 37922 19616
rect 37606 19551 37922 19552
rect 1946 19072 2262 19073
rect 1946 19008 1952 19072
rect 2016 19008 2032 19072
rect 2096 19008 2112 19072
rect 2176 19008 2192 19072
rect 2256 19008 2262 19072
rect 1946 19007 2262 19008
rect 6946 19072 7262 19073
rect 6946 19008 6952 19072
rect 7016 19008 7032 19072
rect 7096 19008 7112 19072
rect 7176 19008 7192 19072
rect 7256 19008 7262 19072
rect 6946 19007 7262 19008
rect 11946 19072 12262 19073
rect 11946 19008 11952 19072
rect 12016 19008 12032 19072
rect 12096 19008 12112 19072
rect 12176 19008 12192 19072
rect 12256 19008 12262 19072
rect 11946 19007 12262 19008
rect 16946 19072 17262 19073
rect 16946 19008 16952 19072
rect 17016 19008 17032 19072
rect 17096 19008 17112 19072
rect 17176 19008 17192 19072
rect 17256 19008 17262 19072
rect 16946 19007 17262 19008
rect 21946 19072 22262 19073
rect 21946 19008 21952 19072
rect 22016 19008 22032 19072
rect 22096 19008 22112 19072
rect 22176 19008 22192 19072
rect 22256 19008 22262 19072
rect 21946 19007 22262 19008
rect 26946 19072 27262 19073
rect 26946 19008 26952 19072
rect 27016 19008 27032 19072
rect 27096 19008 27112 19072
rect 27176 19008 27192 19072
rect 27256 19008 27262 19072
rect 26946 19007 27262 19008
rect 31946 19072 32262 19073
rect 31946 19008 31952 19072
rect 32016 19008 32032 19072
rect 32096 19008 32112 19072
rect 32176 19008 32192 19072
rect 32256 19008 32262 19072
rect 31946 19007 32262 19008
rect 36946 19072 37262 19073
rect 36946 19008 36952 19072
rect 37016 19008 37032 19072
rect 37096 19008 37112 19072
rect 37176 19008 37192 19072
rect 37256 19008 37262 19072
rect 36946 19007 37262 19008
rect 2606 18528 2922 18529
rect 2606 18464 2612 18528
rect 2676 18464 2692 18528
rect 2756 18464 2772 18528
rect 2836 18464 2852 18528
rect 2916 18464 2922 18528
rect 2606 18463 2922 18464
rect 7606 18528 7922 18529
rect 7606 18464 7612 18528
rect 7676 18464 7692 18528
rect 7756 18464 7772 18528
rect 7836 18464 7852 18528
rect 7916 18464 7922 18528
rect 7606 18463 7922 18464
rect 12606 18528 12922 18529
rect 12606 18464 12612 18528
rect 12676 18464 12692 18528
rect 12756 18464 12772 18528
rect 12836 18464 12852 18528
rect 12916 18464 12922 18528
rect 12606 18463 12922 18464
rect 17606 18528 17922 18529
rect 17606 18464 17612 18528
rect 17676 18464 17692 18528
rect 17756 18464 17772 18528
rect 17836 18464 17852 18528
rect 17916 18464 17922 18528
rect 17606 18463 17922 18464
rect 22606 18528 22922 18529
rect 22606 18464 22612 18528
rect 22676 18464 22692 18528
rect 22756 18464 22772 18528
rect 22836 18464 22852 18528
rect 22916 18464 22922 18528
rect 22606 18463 22922 18464
rect 27606 18528 27922 18529
rect 27606 18464 27612 18528
rect 27676 18464 27692 18528
rect 27756 18464 27772 18528
rect 27836 18464 27852 18528
rect 27916 18464 27922 18528
rect 27606 18463 27922 18464
rect 32606 18528 32922 18529
rect 32606 18464 32612 18528
rect 32676 18464 32692 18528
rect 32756 18464 32772 18528
rect 32836 18464 32852 18528
rect 32916 18464 32922 18528
rect 32606 18463 32922 18464
rect 37606 18528 37922 18529
rect 37606 18464 37612 18528
rect 37676 18464 37692 18528
rect 37756 18464 37772 18528
rect 37836 18464 37852 18528
rect 37916 18464 37922 18528
rect 37606 18463 37922 18464
rect 1946 17984 2262 17985
rect 1946 17920 1952 17984
rect 2016 17920 2032 17984
rect 2096 17920 2112 17984
rect 2176 17920 2192 17984
rect 2256 17920 2262 17984
rect 1946 17919 2262 17920
rect 6946 17984 7262 17985
rect 6946 17920 6952 17984
rect 7016 17920 7032 17984
rect 7096 17920 7112 17984
rect 7176 17920 7192 17984
rect 7256 17920 7262 17984
rect 6946 17919 7262 17920
rect 11946 17984 12262 17985
rect 11946 17920 11952 17984
rect 12016 17920 12032 17984
rect 12096 17920 12112 17984
rect 12176 17920 12192 17984
rect 12256 17920 12262 17984
rect 11946 17919 12262 17920
rect 16946 17984 17262 17985
rect 16946 17920 16952 17984
rect 17016 17920 17032 17984
rect 17096 17920 17112 17984
rect 17176 17920 17192 17984
rect 17256 17920 17262 17984
rect 16946 17919 17262 17920
rect 21946 17984 22262 17985
rect 21946 17920 21952 17984
rect 22016 17920 22032 17984
rect 22096 17920 22112 17984
rect 22176 17920 22192 17984
rect 22256 17920 22262 17984
rect 21946 17919 22262 17920
rect 26946 17984 27262 17985
rect 26946 17920 26952 17984
rect 27016 17920 27032 17984
rect 27096 17920 27112 17984
rect 27176 17920 27192 17984
rect 27256 17920 27262 17984
rect 26946 17919 27262 17920
rect 31946 17984 32262 17985
rect 31946 17920 31952 17984
rect 32016 17920 32032 17984
rect 32096 17920 32112 17984
rect 32176 17920 32192 17984
rect 32256 17920 32262 17984
rect 31946 17919 32262 17920
rect 36946 17984 37262 17985
rect 36946 17920 36952 17984
rect 37016 17920 37032 17984
rect 37096 17920 37112 17984
rect 37176 17920 37192 17984
rect 37256 17920 37262 17984
rect 36946 17919 37262 17920
rect 2606 17440 2922 17441
rect 2606 17376 2612 17440
rect 2676 17376 2692 17440
rect 2756 17376 2772 17440
rect 2836 17376 2852 17440
rect 2916 17376 2922 17440
rect 2606 17375 2922 17376
rect 7606 17440 7922 17441
rect 7606 17376 7612 17440
rect 7676 17376 7692 17440
rect 7756 17376 7772 17440
rect 7836 17376 7852 17440
rect 7916 17376 7922 17440
rect 7606 17375 7922 17376
rect 12606 17440 12922 17441
rect 12606 17376 12612 17440
rect 12676 17376 12692 17440
rect 12756 17376 12772 17440
rect 12836 17376 12852 17440
rect 12916 17376 12922 17440
rect 12606 17375 12922 17376
rect 17606 17440 17922 17441
rect 17606 17376 17612 17440
rect 17676 17376 17692 17440
rect 17756 17376 17772 17440
rect 17836 17376 17852 17440
rect 17916 17376 17922 17440
rect 17606 17375 17922 17376
rect 22606 17440 22922 17441
rect 22606 17376 22612 17440
rect 22676 17376 22692 17440
rect 22756 17376 22772 17440
rect 22836 17376 22852 17440
rect 22916 17376 22922 17440
rect 22606 17375 22922 17376
rect 27606 17440 27922 17441
rect 27606 17376 27612 17440
rect 27676 17376 27692 17440
rect 27756 17376 27772 17440
rect 27836 17376 27852 17440
rect 27916 17376 27922 17440
rect 27606 17375 27922 17376
rect 32606 17440 32922 17441
rect 32606 17376 32612 17440
rect 32676 17376 32692 17440
rect 32756 17376 32772 17440
rect 32836 17376 32852 17440
rect 32916 17376 32922 17440
rect 32606 17375 32922 17376
rect 37606 17440 37922 17441
rect 37606 17376 37612 17440
rect 37676 17376 37692 17440
rect 37756 17376 37772 17440
rect 37836 17376 37852 17440
rect 37916 17376 37922 17440
rect 37606 17375 37922 17376
rect 1946 16896 2262 16897
rect 1946 16832 1952 16896
rect 2016 16832 2032 16896
rect 2096 16832 2112 16896
rect 2176 16832 2192 16896
rect 2256 16832 2262 16896
rect 1946 16831 2262 16832
rect 6946 16896 7262 16897
rect 6946 16832 6952 16896
rect 7016 16832 7032 16896
rect 7096 16832 7112 16896
rect 7176 16832 7192 16896
rect 7256 16832 7262 16896
rect 6946 16831 7262 16832
rect 11946 16896 12262 16897
rect 11946 16832 11952 16896
rect 12016 16832 12032 16896
rect 12096 16832 12112 16896
rect 12176 16832 12192 16896
rect 12256 16832 12262 16896
rect 11946 16831 12262 16832
rect 16946 16896 17262 16897
rect 16946 16832 16952 16896
rect 17016 16832 17032 16896
rect 17096 16832 17112 16896
rect 17176 16832 17192 16896
rect 17256 16832 17262 16896
rect 16946 16831 17262 16832
rect 21946 16896 22262 16897
rect 21946 16832 21952 16896
rect 22016 16832 22032 16896
rect 22096 16832 22112 16896
rect 22176 16832 22192 16896
rect 22256 16832 22262 16896
rect 21946 16831 22262 16832
rect 26946 16896 27262 16897
rect 26946 16832 26952 16896
rect 27016 16832 27032 16896
rect 27096 16832 27112 16896
rect 27176 16832 27192 16896
rect 27256 16832 27262 16896
rect 26946 16831 27262 16832
rect 31946 16896 32262 16897
rect 31946 16832 31952 16896
rect 32016 16832 32032 16896
rect 32096 16832 32112 16896
rect 32176 16832 32192 16896
rect 32256 16832 32262 16896
rect 31946 16831 32262 16832
rect 36946 16896 37262 16897
rect 36946 16832 36952 16896
rect 37016 16832 37032 16896
rect 37096 16832 37112 16896
rect 37176 16832 37192 16896
rect 37256 16832 37262 16896
rect 36946 16831 37262 16832
rect 2606 16352 2922 16353
rect 2606 16288 2612 16352
rect 2676 16288 2692 16352
rect 2756 16288 2772 16352
rect 2836 16288 2852 16352
rect 2916 16288 2922 16352
rect 2606 16287 2922 16288
rect 7606 16352 7922 16353
rect 7606 16288 7612 16352
rect 7676 16288 7692 16352
rect 7756 16288 7772 16352
rect 7836 16288 7852 16352
rect 7916 16288 7922 16352
rect 7606 16287 7922 16288
rect 12606 16352 12922 16353
rect 12606 16288 12612 16352
rect 12676 16288 12692 16352
rect 12756 16288 12772 16352
rect 12836 16288 12852 16352
rect 12916 16288 12922 16352
rect 12606 16287 12922 16288
rect 17606 16352 17922 16353
rect 17606 16288 17612 16352
rect 17676 16288 17692 16352
rect 17756 16288 17772 16352
rect 17836 16288 17852 16352
rect 17916 16288 17922 16352
rect 17606 16287 17922 16288
rect 22606 16352 22922 16353
rect 22606 16288 22612 16352
rect 22676 16288 22692 16352
rect 22756 16288 22772 16352
rect 22836 16288 22852 16352
rect 22916 16288 22922 16352
rect 22606 16287 22922 16288
rect 27606 16352 27922 16353
rect 27606 16288 27612 16352
rect 27676 16288 27692 16352
rect 27756 16288 27772 16352
rect 27836 16288 27852 16352
rect 27916 16288 27922 16352
rect 27606 16287 27922 16288
rect 32606 16352 32922 16353
rect 32606 16288 32612 16352
rect 32676 16288 32692 16352
rect 32756 16288 32772 16352
rect 32836 16288 32852 16352
rect 32916 16288 32922 16352
rect 32606 16287 32922 16288
rect 37606 16352 37922 16353
rect 37606 16288 37612 16352
rect 37676 16288 37692 16352
rect 37756 16288 37772 16352
rect 37836 16288 37852 16352
rect 37916 16288 37922 16352
rect 37606 16287 37922 16288
rect 1946 15808 2262 15809
rect 1946 15744 1952 15808
rect 2016 15744 2032 15808
rect 2096 15744 2112 15808
rect 2176 15744 2192 15808
rect 2256 15744 2262 15808
rect 1946 15743 2262 15744
rect 6946 15808 7262 15809
rect 6946 15744 6952 15808
rect 7016 15744 7032 15808
rect 7096 15744 7112 15808
rect 7176 15744 7192 15808
rect 7256 15744 7262 15808
rect 6946 15743 7262 15744
rect 11946 15808 12262 15809
rect 11946 15744 11952 15808
rect 12016 15744 12032 15808
rect 12096 15744 12112 15808
rect 12176 15744 12192 15808
rect 12256 15744 12262 15808
rect 11946 15743 12262 15744
rect 16946 15808 17262 15809
rect 16946 15744 16952 15808
rect 17016 15744 17032 15808
rect 17096 15744 17112 15808
rect 17176 15744 17192 15808
rect 17256 15744 17262 15808
rect 16946 15743 17262 15744
rect 21946 15808 22262 15809
rect 21946 15744 21952 15808
rect 22016 15744 22032 15808
rect 22096 15744 22112 15808
rect 22176 15744 22192 15808
rect 22256 15744 22262 15808
rect 21946 15743 22262 15744
rect 26946 15808 27262 15809
rect 26946 15744 26952 15808
rect 27016 15744 27032 15808
rect 27096 15744 27112 15808
rect 27176 15744 27192 15808
rect 27256 15744 27262 15808
rect 26946 15743 27262 15744
rect 31946 15808 32262 15809
rect 31946 15744 31952 15808
rect 32016 15744 32032 15808
rect 32096 15744 32112 15808
rect 32176 15744 32192 15808
rect 32256 15744 32262 15808
rect 31946 15743 32262 15744
rect 36946 15808 37262 15809
rect 36946 15744 36952 15808
rect 37016 15744 37032 15808
rect 37096 15744 37112 15808
rect 37176 15744 37192 15808
rect 37256 15744 37262 15808
rect 36946 15743 37262 15744
rect 2606 15264 2922 15265
rect 2606 15200 2612 15264
rect 2676 15200 2692 15264
rect 2756 15200 2772 15264
rect 2836 15200 2852 15264
rect 2916 15200 2922 15264
rect 2606 15199 2922 15200
rect 7606 15264 7922 15265
rect 7606 15200 7612 15264
rect 7676 15200 7692 15264
rect 7756 15200 7772 15264
rect 7836 15200 7852 15264
rect 7916 15200 7922 15264
rect 7606 15199 7922 15200
rect 12606 15264 12922 15265
rect 12606 15200 12612 15264
rect 12676 15200 12692 15264
rect 12756 15200 12772 15264
rect 12836 15200 12852 15264
rect 12916 15200 12922 15264
rect 12606 15199 12922 15200
rect 17606 15264 17922 15265
rect 17606 15200 17612 15264
rect 17676 15200 17692 15264
rect 17756 15200 17772 15264
rect 17836 15200 17852 15264
rect 17916 15200 17922 15264
rect 17606 15199 17922 15200
rect 22606 15264 22922 15265
rect 22606 15200 22612 15264
rect 22676 15200 22692 15264
rect 22756 15200 22772 15264
rect 22836 15200 22852 15264
rect 22916 15200 22922 15264
rect 22606 15199 22922 15200
rect 27606 15264 27922 15265
rect 27606 15200 27612 15264
rect 27676 15200 27692 15264
rect 27756 15200 27772 15264
rect 27836 15200 27852 15264
rect 27916 15200 27922 15264
rect 27606 15199 27922 15200
rect 32606 15264 32922 15265
rect 32606 15200 32612 15264
rect 32676 15200 32692 15264
rect 32756 15200 32772 15264
rect 32836 15200 32852 15264
rect 32916 15200 32922 15264
rect 32606 15199 32922 15200
rect 37606 15264 37922 15265
rect 37606 15200 37612 15264
rect 37676 15200 37692 15264
rect 37756 15200 37772 15264
rect 37836 15200 37852 15264
rect 37916 15200 37922 15264
rect 37606 15199 37922 15200
rect 1946 14720 2262 14721
rect 1946 14656 1952 14720
rect 2016 14656 2032 14720
rect 2096 14656 2112 14720
rect 2176 14656 2192 14720
rect 2256 14656 2262 14720
rect 1946 14655 2262 14656
rect 6946 14720 7262 14721
rect 6946 14656 6952 14720
rect 7016 14656 7032 14720
rect 7096 14656 7112 14720
rect 7176 14656 7192 14720
rect 7256 14656 7262 14720
rect 6946 14655 7262 14656
rect 11946 14720 12262 14721
rect 11946 14656 11952 14720
rect 12016 14656 12032 14720
rect 12096 14656 12112 14720
rect 12176 14656 12192 14720
rect 12256 14656 12262 14720
rect 11946 14655 12262 14656
rect 16946 14720 17262 14721
rect 16946 14656 16952 14720
rect 17016 14656 17032 14720
rect 17096 14656 17112 14720
rect 17176 14656 17192 14720
rect 17256 14656 17262 14720
rect 16946 14655 17262 14656
rect 21946 14720 22262 14721
rect 21946 14656 21952 14720
rect 22016 14656 22032 14720
rect 22096 14656 22112 14720
rect 22176 14656 22192 14720
rect 22256 14656 22262 14720
rect 21946 14655 22262 14656
rect 26946 14720 27262 14721
rect 26946 14656 26952 14720
rect 27016 14656 27032 14720
rect 27096 14656 27112 14720
rect 27176 14656 27192 14720
rect 27256 14656 27262 14720
rect 26946 14655 27262 14656
rect 31946 14720 32262 14721
rect 31946 14656 31952 14720
rect 32016 14656 32032 14720
rect 32096 14656 32112 14720
rect 32176 14656 32192 14720
rect 32256 14656 32262 14720
rect 31946 14655 32262 14656
rect 36946 14720 37262 14721
rect 36946 14656 36952 14720
rect 37016 14656 37032 14720
rect 37096 14656 37112 14720
rect 37176 14656 37192 14720
rect 37256 14656 37262 14720
rect 36946 14655 37262 14656
rect 33910 14316 33916 14380
rect 33980 14378 33986 14380
rect 38929 14378 38995 14381
rect 33980 14376 38995 14378
rect 33980 14320 38934 14376
rect 38990 14320 38995 14376
rect 33980 14318 38995 14320
rect 33980 14316 33986 14318
rect 38929 14315 38995 14318
rect 2606 14176 2922 14177
rect 2606 14112 2612 14176
rect 2676 14112 2692 14176
rect 2756 14112 2772 14176
rect 2836 14112 2852 14176
rect 2916 14112 2922 14176
rect 2606 14111 2922 14112
rect 7606 14176 7922 14177
rect 7606 14112 7612 14176
rect 7676 14112 7692 14176
rect 7756 14112 7772 14176
rect 7836 14112 7852 14176
rect 7916 14112 7922 14176
rect 7606 14111 7922 14112
rect 12606 14176 12922 14177
rect 12606 14112 12612 14176
rect 12676 14112 12692 14176
rect 12756 14112 12772 14176
rect 12836 14112 12852 14176
rect 12916 14112 12922 14176
rect 12606 14111 12922 14112
rect 17606 14176 17922 14177
rect 17606 14112 17612 14176
rect 17676 14112 17692 14176
rect 17756 14112 17772 14176
rect 17836 14112 17852 14176
rect 17916 14112 17922 14176
rect 17606 14111 17922 14112
rect 22606 14176 22922 14177
rect 22606 14112 22612 14176
rect 22676 14112 22692 14176
rect 22756 14112 22772 14176
rect 22836 14112 22852 14176
rect 22916 14112 22922 14176
rect 22606 14111 22922 14112
rect 27606 14176 27922 14177
rect 27606 14112 27612 14176
rect 27676 14112 27692 14176
rect 27756 14112 27772 14176
rect 27836 14112 27852 14176
rect 27916 14112 27922 14176
rect 27606 14111 27922 14112
rect 32606 14176 32922 14177
rect 32606 14112 32612 14176
rect 32676 14112 32692 14176
rect 32756 14112 32772 14176
rect 32836 14112 32852 14176
rect 32916 14112 32922 14176
rect 32606 14111 32922 14112
rect 37606 14176 37922 14177
rect 37606 14112 37612 14176
rect 37676 14112 37692 14176
rect 37756 14112 37772 14176
rect 37836 14112 37852 14176
rect 37916 14112 37922 14176
rect 37606 14111 37922 14112
rect 1946 13632 2262 13633
rect 1946 13568 1952 13632
rect 2016 13568 2032 13632
rect 2096 13568 2112 13632
rect 2176 13568 2192 13632
rect 2256 13568 2262 13632
rect 1946 13567 2262 13568
rect 6946 13632 7262 13633
rect 6946 13568 6952 13632
rect 7016 13568 7032 13632
rect 7096 13568 7112 13632
rect 7176 13568 7192 13632
rect 7256 13568 7262 13632
rect 6946 13567 7262 13568
rect 11946 13632 12262 13633
rect 11946 13568 11952 13632
rect 12016 13568 12032 13632
rect 12096 13568 12112 13632
rect 12176 13568 12192 13632
rect 12256 13568 12262 13632
rect 11946 13567 12262 13568
rect 16946 13632 17262 13633
rect 16946 13568 16952 13632
rect 17016 13568 17032 13632
rect 17096 13568 17112 13632
rect 17176 13568 17192 13632
rect 17256 13568 17262 13632
rect 16946 13567 17262 13568
rect 21946 13632 22262 13633
rect 21946 13568 21952 13632
rect 22016 13568 22032 13632
rect 22096 13568 22112 13632
rect 22176 13568 22192 13632
rect 22256 13568 22262 13632
rect 21946 13567 22262 13568
rect 26946 13632 27262 13633
rect 26946 13568 26952 13632
rect 27016 13568 27032 13632
rect 27096 13568 27112 13632
rect 27176 13568 27192 13632
rect 27256 13568 27262 13632
rect 26946 13567 27262 13568
rect 31946 13632 32262 13633
rect 31946 13568 31952 13632
rect 32016 13568 32032 13632
rect 32096 13568 32112 13632
rect 32176 13568 32192 13632
rect 32256 13568 32262 13632
rect 31946 13567 32262 13568
rect 36946 13632 37262 13633
rect 36946 13568 36952 13632
rect 37016 13568 37032 13632
rect 37096 13568 37112 13632
rect 37176 13568 37192 13632
rect 37256 13568 37262 13632
rect 36946 13567 37262 13568
rect 2606 13088 2922 13089
rect 2606 13024 2612 13088
rect 2676 13024 2692 13088
rect 2756 13024 2772 13088
rect 2836 13024 2852 13088
rect 2916 13024 2922 13088
rect 2606 13023 2922 13024
rect 7606 13088 7922 13089
rect 7606 13024 7612 13088
rect 7676 13024 7692 13088
rect 7756 13024 7772 13088
rect 7836 13024 7852 13088
rect 7916 13024 7922 13088
rect 7606 13023 7922 13024
rect 12606 13088 12922 13089
rect 12606 13024 12612 13088
rect 12676 13024 12692 13088
rect 12756 13024 12772 13088
rect 12836 13024 12852 13088
rect 12916 13024 12922 13088
rect 12606 13023 12922 13024
rect 17606 13088 17922 13089
rect 17606 13024 17612 13088
rect 17676 13024 17692 13088
rect 17756 13024 17772 13088
rect 17836 13024 17852 13088
rect 17916 13024 17922 13088
rect 17606 13023 17922 13024
rect 22606 13088 22922 13089
rect 22606 13024 22612 13088
rect 22676 13024 22692 13088
rect 22756 13024 22772 13088
rect 22836 13024 22852 13088
rect 22916 13024 22922 13088
rect 22606 13023 22922 13024
rect 27606 13088 27922 13089
rect 27606 13024 27612 13088
rect 27676 13024 27692 13088
rect 27756 13024 27772 13088
rect 27836 13024 27852 13088
rect 27916 13024 27922 13088
rect 27606 13023 27922 13024
rect 32606 13088 32922 13089
rect 32606 13024 32612 13088
rect 32676 13024 32692 13088
rect 32756 13024 32772 13088
rect 32836 13024 32852 13088
rect 32916 13024 32922 13088
rect 32606 13023 32922 13024
rect 37606 13088 37922 13089
rect 37606 13024 37612 13088
rect 37676 13024 37692 13088
rect 37756 13024 37772 13088
rect 37836 13024 37852 13088
rect 37916 13024 37922 13088
rect 37606 13023 37922 13024
rect 1946 12544 2262 12545
rect 1946 12480 1952 12544
rect 2016 12480 2032 12544
rect 2096 12480 2112 12544
rect 2176 12480 2192 12544
rect 2256 12480 2262 12544
rect 1946 12479 2262 12480
rect 6946 12544 7262 12545
rect 6946 12480 6952 12544
rect 7016 12480 7032 12544
rect 7096 12480 7112 12544
rect 7176 12480 7192 12544
rect 7256 12480 7262 12544
rect 6946 12479 7262 12480
rect 11946 12544 12262 12545
rect 11946 12480 11952 12544
rect 12016 12480 12032 12544
rect 12096 12480 12112 12544
rect 12176 12480 12192 12544
rect 12256 12480 12262 12544
rect 11946 12479 12262 12480
rect 16946 12544 17262 12545
rect 16946 12480 16952 12544
rect 17016 12480 17032 12544
rect 17096 12480 17112 12544
rect 17176 12480 17192 12544
rect 17256 12480 17262 12544
rect 16946 12479 17262 12480
rect 21946 12544 22262 12545
rect 21946 12480 21952 12544
rect 22016 12480 22032 12544
rect 22096 12480 22112 12544
rect 22176 12480 22192 12544
rect 22256 12480 22262 12544
rect 21946 12479 22262 12480
rect 26946 12544 27262 12545
rect 26946 12480 26952 12544
rect 27016 12480 27032 12544
rect 27096 12480 27112 12544
rect 27176 12480 27192 12544
rect 27256 12480 27262 12544
rect 26946 12479 27262 12480
rect 31946 12544 32262 12545
rect 31946 12480 31952 12544
rect 32016 12480 32032 12544
rect 32096 12480 32112 12544
rect 32176 12480 32192 12544
rect 32256 12480 32262 12544
rect 31946 12479 32262 12480
rect 36946 12544 37262 12545
rect 36946 12480 36952 12544
rect 37016 12480 37032 12544
rect 37096 12480 37112 12544
rect 37176 12480 37192 12544
rect 37256 12480 37262 12544
rect 36946 12479 37262 12480
rect 2606 12000 2922 12001
rect 2606 11936 2612 12000
rect 2676 11936 2692 12000
rect 2756 11936 2772 12000
rect 2836 11936 2852 12000
rect 2916 11936 2922 12000
rect 2606 11935 2922 11936
rect 7606 12000 7922 12001
rect 7606 11936 7612 12000
rect 7676 11936 7692 12000
rect 7756 11936 7772 12000
rect 7836 11936 7852 12000
rect 7916 11936 7922 12000
rect 7606 11935 7922 11936
rect 12606 12000 12922 12001
rect 12606 11936 12612 12000
rect 12676 11936 12692 12000
rect 12756 11936 12772 12000
rect 12836 11936 12852 12000
rect 12916 11936 12922 12000
rect 12606 11935 12922 11936
rect 17606 12000 17922 12001
rect 17606 11936 17612 12000
rect 17676 11936 17692 12000
rect 17756 11936 17772 12000
rect 17836 11936 17852 12000
rect 17916 11936 17922 12000
rect 17606 11935 17922 11936
rect 22606 12000 22922 12001
rect 22606 11936 22612 12000
rect 22676 11936 22692 12000
rect 22756 11936 22772 12000
rect 22836 11936 22852 12000
rect 22916 11936 22922 12000
rect 22606 11935 22922 11936
rect 27606 12000 27922 12001
rect 27606 11936 27612 12000
rect 27676 11936 27692 12000
rect 27756 11936 27772 12000
rect 27836 11936 27852 12000
rect 27916 11936 27922 12000
rect 27606 11935 27922 11936
rect 32606 12000 32922 12001
rect 32606 11936 32612 12000
rect 32676 11936 32692 12000
rect 32756 11936 32772 12000
rect 32836 11936 32852 12000
rect 32916 11936 32922 12000
rect 32606 11935 32922 11936
rect 37606 12000 37922 12001
rect 37606 11936 37612 12000
rect 37676 11936 37692 12000
rect 37756 11936 37772 12000
rect 37836 11936 37852 12000
rect 37916 11936 37922 12000
rect 37606 11935 37922 11936
rect 1946 11456 2262 11457
rect 1946 11392 1952 11456
rect 2016 11392 2032 11456
rect 2096 11392 2112 11456
rect 2176 11392 2192 11456
rect 2256 11392 2262 11456
rect 1946 11391 2262 11392
rect 6946 11456 7262 11457
rect 6946 11392 6952 11456
rect 7016 11392 7032 11456
rect 7096 11392 7112 11456
rect 7176 11392 7192 11456
rect 7256 11392 7262 11456
rect 6946 11391 7262 11392
rect 11946 11456 12262 11457
rect 11946 11392 11952 11456
rect 12016 11392 12032 11456
rect 12096 11392 12112 11456
rect 12176 11392 12192 11456
rect 12256 11392 12262 11456
rect 11946 11391 12262 11392
rect 16946 11456 17262 11457
rect 16946 11392 16952 11456
rect 17016 11392 17032 11456
rect 17096 11392 17112 11456
rect 17176 11392 17192 11456
rect 17256 11392 17262 11456
rect 16946 11391 17262 11392
rect 21946 11456 22262 11457
rect 21946 11392 21952 11456
rect 22016 11392 22032 11456
rect 22096 11392 22112 11456
rect 22176 11392 22192 11456
rect 22256 11392 22262 11456
rect 21946 11391 22262 11392
rect 26946 11456 27262 11457
rect 26946 11392 26952 11456
rect 27016 11392 27032 11456
rect 27096 11392 27112 11456
rect 27176 11392 27192 11456
rect 27256 11392 27262 11456
rect 26946 11391 27262 11392
rect 31946 11456 32262 11457
rect 31946 11392 31952 11456
rect 32016 11392 32032 11456
rect 32096 11392 32112 11456
rect 32176 11392 32192 11456
rect 32256 11392 32262 11456
rect 31946 11391 32262 11392
rect 36946 11456 37262 11457
rect 36946 11392 36952 11456
rect 37016 11392 37032 11456
rect 37096 11392 37112 11456
rect 37176 11392 37192 11456
rect 37256 11392 37262 11456
rect 36946 11391 37262 11392
rect 33133 10980 33199 10981
rect 33133 10976 33180 10980
rect 33244 10978 33250 10980
rect 33133 10920 33138 10976
rect 33133 10916 33180 10920
rect 33244 10918 33290 10978
rect 33244 10916 33250 10918
rect 33133 10915 33199 10916
rect 2606 10912 2922 10913
rect 2606 10848 2612 10912
rect 2676 10848 2692 10912
rect 2756 10848 2772 10912
rect 2836 10848 2852 10912
rect 2916 10848 2922 10912
rect 2606 10847 2922 10848
rect 7606 10912 7922 10913
rect 7606 10848 7612 10912
rect 7676 10848 7692 10912
rect 7756 10848 7772 10912
rect 7836 10848 7852 10912
rect 7916 10848 7922 10912
rect 7606 10847 7922 10848
rect 12606 10912 12922 10913
rect 12606 10848 12612 10912
rect 12676 10848 12692 10912
rect 12756 10848 12772 10912
rect 12836 10848 12852 10912
rect 12916 10848 12922 10912
rect 12606 10847 12922 10848
rect 17606 10912 17922 10913
rect 17606 10848 17612 10912
rect 17676 10848 17692 10912
rect 17756 10848 17772 10912
rect 17836 10848 17852 10912
rect 17916 10848 17922 10912
rect 17606 10847 17922 10848
rect 22606 10912 22922 10913
rect 22606 10848 22612 10912
rect 22676 10848 22692 10912
rect 22756 10848 22772 10912
rect 22836 10848 22852 10912
rect 22916 10848 22922 10912
rect 22606 10847 22922 10848
rect 27606 10912 27922 10913
rect 27606 10848 27612 10912
rect 27676 10848 27692 10912
rect 27756 10848 27772 10912
rect 27836 10848 27852 10912
rect 27916 10848 27922 10912
rect 27606 10847 27922 10848
rect 32606 10912 32922 10913
rect 32606 10848 32612 10912
rect 32676 10848 32692 10912
rect 32756 10848 32772 10912
rect 32836 10848 32852 10912
rect 32916 10848 32922 10912
rect 32606 10847 32922 10848
rect 37606 10912 37922 10913
rect 37606 10848 37612 10912
rect 37676 10848 37692 10912
rect 37756 10848 37772 10912
rect 37836 10848 37852 10912
rect 37916 10848 37922 10912
rect 37606 10847 37922 10848
rect 1946 10368 2262 10369
rect 1946 10304 1952 10368
rect 2016 10304 2032 10368
rect 2096 10304 2112 10368
rect 2176 10304 2192 10368
rect 2256 10304 2262 10368
rect 1946 10303 2262 10304
rect 6946 10368 7262 10369
rect 6946 10304 6952 10368
rect 7016 10304 7032 10368
rect 7096 10304 7112 10368
rect 7176 10304 7192 10368
rect 7256 10304 7262 10368
rect 6946 10303 7262 10304
rect 11946 10368 12262 10369
rect 11946 10304 11952 10368
rect 12016 10304 12032 10368
rect 12096 10304 12112 10368
rect 12176 10304 12192 10368
rect 12256 10304 12262 10368
rect 11946 10303 12262 10304
rect 16946 10368 17262 10369
rect 16946 10304 16952 10368
rect 17016 10304 17032 10368
rect 17096 10304 17112 10368
rect 17176 10304 17192 10368
rect 17256 10304 17262 10368
rect 16946 10303 17262 10304
rect 21946 10368 22262 10369
rect 21946 10304 21952 10368
rect 22016 10304 22032 10368
rect 22096 10304 22112 10368
rect 22176 10304 22192 10368
rect 22256 10304 22262 10368
rect 21946 10303 22262 10304
rect 26946 10368 27262 10369
rect 26946 10304 26952 10368
rect 27016 10304 27032 10368
rect 27096 10304 27112 10368
rect 27176 10304 27192 10368
rect 27256 10304 27262 10368
rect 26946 10303 27262 10304
rect 31946 10368 32262 10369
rect 31946 10304 31952 10368
rect 32016 10304 32032 10368
rect 32096 10304 32112 10368
rect 32176 10304 32192 10368
rect 32256 10304 32262 10368
rect 31946 10303 32262 10304
rect 36946 10368 37262 10369
rect 36946 10304 36952 10368
rect 37016 10304 37032 10368
rect 37096 10304 37112 10368
rect 37176 10304 37192 10368
rect 37256 10304 37262 10368
rect 36946 10303 37262 10304
rect 2606 9824 2922 9825
rect 2606 9760 2612 9824
rect 2676 9760 2692 9824
rect 2756 9760 2772 9824
rect 2836 9760 2852 9824
rect 2916 9760 2922 9824
rect 2606 9759 2922 9760
rect 7606 9824 7922 9825
rect 7606 9760 7612 9824
rect 7676 9760 7692 9824
rect 7756 9760 7772 9824
rect 7836 9760 7852 9824
rect 7916 9760 7922 9824
rect 7606 9759 7922 9760
rect 12606 9824 12922 9825
rect 12606 9760 12612 9824
rect 12676 9760 12692 9824
rect 12756 9760 12772 9824
rect 12836 9760 12852 9824
rect 12916 9760 12922 9824
rect 12606 9759 12922 9760
rect 17606 9824 17922 9825
rect 17606 9760 17612 9824
rect 17676 9760 17692 9824
rect 17756 9760 17772 9824
rect 17836 9760 17852 9824
rect 17916 9760 17922 9824
rect 17606 9759 17922 9760
rect 22606 9824 22922 9825
rect 22606 9760 22612 9824
rect 22676 9760 22692 9824
rect 22756 9760 22772 9824
rect 22836 9760 22852 9824
rect 22916 9760 22922 9824
rect 22606 9759 22922 9760
rect 27606 9824 27922 9825
rect 27606 9760 27612 9824
rect 27676 9760 27692 9824
rect 27756 9760 27772 9824
rect 27836 9760 27852 9824
rect 27916 9760 27922 9824
rect 27606 9759 27922 9760
rect 32606 9824 32922 9825
rect 32606 9760 32612 9824
rect 32676 9760 32692 9824
rect 32756 9760 32772 9824
rect 32836 9760 32852 9824
rect 32916 9760 32922 9824
rect 32606 9759 32922 9760
rect 37606 9824 37922 9825
rect 37606 9760 37612 9824
rect 37676 9760 37692 9824
rect 37756 9760 37772 9824
rect 37836 9760 37852 9824
rect 37916 9760 37922 9824
rect 37606 9759 37922 9760
rect 7557 9618 7623 9621
rect 33358 9618 33364 9620
rect 7557 9616 33364 9618
rect 7557 9560 7562 9616
rect 7618 9560 33364 9616
rect 7557 9558 33364 9560
rect 7557 9555 7623 9558
rect 33358 9556 33364 9558
rect 33428 9556 33434 9620
rect 1946 9280 2262 9281
rect 1946 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2262 9280
rect 1946 9215 2262 9216
rect 6946 9280 7262 9281
rect 6946 9216 6952 9280
rect 7016 9216 7032 9280
rect 7096 9216 7112 9280
rect 7176 9216 7192 9280
rect 7256 9216 7262 9280
rect 6946 9215 7262 9216
rect 11946 9280 12262 9281
rect 11946 9216 11952 9280
rect 12016 9216 12032 9280
rect 12096 9216 12112 9280
rect 12176 9216 12192 9280
rect 12256 9216 12262 9280
rect 11946 9215 12262 9216
rect 16946 9280 17262 9281
rect 16946 9216 16952 9280
rect 17016 9216 17032 9280
rect 17096 9216 17112 9280
rect 17176 9216 17192 9280
rect 17256 9216 17262 9280
rect 16946 9215 17262 9216
rect 21946 9280 22262 9281
rect 21946 9216 21952 9280
rect 22016 9216 22032 9280
rect 22096 9216 22112 9280
rect 22176 9216 22192 9280
rect 22256 9216 22262 9280
rect 21946 9215 22262 9216
rect 26946 9280 27262 9281
rect 26946 9216 26952 9280
rect 27016 9216 27032 9280
rect 27096 9216 27112 9280
rect 27176 9216 27192 9280
rect 27256 9216 27262 9280
rect 26946 9215 27262 9216
rect 31946 9280 32262 9281
rect 31946 9216 31952 9280
rect 32016 9216 32032 9280
rect 32096 9216 32112 9280
rect 32176 9216 32192 9280
rect 32256 9216 32262 9280
rect 31946 9215 32262 9216
rect 36946 9280 37262 9281
rect 36946 9216 36952 9280
rect 37016 9216 37032 9280
rect 37096 9216 37112 9280
rect 37176 9216 37192 9280
rect 37256 9216 37262 9280
rect 36946 9215 37262 9216
rect 2606 8736 2922 8737
rect 2606 8672 2612 8736
rect 2676 8672 2692 8736
rect 2756 8672 2772 8736
rect 2836 8672 2852 8736
rect 2916 8672 2922 8736
rect 2606 8671 2922 8672
rect 7606 8736 7922 8737
rect 7606 8672 7612 8736
rect 7676 8672 7692 8736
rect 7756 8672 7772 8736
rect 7836 8672 7852 8736
rect 7916 8672 7922 8736
rect 7606 8671 7922 8672
rect 12606 8736 12922 8737
rect 12606 8672 12612 8736
rect 12676 8672 12692 8736
rect 12756 8672 12772 8736
rect 12836 8672 12852 8736
rect 12916 8672 12922 8736
rect 12606 8671 12922 8672
rect 17606 8736 17922 8737
rect 17606 8672 17612 8736
rect 17676 8672 17692 8736
rect 17756 8672 17772 8736
rect 17836 8672 17852 8736
rect 17916 8672 17922 8736
rect 17606 8671 17922 8672
rect 22606 8736 22922 8737
rect 22606 8672 22612 8736
rect 22676 8672 22692 8736
rect 22756 8672 22772 8736
rect 22836 8672 22852 8736
rect 22916 8672 22922 8736
rect 22606 8671 22922 8672
rect 27606 8736 27922 8737
rect 27606 8672 27612 8736
rect 27676 8672 27692 8736
rect 27756 8672 27772 8736
rect 27836 8672 27852 8736
rect 27916 8672 27922 8736
rect 27606 8671 27922 8672
rect 32606 8736 32922 8737
rect 32606 8672 32612 8736
rect 32676 8672 32692 8736
rect 32756 8672 32772 8736
rect 32836 8672 32852 8736
rect 32916 8672 32922 8736
rect 32606 8671 32922 8672
rect 37606 8736 37922 8737
rect 37606 8672 37612 8736
rect 37676 8672 37692 8736
rect 37756 8672 37772 8736
rect 37836 8672 37852 8736
rect 37916 8672 37922 8736
rect 37606 8671 37922 8672
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 6946 8192 7262 8193
rect 6946 8128 6952 8192
rect 7016 8128 7032 8192
rect 7096 8128 7112 8192
rect 7176 8128 7192 8192
rect 7256 8128 7262 8192
rect 6946 8127 7262 8128
rect 11946 8192 12262 8193
rect 11946 8128 11952 8192
rect 12016 8128 12032 8192
rect 12096 8128 12112 8192
rect 12176 8128 12192 8192
rect 12256 8128 12262 8192
rect 11946 8127 12262 8128
rect 16946 8192 17262 8193
rect 16946 8128 16952 8192
rect 17016 8128 17032 8192
rect 17096 8128 17112 8192
rect 17176 8128 17192 8192
rect 17256 8128 17262 8192
rect 16946 8127 17262 8128
rect 21946 8192 22262 8193
rect 21946 8128 21952 8192
rect 22016 8128 22032 8192
rect 22096 8128 22112 8192
rect 22176 8128 22192 8192
rect 22256 8128 22262 8192
rect 21946 8127 22262 8128
rect 26946 8192 27262 8193
rect 26946 8128 26952 8192
rect 27016 8128 27032 8192
rect 27096 8128 27112 8192
rect 27176 8128 27192 8192
rect 27256 8128 27262 8192
rect 26946 8127 27262 8128
rect 31946 8192 32262 8193
rect 31946 8128 31952 8192
rect 32016 8128 32032 8192
rect 32096 8128 32112 8192
rect 32176 8128 32192 8192
rect 32256 8128 32262 8192
rect 31946 8127 32262 8128
rect 36946 8192 37262 8193
rect 36946 8128 36952 8192
rect 37016 8128 37032 8192
rect 37096 8128 37112 8192
rect 37176 8128 37192 8192
rect 37256 8128 37262 8192
rect 36946 8127 37262 8128
rect 18873 7850 18939 7853
rect 33542 7850 33548 7852
rect 18873 7848 33548 7850
rect 18873 7792 18878 7848
rect 18934 7792 33548 7848
rect 18873 7790 33548 7792
rect 18873 7787 18939 7790
rect 33542 7788 33548 7790
rect 33612 7788 33618 7852
rect 2606 7648 2922 7649
rect 2606 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2922 7648
rect 2606 7583 2922 7584
rect 7606 7648 7922 7649
rect 7606 7584 7612 7648
rect 7676 7584 7692 7648
rect 7756 7584 7772 7648
rect 7836 7584 7852 7648
rect 7916 7584 7922 7648
rect 7606 7583 7922 7584
rect 12606 7648 12922 7649
rect 12606 7584 12612 7648
rect 12676 7584 12692 7648
rect 12756 7584 12772 7648
rect 12836 7584 12852 7648
rect 12916 7584 12922 7648
rect 12606 7583 12922 7584
rect 17606 7648 17922 7649
rect 17606 7584 17612 7648
rect 17676 7584 17692 7648
rect 17756 7584 17772 7648
rect 17836 7584 17852 7648
rect 17916 7584 17922 7648
rect 17606 7583 17922 7584
rect 22606 7648 22922 7649
rect 22606 7584 22612 7648
rect 22676 7584 22692 7648
rect 22756 7584 22772 7648
rect 22836 7584 22852 7648
rect 22916 7584 22922 7648
rect 22606 7583 22922 7584
rect 27606 7648 27922 7649
rect 27606 7584 27612 7648
rect 27676 7584 27692 7648
rect 27756 7584 27772 7648
rect 27836 7584 27852 7648
rect 27916 7584 27922 7648
rect 27606 7583 27922 7584
rect 32606 7648 32922 7649
rect 32606 7584 32612 7648
rect 32676 7584 32692 7648
rect 32756 7584 32772 7648
rect 32836 7584 32852 7648
rect 32916 7584 32922 7648
rect 32606 7583 32922 7584
rect 37606 7648 37922 7649
rect 37606 7584 37612 7648
rect 37676 7584 37692 7648
rect 37756 7584 37772 7648
rect 37836 7584 37852 7648
rect 37916 7584 37922 7648
rect 37606 7583 37922 7584
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 6946 7104 7262 7105
rect 6946 7040 6952 7104
rect 7016 7040 7032 7104
rect 7096 7040 7112 7104
rect 7176 7040 7192 7104
rect 7256 7040 7262 7104
rect 6946 7039 7262 7040
rect 11946 7104 12262 7105
rect 11946 7040 11952 7104
rect 12016 7040 12032 7104
rect 12096 7040 12112 7104
rect 12176 7040 12192 7104
rect 12256 7040 12262 7104
rect 11946 7039 12262 7040
rect 16946 7104 17262 7105
rect 16946 7040 16952 7104
rect 17016 7040 17032 7104
rect 17096 7040 17112 7104
rect 17176 7040 17192 7104
rect 17256 7040 17262 7104
rect 16946 7039 17262 7040
rect 21946 7104 22262 7105
rect 21946 7040 21952 7104
rect 22016 7040 22032 7104
rect 22096 7040 22112 7104
rect 22176 7040 22192 7104
rect 22256 7040 22262 7104
rect 21946 7039 22262 7040
rect 26946 7104 27262 7105
rect 26946 7040 26952 7104
rect 27016 7040 27032 7104
rect 27096 7040 27112 7104
rect 27176 7040 27192 7104
rect 27256 7040 27262 7104
rect 26946 7039 27262 7040
rect 31946 7104 32262 7105
rect 31946 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32262 7104
rect 31946 7039 32262 7040
rect 36946 7104 37262 7105
rect 36946 7040 36952 7104
rect 37016 7040 37032 7104
rect 37096 7040 37112 7104
rect 37176 7040 37192 7104
rect 37256 7040 37262 7104
rect 36946 7039 37262 7040
rect 2606 6560 2922 6561
rect 2606 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2922 6560
rect 2606 6495 2922 6496
rect 7606 6560 7922 6561
rect 7606 6496 7612 6560
rect 7676 6496 7692 6560
rect 7756 6496 7772 6560
rect 7836 6496 7852 6560
rect 7916 6496 7922 6560
rect 7606 6495 7922 6496
rect 12606 6560 12922 6561
rect 12606 6496 12612 6560
rect 12676 6496 12692 6560
rect 12756 6496 12772 6560
rect 12836 6496 12852 6560
rect 12916 6496 12922 6560
rect 12606 6495 12922 6496
rect 17606 6560 17922 6561
rect 17606 6496 17612 6560
rect 17676 6496 17692 6560
rect 17756 6496 17772 6560
rect 17836 6496 17852 6560
rect 17916 6496 17922 6560
rect 17606 6495 17922 6496
rect 22606 6560 22922 6561
rect 22606 6496 22612 6560
rect 22676 6496 22692 6560
rect 22756 6496 22772 6560
rect 22836 6496 22852 6560
rect 22916 6496 22922 6560
rect 22606 6495 22922 6496
rect 27606 6560 27922 6561
rect 27606 6496 27612 6560
rect 27676 6496 27692 6560
rect 27756 6496 27772 6560
rect 27836 6496 27852 6560
rect 27916 6496 27922 6560
rect 27606 6495 27922 6496
rect 32606 6560 32922 6561
rect 32606 6496 32612 6560
rect 32676 6496 32692 6560
rect 32756 6496 32772 6560
rect 32836 6496 32852 6560
rect 32916 6496 32922 6560
rect 32606 6495 32922 6496
rect 37606 6560 37922 6561
rect 37606 6496 37612 6560
rect 37676 6496 37692 6560
rect 37756 6496 37772 6560
rect 37836 6496 37852 6560
rect 37916 6496 37922 6560
rect 37606 6495 37922 6496
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 6946 6016 7262 6017
rect 6946 5952 6952 6016
rect 7016 5952 7032 6016
rect 7096 5952 7112 6016
rect 7176 5952 7192 6016
rect 7256 5952 7262 6016
rect 6946 5951 7262 5952
rect 11946 6016 12262 6017
rect 11946 5952 11952 6016
rect 12016 5952 12032 6016
rect 12096 5952 12112 6016
rect 12176 5952 12192 6016
rect 12256 5952 12262 6016
rect 11946 5951 12262 5952
rect 16946 6016 17262 6017
rect 16946 5952 16952 6016
rect 17016 5952 17032 6016
rect 17096 5952 17112 6016
rect 17176 5952 17192 6016
rect 17256 5952 17262 6016
rect 16946 5951 17262 5952
rect 21946 6016 22262 6017
rect 21946 5952 21952 6016
rect 22016 5952 22032 6016
rect 22096 5952 22112 6016
rect 22176 5952 22192 6016
rect 22256 5952 22262 6016
rect 21946 5951 22262 5952
rect 26946 6016 27262 6017
rect 26946 5952 26952 6016
rect 27016 5952 27032 6016
rect 27096 5952 27112 6016
rect 27176 5952 27192 6016
rect 27256 5952 27262 6016
rect 26946 5951 27262 5952
rect 31946 6016 32262 6017
rect 31946 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32262 6016
rect 31946 5951 32262 5952
rect 36946 6016 37262 6017
rect 36946 5952 36952 6016
rect 37016 5952 37032 6016
rect 37096 5952 37112 6016
rect 37176 5952 37192 6016
rect 37256 5952 37262 6016
rect 36946 5951 37262 5952
rect 2606 5472 2922 5473
rect 2606 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2922 5472
rect 2606 5407 2922 5408
rect 7606 5472 7922 5473
rect 7606 5408 7612 5472
rect 7676 5408 7692 5472
rect 7756 5408 7772 5472
rect 7836 5408 7852 5472
rect 7916 5408 7922 5472
rect 7606 5407 7922 5408
rect 12606 5472 12922 5473
rect 12606 5408 12612 5472
rect 12676 5408 12692 5472
rect 12756 5408 12772 5472
rect 12836 5408 12852 5472
rect 12916 5408 12922 5472
rect 12606 5407 12922 5408
rect 17606 5472 17922 5473
rect 17606 5408 17612 5472
rect 17676 5408 17692 5472
rect 17756 5408 17772 5472
rect 17836 5408 17852 5472
rect 17916 5408 17922 5472
rect 17606 5407 17922 5408
rect 22606 5472 22922 5473
rect 22606 5408 22612 5472
rect 22676 5408 22692 5472
rect 22756 5408 22772 5472
rect 22836 5408 22852 5472
rect 22916 5408 22922 5472
rect 22606 5407 22922 5408
rect 27606 5472 27922 5473
rect 27606 5408 27612 5472
rect 27676 5408 27692 5472
rect 27756 5408 27772 5472
rect 27836 5408 27852 5472
rect 27916 5408 27922 5472
rect 27606 5407 27922 5408
rect 32606 5472 32922 5473
rect 32606 5408 32612 5472
rect 32676 5408 32692 5472
rect 32756 5408 32772 5472
rect 32836 5408 32852 5472
rect 32916 5408 32922 5472
rect 32606 5407 32922 5408
rect 37606 5472 37922 5473
rect 37606 5408 37612 5472
rect 37676 5408 37692 5472
rect 37756 5408 37772 5472
rect 37836 5408 37852 5472
rect 37916 5408 37922 5472
rect 37606 5407 37922 5408
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 1946 4863 2262 4864
rect 6946 4928 7262 4929
rect 6946 4864 6952 4928
rect 7016 4864 7032 4928
rect 7096 4864 7112 4928
rect 7176 4864 7192 4928
rect 7256 4864 7262 4928
rect 6946 4863 7262 4864
rect 11946 4928 12262 4929
rect 11946 4864 11952 4928
rect 12016 4864 12032 4928
rect 12096 4864 12112 4928
rect 12176 4864 12192 4928
rect 12256 4864 12262 4928
rect 11946 4863 12262 4864
rect 16946 4928 17262 4929
rect 16946 4864 16952 4928
rect 17016 4864 17032 4928
rect 17096 4864 17112 4928
rect 17176 4864 17192 4928
rect 17256 4864 17262 4928
rect 16946 4863 17262 4864
rect 21946 4928 22262 4929
rect 21946 4864 21952 4928
rect 22016 4864 22032 4928
rect 22096 4864 22112 4928
rect 22176 4864 22192 4928
rect 22256 4864 22262 4928
rect 21946 4863 22262 4864
rect 26946 4928 27262 4929
rect 26946 4864 26952 4928
rect 27016 4864 27032 4928
rect 27096 4864 27112 4928
rect 27176 4864 27192 4928
rect 27256 4864 27262 4928
rect 26946 4863 27262 4864
rect 31946 4928 32262 4929
rect 31946 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32262 4928
rect 31946 4863 32262 4864
rect 36946 4928 37262 4929
rect 36946 4864 36952 4928
rect 37016 4864 37032 4928
rect 37096 4864 37112 4928
rect 37176 4864 37192 4928
rect 37256 4864 37262 4928
rect 36946 4863 37262 4864
rect 2606 4384 2922 4385
rect 2606 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2922 4384
rect 2606 4319 2922 4320
rect 7606 4384 7922 4385
rect 7606 4320 7612 4384
rect 7676 4320 7692 4384
rect 7756 4320 7772 4384
rect 7836 4320 7852 4384
rect 7916 4320 7922 4384
rect 7606 4319 7922 4320
rect 12606 4384 12922 4385
rect 12606 4320 12612 4384
rect 12676 4320 12692 4384
rect 12756 4320 12772 4384
rect 12836 4320 12852 4384
rect 12916 4320 12922 4384
rect 12606 4319 12922 4320
rect 17606 4384 17922 4385
rect 17606 4320 17612 4384
rect 17676 4320 17692 4384
rect 17756 4320 17772 4384
rect 17836 4320 17852 4384
rect 17916 4320 17922 4384
rect 17606 4319 17922 4320
rect 22606 4384 22922 4385
rect 22606 4320 22612 4384
rect 22676 4320 22692 4384
rect 22756 4320 22772 4384
rect 22836 4320 22852 4384
rect 22916 4320 22922 4384
rect 22606 4319 22922 4320
rect 27606 4384 27922 4385
rect 27606 4320 27612 4384
rect 27676 4320 27692 4384
rect 27756 4320 27772 4384
rect 27836 4320 27852 4384
rect 27916 4320 27922 4384
rect 27606 4319 27922 4320
rect 32606 4384 32922 4385
rect 32606 4320 32612 4384
rect 32676 4320 32692 4384
rect 32756 4320 32772 4384
rect 32836 4320 32852 4384
rect 32916 4320 32922 4384
rect 32606 4319 32922 4320
rect 37606 4384 37922 4385
rect 37606 4320 37612 4384
rect 37676 4320 37692 4384
rect 37756 4320 37772 4384
rect 37836 4320 37852 4384
rect 37916 4320 37922 4384
rect 37606 4319 37922 4320
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 6946 3840 7262 3841
rect 6946 3776 6952 3840
rect 7016 3776 7032 3840
rect 7096 3776 7112 3840
rect 7176 3776 7192 3840
rect 7256 3776 7262 3840
rect 6946 3775 7262 3776
rect 11946 3840 12262 3841
rect 11946 3776 11952 3840
rect 12016 3776 12032 3840
rect 12096 3776 12112 3840
rect 12176 3776 12192 3840
rect 12256 3776 12262 3840
rect 11946 3775 12262 3776
rect 16946 3840 17262 3841
rect 16946 3776 16952 3840
rect 17016 3776 17032 3840
rect 17096 3776 17112 3840
rect 17176 3776 17192 3840
rect 17256 3776 17262 3840
rect 16946 3775 17262 3776
rect 21946 3840 22262 3841
rect 21946 3776 21952 3840
rect 22016 3776 22032 3840
rect 22096 3776 22112 3840
rect 22176 3776 22192 3840
rect 22256 3776 22262 3840
rect 21946 3775 22262 3776
rect 26946 3840 27262 3841
rect 26946 3776 26952 3840
rect 27016 3776 27032 3840
rect 27096 3776 27112 3840
rect 27176 3776 27192 3840
rect 27256 3776 27262 3840
rect 26946 3775 27262 3776
rect 31946 3840 32262 3841
rect 31946 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32262 3840
rect 31946 3775 32262 3776
rect 36946 3840 37262 3841
rect 36946 3776 36952 3840
rect 37016 3776 37032 3840
rect 37096 3776 37112 3840
rect 37176 3776 37192 3840
rect 37256 3776 37262 3840
rect 36946 3775 37262 3776
rect 2606 3296 2922 3297
rect 2606 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2922 3296
rect 2606 3231 2922 3232
rect 7606 3296 7922 3297
rect 7606 3232 7612 3296
rect 7676 3232 7692 3296
rect 7756 3232 7772 3296
rect 7836 3232 7852 3296
rect 7916 3232 7922 3296
rect 7606 3231 7922 3232
rect 12606 3296 12922 3297
rect 12606 3232 12612 3296
rect 12676 3232 12692 3296
rect 12756 3232 12772 3296
rect 12836 3232 12852 3296
rect 12916 3232 12922 3296
rect 12606 3231 12922 3232
rect 17606 3296 17922 3297
rect 17606 3232 17612 3296
rect 17676 3232 17692 3296
rect 17756 3232 17772 3296
rect 17836 3232 17852 3296
rect 17916 3232 17922 3296
rect 17606 3231 17922 3232
rect 22606 3296 22922 3297
rect 22606 3232 22612 3296
rect 22676 3232 22692 3296
rect 22756 3232 22772 3296
rect 22836 3232 22852 3296
rect 22916 3232 22922 3296
rect 22606 3231 22922 3232
rect 27606 3296 27922 3297
rect 27606 3232 27612 3296
rect 27676 3232 27692 3296
rect 27756 3232 27772 3296
rect 27836 3232 27852 3296
rect 27916 3232 27922 3296
rect 27606 3231 27922 3232
rect 32606 3296 32922 3297
rect 32606 3232 32612 3296
rect 32676 3232 32692 3296
rect 32756 3232 32772 3296
rect 32836 3232 32852 3296
rect 32916 3232 32922 3296
rect 32606 3231 32922 3232
rect 37606 3296 37922 3297
rect 37606 3232 37612 3296
rect 37676 3232 37692 3296
rect 37756 3232 37772 3296
rect 37836 3232 37852 3296
rect 37916 3232 37922 3296
rect 37606 3231 37922 3232
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 6946 2752 7262 2753
rect 6946 2688 6952 2752
rect 7016 2688 7032 2752
rect 7096 2688 7112 2752
rect 7176 2688 7192 2752
rect 7256 2688 7262 2752
rect 6946 2687 7262 2688
rect 11946 2752 12262 2753
rect 11946 2688 11952 2752
rect 12016 2688 12032 2752
rect 12096 2688 12112 2752
rect 12176 2688 12192 2752
rect 12256 2688 12262 2752
rect 11946 2687 12262 2688
rect 16946 2752 17262 2753
rect 16946 2688 16952 2752
rect 17016 2688 17032 2752
rect 17096 2688 17112 2752
rect 17176 2688 17192 2752
rect 17256 2688 17262 2752
rect 16946 2687 17262 2688
rect 21946 2752 22262 2753
rect 21946 2688 21952 2752
rect 22016 2688 22032 2752
rect 22096 2688 22112 2752
rect 22176 2688 22192 2752
rect 22256 2688 22262 2752
rect 21946 2687 22262 2688
rect 26946 2752 27262 2753
rect 26946 2688 26952 2752
rect 27016 2688 27032 2752
rect 27096 2688 27112 2752
rect 27176 2688 27192 2752
rect 27256 2688 27262 2752
rect 26946 2687 27262 2688
rect 31946 2752 32262 2753
rect 31946 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32262 2752
rect 31946 2687 32262 2688
rect 36946 2752 37262 2753
rect 36946 2688 36952 2752
rect 37016 2688 37032 2752
rect 37096 2688 37112 2752
rect 37176 2688 37192 2752
rect 37256 2688 37262 2752
rect 36946 2687 37262 2688
rect 2606 2208 2922 2209
rect 2606 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2922 2208
rect 2606 2143 2922 2144
rect 7606 2208 7922 2209
rect 7606 2144 7612 2208
rect 7676 2144 7692 2208
rect 7756 2144 7772 2208
rect 7836 2144 7852 2208
rect 7916 2144 7922 2208
rect 7606 2143 7922 2144
rect 12606 2208 12922 2209
rect 12606 2144 12612 2208
rect 12676 2144 12692 2208
rect 12756 2144 12772 2208
rect 12836 2144 12852 2208
rect 12916 2144 12922 2208
rect 12606 2143 12922 2144
rect 17606 2208 17922 2209
rect 17606 2144 17612 2208
rect 17676 2144 17692 2208
rect 17756 2144 17772 2208
rect 17836 2144 17852 2208
rect 17916 2144 17922 2208
rect 17606 2143 17922 2144
rect 22606 2208 22922 2209
rect 22606 2144 22612 2208
rect 22676 2144 22692 2208
rect 22756 2144 22772 2208
rect 22836 2144 22852 2208
rect 22916 2144 22922 2208
rect 22606 2143 22922 2144
rect 27606 2208 27922 2209
rect 27606 2144 27612 2208
rect 27676 2144 27692 2208
rect 27756 2144 27772 2208
rect 27836 2144 27852 2208
rect 27916 2144 27922 2208
rect 27606 2143 27922 2144
rect 32606 2208 32922 2209
rect 32606 2144 32612 2208
rect 32676 2144 32692 2208
rect 32756 2144 32772 2208
rect 32836 2144 32852 2208
rect 32916 2144 32922 2208
rect 32606 2143 32922 2144
rect 37606 2208 37922 2209
rect 37606 2144 37612 2208
rect 37676 2144 37692 2208
rect 37756 2144 37772 2208
rect 37836 2144 37852 2208
rect 37916 2144 37922 2208
rect 37606 2143 37922 2144
<< via3 >>
rect 2612 69660 2676 69664
rect 2612 69604 2616 69660
rect 2616 69604 2672 69660
rect 2672 69604 2676 69660
rect 2612 69600 2676 69604
rect 2692 69660 2756 69664
rect 2692 69604 2696 69660
rect 2696 69604 2752 69660
rect 2752 69604 2756 69660
rect 2692 69600 2756 69604
rect 2772 69660 2836 69664
rect 2772 69604 2776 69660
rect 2776 69604 2832 69660
rect 2832 69604 2836 69660
rect 2772 69600 2836 69604
rect 2852 69660 2916 69664
rect 2852 69604 2856 69660
rect 2856 69604 2912 69660
rect 2912 69604 2916 69660
rect 2852 69600 2916 69604
rect 7612 69660 7676 69664
rect 7612 69604 7616 69660
rect 7616 69604 7672 69660
rect 7672 69604 7676 69660
rect 7612 69600 7676 69604
rect 7692 69660 7756 69664
rect 7692 69604 7696 69660
rect 7696 69604 7752 69660
rect 7752 69604 7756 69660
rect 7692 69600 7756 69604
rect 7772 69660 7836 69664
rect 7772 69604 7776 69660
rect 7776 69604 7832 69660
rect 7832 69604 7836 69660
rect 7772 69600 7836 69604
rect 7852 69660 7916 69664
rect 7852 69604 7856 69660
rect 7856 69604 7912 69660
rect 7912 69604 7916 69660
rect 7852 69600 7916 69604
rect 12612 69660 12676 69664
rect 12612 69604 12616 69660
rect 12616 69604 12672 69660
rect 12672 69604 12676 69660
rect 12612 69600 12676 69604
rect 12692 69660 12756 69664
rect 12692 69604 12696 69660
rect 12696 69604 12752 69660
rect 12752 69604 12756 69660
rect 12692 69600 12756 69604
rect 12772 69660 12836 69664
rect 12772 69604 12776 69660
rect 12776 69604 12832 69660
rect 12832 69604 12836 69660
rect 12772 69600 12836 69604
rect 12852 69660 12916 69664
rect 12852 69604 12856 69660
rect 12856 69604 12912 69660
rect 12912 69604 12916 69660
rect 12852 69600 12916 69604
rect 17612 69660 17676 69664
rect 17612 69604 17616 69660
rect 17616 69604 17672 69660
rect 17672 69604 17676 69660
rect 17612 69600 17676 69604
rect 17692 69660 17756 69664
rect 17692 69604 17696 69660
rect 17696 69604 17752 69660
rect 17752 69604 17756 69660
rect 17692 69600 17756 69604
rect 17772 69660 17836 69664
rect 17772 69604 17776 69660
rect 17776 69604 17832 69660
rect 17832 69604 17836 69660
rect 17772 69600 17836 69604
rect 17852 69660 17916 69664
rect 17852 69604 17856 69660
rect 17856 69604 17912 69660
rect 17912 69604 17916 69660
rect 17852 69600 17916 69604
rect 22612 69660 22676 69664
rect 22612 69604 22616 69660
rect 22616 69604 22672 69660
rect 22672 69604 22676 69660
rect 22612 69600 22676 69604
rect 22692 69660 22756 69664
rect 22692 69604 22696 69660
rect 22696 69604 22752 69660
rect 22752 69604 22756 69660
rect 22692 69600 22756 69604
rect 22772 69660 22836 69664
rect 22772 69604 22776 69660
rect 22776 69604 22832 69660
rect 22832 69604 22836 69660
rect 22772 69600 22836 69604
rect 22852 69660 22916 69664
rect 22852 69604 22856 69660
rect 22856 69604 22912 69660
rect 22912 69604 22916 69660
rect 22852 69600 22916 69604
rect 27612 69660 27676 69664
rect 27612 69604 27616 69660
rect 27616 69604 27672 69660
rect 27672 69604 27676 69660
rect 27612 69600 27676 69604
rect 27692 69660 27756 69664
rect 27692 69604 27696 69660
rect 27696 69604 27752 69660
rect 27752 69604 27756 69660
rect 27692 69600 27756 69604
rect 27772 69660 27836 69664
rect 27772 69604 27776 69660
rect 27776 69604 27832 69660
rect 27832 69604 27836 69660
rect 27772 69600 27836 69604
rect 27852 69660 27916 69664
rect 27852 69604 27856 69660
rect 27856 69604 27912 69660
rect 27912 69604 27916 69660
rect 27852 69600 27916 69604
rect 32612 69660 32676 69664
rect 32612 69604 32616 69660
rect 32616 69604 32672 69660
rect 32672 69604 32676 69660
rect 32612 69600 32676 69604
rect 32692 69660 32756 69664
rect 32692 69604 32696 69660
rect 32696 69604 32752 69660
rect 32752 69604 32756 69660
rect 32692 69600 32756 69604
rect 32772 69660 32836 69664
rect 32772 69604 32776 69660
rect 32776 69604 32832 69660
rect 32832 69604 32836 69660
rect 32772 69600 32836 69604
rect 32852 69660 32916 69664
rect 32852 69604 32856 69660
rect 32856 69604 32912 69660
rect 32912 69604 32916 69660
rect 32852 69600 32916 69604
rect 37612 69660 37676 69664
rect 37612 69604 37616 69660
rect 37616 69604 37672 69660
rect 37672 69604 37676 69660
rect 37612 69600 37676 69604
rect 37692 69660 37756 69664
rect 37692 69604 37696 69660
rect 37696 69604 37752 69660
rect 37752 69604 37756 69660
rect 37692 69600 37756 69604
rect 37772 69660 37836 69664
rect 37772 69604 37776 69660
rect 37776 69604 37832 69660
rect 37832 69604 37836 69660
rect 37772 69600 37836 69604
rect 37852 69660 37916 69664
rect 37852 69604 37856 69660
rect 37856 69604 37912 69660
rect 37912 69604 37916 69660
rect 37852 69600 37916 69604
rect 1952 69116 2016 69120
rect 1952 69060 1956 69116
rect 1956 69060 2012 69116
rect 2012 69060 2016 69116
rect 1952 69056 2016 69060
rect 2032 69116 2096 69120
rect 2032 69060 2036 69116
rect 2036 69060 2092 69116
rect 2092 69060 2096 69116
rect 2032 69056 2096 69060
rect 2112 69116 2176 69120
rect 2112 69060 2116 69116
rect 2116 69060 2172 69116
rect 2172 69060 2176 69116
rect 2112 69056 2176 69060
rect 2192 69116 2256 69120
rect 2192 69060 2196 69116
rect 2196 69060 2252 69116
rect 2252 69060 2256 69116
rect 2192 69056 2256 69060
rect 6952 69116 7016 69120
rect 6952 69060 6956 69116
rect 6956 69060 7012 69116
rect 7012 69060 7016 69116
rect 6952 69056 7016 69060
rect 7032 69116 7096 69120
rect 7032 69060 7036 69116
rect 7036 69060 7092 69116
rect 7092 69060 7096 69116
rect 7032 69056 7096 69060
rect 7112 69116 7176 69120
rect 7112 69060 7116 69116
rect 7116 69060 7172 69116
rect 7172 69060 7176 69116
rect 7112 69056 7176 69060
rect 7192 69116 7256 69120
rect 7192 69060 7196 69116
rect 7196 69060 7252 69116
rect 7252 69060 7256 69116
rect 7192 69056 7256 69060
rect 11952 69116 12016 69120
rect 11952 69060 11956 69116
rect 11956 69060 12012 69116
rect 12012 69060 12016 69116
rect 11952 69056 12016 69060
rect 12032 69116 12096 69120
rect 12032 69060 12036 69116
rect 12036 69060 12092 69116
rect 12092 69060 12096 69116
rect 12032 69056 12096 69060
rect 12112 69116 12176 69120
rect 12112 69060 12116 69116
rect 12116 69060 12172 69116
rect 12172 69060 12176 69116
rect 12112 69056 12176 69060
rect 12192 69116 12256 69120
rect 12192 69060 12196 69116
rect 12196 69060 12252 69116
rect 12252 69060 12256 69116
rect 12192 69056 12256 69060
rect 16952 69116 17016 69120
rect 16952 69060 16956 69116
rect 16956 69060 17012 69116
rect 17012 69060 17016 69116
rect 16952 69056 17016 69060
rect 17032 69116 17096 69120
rect 17032 69060 17036 69116
rect 17036 69060 17092 69116
rect 17092 69060 17096 69116
rect 17032 69056 17096 69060
rect 17112 69116 17176 69120
rect 17112 69060 17116 69116
rect 17116 69060 17172 69116
rect 17172 69060 17176 69116
rect 17112 69056 17176 69060
rect 17192 69116 17256 69120
rect 17192 69060 17196 69116
rect 17196 69060 17252 69116
rect 17252 69060 17256 69116
rect 17192 69056 17256 69060
rect 21952 69116 22016 69120
rect 21952 69060 21956 69116
rect 21956 69060 22012 69116
rect 22012 69060 22016 69116
rect 21952 69056 22016 69060
rect 22032 69116 22096 69120
rect 22032 69060 22036 69116
rect 22036 69060 22092 69116
rect 22092 69060 22096 69116
rect 22032 69056 22096 69060
rect 22112 69116 22176 69120
rect 22112 69060 22116 69116
rect 22116 69060 22172 69116
rect 22172 69060 22176 69116
rect 22112 69056 22176 69060
rect 22192 69116 22256 69120
rect 22192 69060 22196 69116
rect 22196 69060 22252 69116
rect 22252 69060 22256 69116
rect 22192 69056 22256 69060
rect 26952 69116 27016 69120
rect 26952 69060 26956 69116
rect 26956 69060 27012 69116
rect 27012 69060 27016 69116
rect 26952 69056 27016 69060
rect 27032 69116 27096 69120
rect 27032 69060 27036 69116
rect 27036 69060 27092 69116
rect 27092 69060 27096 69116
rect 27032 69056 27096 69060
rect 27112 69116 27176 69120
rect 27112 69060 27116 69116
rect 27116 69060 27172 69116
rect 27172 69060 27176 69116
rect 27112 69056 27176 69060
rect 27192 69116 27256 69120
rect 27192 69060 27196 69116
rect 27196 69060 27252 69116
rect 27252 69060 27256 69116
rect 27192 69056 27256 69060
rect 31952 69116 32016 69120
rect 31952 69060 31956 69116
rect 31956 69060 32012 69116
rect 32012 69060 32016 69116
rect 31952 69056 32016 69060
rect 32032 69116 32096 69120
rect 32032 69060 32036 69116
rect 32036 69060 32092 69116
rect 32092 69060 32096 69116
rect 32032 69056 32096 69060
rect 32112 69116 32176 69120
rect 32112 69060 32116 69116
rect 32116 69060 32172 69116
rect 32172 69060 32176 69116
rect 32112 69056 32176 69060
rect 32192 69116 32256 69120
rect 32192 69060 32196 69116
rect 32196 69060 32252 69116
rect 32252 69060 32256 69116
rect 32192 69056 32256 69060
rect 36952 69116 37016 69120
rect 36952 69060 36956 69116
rect 36956 69060 37012 69116
rect 37012 69060 37016 69116
rect 36952 69056 37016 69060
rect 37032 69116 37096 69120
rect 37032 69060 37036 69116
rect 37036 69060 37092 69116
rect 37092 69060 37096 69116
rect 37032 69056 37096 69060
rect 37112 69116 37176 69120
rect 37112 69060 37116 69116
rect 37116 69060 37172 69116
rect 37172 69060 37176 69116
rect 37112 69056 37176 69060
rect 37192 69116 37256 69120
rect 37192 69060 37196 69116
rect 37196 69060 37252 69116
rect 37252 69060 37256 69116
rect 37192 69056 37256 69060
rect 2612 68572 2676 68576
rect 2612 68516 2616 68572
rect 2616 68516 2672 68572
rect 2672 68516 2676 68572
rect 2612 68512 2676 68516
rect 2692 68572 2756 68576
rect 2692 68516 2696 68572
rect 2696 68516 2752 68572
rect 2752 68516 2756 68572
rect 2692 68512 2756 68516
rect 2772 68572 2836 68576
rect 2772 68516 2776 68572
rect 2776 68516 2832 68572
rect 2832 68516 2836 68572
rect 2772 68512 2836 68516
rect 2852 68572 2916 68576
rect 2852 68516 2856 68572
rect 2856 68516 2912 68572
rect 2912 68516 2916 68572
rect 2852 68512 2916 68516
rect 7612 68572 7676 68576
rect 7612 68516 7616 68572
rect 7616 68516 7672 68572
rect 7672 68516 7676 68572
rect 7612 68512 7676 68516
rect 7692 68572 7756 68576
rect 7692 68516 7696 68572
rect 7696 68516 7752 68572
rect 7752 68516 7756 68572
rect 7692 68512 7756 68516
rect 7772 68572 7836 68576
rect 7772 68516 7776 68572
rect 7776 68516 7832 68572
rect 7832 68516 7836 68572
rect 7772 68512 7836 68516
rect 7852 68572 7916 68576
rect 7852 68516 7856 68572
rect 7856 68516 7912 68572
rect 7912 68516 7916 68572
rect 7852 68512 7916 68516
rect 12612 68572 12676 68576
rect 12612 68516 12616 68572
rect 12616 68516 12672 68572
rect 12672 68516 12676 68572
rect 12612 68512 12676 68516
rect 12692 68572 12756 68576
rect 12692 68516 12696 68572
rect 12696 68516 12752 68572
rect 12752 68516 12756 68572
rect 12692 68512 12756 68516
rect 12772 68572 12836 68576
rect 12772 68516 12776 68572
rect 12776 68516 12832 68572
rect 12832 68516 12836 68572
rect 12772 68512 12836 68516
rect 12852 68572 12916 68576
rect 12852 68516 12856 68572
rect 12856 68516 12912 68572
rect 12912 68516 12916 68572
rect 12852 68512 12916 68516
rect 17612 68572 17676 68576
rect 17612 68516 17616 68572
rect 17616 68516 17672 68572
rect 17672 68516 17676 68572
rect 17612 68512 17676 68516
rect 17692 68572 17756 68576
rect 17692 68516 17696 68572
rect 17696 68516 17752 68572
rect 17752 68516 17756 68572
rect 17692 68512 17756 68516
rect 17772 68572 17836 68576
rect 17772 68516 17776 68572
rect 17776 68516 17832 68572
rect 17832 68516 17836 68572
rect 17772 68512 17836 68516
rect 17852 68572 17916 68576
rect 17852 68516 17856 68572
rect 17856 68516 17912 68572
rect 17912 68516 17916 68572
rect 17852 68512 17916 68516
rect 22612 68572 22676 68576
rect 22612 68516 22616 68572
rect 22616 68516 22672 68572
rect 22672 68516 22676 68572
rect 22612 68512 22676 68516
rect 22692 68572 22756 68576
rect 22692 68516 22696 68572
rect 22696 68516 22752 68572
rect 22752 68516 22756 68572
rect 22692 68512 22756 68516
rect 22772 68572 22836 68576
rect 22772 68516 22776 68572
rect 22776 68516 22832 68572
rect 22832 68516 22836 68572
rect 22772 68512 22836 68516
rect 22852 68572 22916 68576
rect 22852 68516 22856 68572
rect 22856 68516 22912 68572
rect 22912 68516 22916 68572
rect 22852 68512 22916 68516
rect 27612 68572 27676 68576
rect 27612 68516 27616 68572
rect 27616 68516 27672 68572
rect 27672 68516 27676 68572
rect 27612 68512 27676 68516
rect 27692 68572 27756 68576
rect 27692 68516 27696 68572
rect 27696 68516 27752 68572
rect 27752 68516 27756 68572
rect 27692 68512 27756 68516
rect 27772 68572 27836 68576
rect 27772 68516 27776 68572
rect 27776 68516 27832 68572
rect 27832 68516 27836 68572
rect 27772 68512 27836 68516
rect 27852 68572 27916 68576
rect 27852 68516 27856 68572
rect 27856 68516 27912 68572
rect 27912 68516 27916 68572
rect 27852 68512 27916 68516
rect 32612 68572 32676 68576
rect 32612 68516 32616 68572
rect 32616 68516 32672 68572
rect 32672 68516 32676 68572
rect 32612 68512 32676 68516
rect 32692 68572 32756 68576
rect 32692 68516 32696 68572
rect 32696 68516 32752 68572
rect 32752 68516 32756 68572
rect 32692 68512 32756 68516
rect 32772 68572 32836 68576
rect 32772 68516 32776 68572
rect 32776 68516 32832 68572
rect 32832 68516 32836 68572
rect 32772 68512 32836 68516
rect 32852 68572 32916 68576
rect 32852 68516 32856 68572
rect 32856 68516 32912 68572
rect 32912 68516 32916 68572
rect 32852 68512 32916 68516
rect 37612 68572 37676 68576
rect 37612 68516 37616 68572
rect 37616 68516 37672 68572
rect 37672 68516 37676 68572
rect 37612 68512 37676 68516
rect 37692 68572 37756 68576
rect 37692 68516 37696 68572
rect 37696 68516 37752 68572
rect 37752 68516 37756 68572
rect 37692 68512 37756 68516
rect 37772 68572 37836 68576
rect 37772 68516 37776 68572
rect 37776 68516 37832 68572
rect 37832 68516 37836 68572
rect 37772 68512 37836 68516
rect 37852 68572 37916 68576
rect 37852 68516 37856 68572
rect 37856 68516 37912 68572
rect 37912 68516 37916 68572
rect 37852 68512 37916 68516
rect 1952 68028 2016 68032
rect 1952 67972 1956 68028
rect 1956 67972 2012 68028
rect 2012 67972 2016 68028
rect 1952 67968 2016 67972
rect 2032 68028 2096 68032
rect 2032 67972 2036 68028
rect 2036 67972 2092 68028
rect 2092 67972 2096 68028
rect 2032 67968 2096 67972
rect 2112 68028 2176 68032
rect 2112 67972 2116 68028
rect 2116 67972 2172 68028
rect 2172 67972 2176 68028
rect 2112 67968 2176 67972
rect 2192 68028 2256 68032
rect 2192 67972 2196 68028
rect 2196 67972 2252 68028
rect 2252 67972 2256 68028
rect 2192 67968 2256 67972
rect 6952 68028 7016 68032
rect 6952 67972 6956 68028
rect 6956 67972 7012 68028
rect 7012 67972 7016 68028
rect 6952 67968 7016 67972
rect 7032 68028 7096 68032
rect 7032 67972 7036 68028
rect 7036 67972 7092 68028
rect 7092 67972 7096 68028
rect 7032 67968 7096 67972
rect 7112 68028 7176 68032
rect 7112 67972 7116 68028
rect 7116 67972 7172 68028
rect 7172 67972 7176 68028
rect 7112 67968 7176 67972
rect 7192 68028 7256 68032
rect 7192 67972 7196 68028
rect 7196 67972 7252 68028
rect 7252 67972 7256 68028
rect 7192 67968 7256 67972
rect 11952 68028 12016 68032
rect 11952 67972 11956 68028
rect 11956 67972 12012 68028
rect 12012 67972 12016 68028
rect 11952 67968 12016 67972
rect 12032 68028 12096 68032
rect 12032 67972 12036 68028
rect 12036 67972 12092 68028
rect 12092 67972 12096 68028
rect 12032 67968 12096 67972
rect 12112 68028 12176 68032
rect 12112 67972 12116 68028
rect 12116 67972 12172 68028
rect 12172 67972 12176 68028
rect 12112 67968 12176 67972
rect 12192 68028 12256 68032
rect 12192 67972 12196 68028
rect 12196 67972 12252 68028
rect 12252 67972 12256 68028
rect 12192 67968 12256 67972
rect 16952 68028 17016 68032
rect 16952 67972 16956 68028
rect 16956 67972 17012 68028
rect 17012 67972 17016 68028
rect 16952 67968 17016 67972
rect 17032 68028 17096 68032
rect 17032 67972 17036 68028
rect 17036 67972 17092 68028
rect 17092 67972 17096 68028
rect 17032 67968 17096 67972
rect 17112 68028 17176 68032
rect 17112 67972 17116 68028
rect 17116 67972 17172 68028
rect 17172 67972 17176 68028
rect 17112 67968 17176 67972
rect 17192 68028 17256 68032
rect 17192 67972 17196 68028
rect 17196 67972 17252 68028
rect 17252 67972 17256 68028
rect 17192 67968 17256 67972
rect 21952 68028 22016 68032
rect 21952 67972 21956 68028
rect 21956 67972 22012 68028
rect 22012 67972 22016 68028
rect 21952 67968 22016 67972
rect 22032 68028 22096 68032
rect 22032 67972 22036 68028
rect 22036 67972 22092 68028
rect 22092 67972 22096 68028
rect 22032 67968 22096 67972
rect 22112 68028 22176 68032
rect 22112 67972 22116 68028
rect 22116 67972 22172 68028
rect 22172 67972 22176 68028
rect 22112 67968 22176 67972
rect 22192 68028 22256 68032
rect 22192 67972 22196 68028
rect 22196 67972 22252 68028
rect 22252 67972 22256 68028
rect 22192 67968 22256 67972
rect 26952 68028 27016 68032
rect 26952 67972 26956 68028
rect 26956 67972 27012 68028
rect 27012 67972 27016 68028
rect 26952 67968 27016 67972
rect 27032 68028 27096 68032
rect 27032 67972 27036 68028
rect 27036 67972 27092 68028
rect 27092 67972 27096 68028
rect 27032 67968 27096 67972
rect 27112 68028 27176 68032
rect 27112 67972 27116 68028
rect 27116 67972 27172 68028
rect 27172 67972 27176 68028
rect 27112 67968 27176 67972
rect 27192 68028 27256 68032
rect 27192 67972 27196 68028
rect 27196 67972 27252 68028
rect 27252 67972 27256 68028
rect 27192 67968 27256 67972
rect 31952 68028 32016 68032
rect 31952 67972 31956 68028
rect 31956 67972 32012 68028
rect 32012 67972 32016 68028
rect 31952 67968 32016 67972
rect 32032 68028 32096 68032
rect 32032 67972 32036 68028
rect 32036 67972 32092 68028
rect 32092 67972 32096 68028
rect 32032 67968 32096 67972
rect 32112 68028 32176 68032
rect 32112 67972 32116 68028
rect 32116 67972 32172 68028
rect 32172 67972 32176 68028
rect 32112 67968 32176 67972
rect 32192 68028 32256 68032
rect 32192 67972 32196 68028
rect 32196 67972 32252 68028
rect 32252 67972 32256 68028
rect 32192 67968 32256 67972
rect 36952 68028 37016 68032
rect 36952 67972 36956 68028
rect 36956 67972 37012 68028
rect 37012 67972 37016 68028
rect 36952 67968 37016 67972
rect 37032 68028 37096 68032
rect 37032 67972 37036 68028
rect 37036 67972 37092 68028
rect 37092 67972 37096 68028
rect 37032 67968 37096 67972
rect 37112 68028 37176 68032
rect 37112 67972 37116 68028
rect 37116 67972 37172 68028
rect 37172 67972 37176 68028
rect 37112 67968 37176 67972
rect 37192 68028 37256 68032
rect 37192 67972 37196 68028
rect 37196 67972 37252 68028
rect 37252 67972 37256 68028
rect 37192 67968 37256 67972
rect 31708 67628 31772 67692
rect 2612 67484 2676 67488
rect 2612 67428 2616 67484
rect 2616 67428 2672 67484
rect 2672 67428 2676 67484
rect 2612 67424 2676 67428
rect 2692 67484 2756 67488
rect 2692 67428 2696 67484
rect 2696 67428 2752 67484
rect 2752 67428 2756 67484
rect 2692 67424 2756 67428
rect 2772 67484 2836 67488
rect 2772 67428 2776 67484
rect 2776 67428 2832 67484
rect 2832 67428 2836 67484
rect 2772 67424 2836 67428
rect 2852 67484 2916 67488
rect 2852 67428 2856 67484
rect 2856 67428 2912 67484
rect 2912 67428 2916 67484
rect 2852 67424 2916 67428
rect 7612 67484 7676 67488
rect 7612 67428 7616 67484
rect 7616 67428 7672 67484
rect 7672 67428 7676 67484
rect 7612 67424 7676 67428
rect 7692 67484 7756 67488
rect 7692 67428 7696 67484
rect 7696 67428 7752 67484
rect 7752 67428 7756 67484
rect 7692 67424 7756 67428
rect 7772 67484 7836 67488
rect 7772 67428 7776 67484
rect 7776 67428 7832 67484
rect 7832 67428 7836 67484
rect 7772 67424 7836 67428
rect 7852 67484 7916 67488
rect 7852 67428 7856 67484
rect 7856 67428 7912 67484
rect 7912 67428 7916 67484
rect 7852 67424 7916 67428
rect 12612 67484 12676 67488
rect 12612 67428 12616 67484
rect 12616 67428 12672 67484
rect 12672 67428 12676 67484
rect 12612 67424 12676 67428
rect 12692 67484 12756 67488
rect 12692 67428 12696 67484
rect 12696 67428 12752 67484
rect 12752 67428 12756 67484
rect 12692 67424 12756 67428
rect 12772 67484 12836 67488
rect 12772 67428 12776 67484
rect 12776 67428 12832 67484
rect 12832 67428 12836 67484
rect 12772 67424 12836 67428
rect 12852 67484 12916 67488
rect 12852 67428 12856 67484
rect 12856 67428 12912 67484
rect 12912 67428 12916 67484
rect 12852 67424 12916 67428
rect 17612 67484 17676 67488
rect 17612 67428 17616 67484
rect 17616 67428 17672 67484
rect 17672 67428 17676 67484
rect 17612 67424 17676 67428
rect 17692 67484 17756 67488
rect 17692 67428 17696 67484
rect 17696 67428 17752 67484
rect 17752 67428 17756 67484
rect 17692 67424 17756 67428
rect 17772 67484 17836 67488
rect 17772 67428 17776 67484
rect 17776 67428 17832 67484
rect 17832 67428 17836 67484
rect 17772 67424 17836 67428
rect 17852 67484 17916 67488
rect 17852 67428 17856 67484
rect 17856 67428 17912 67484
rect 17912 67428 17916 67484
rect 17852 67424 17916 67428
rect 22612 67484 22676 67488
rect 22612 67428 22616 67484
rect 22616 67428 22672 67484
rect 22672 67428 22676 67484
rect 22612 67424 22676 67428
rect 22692 67484 22756 67488
rect 22692 67428 22696 67484
rect 22696 67428 22752 67484
rect 22752 67428 22756 67484
rect 22692 67424 22756 67428
rect 22772 67484 22836 67488
rect 22772 67428 22776 67484
rect 22776 67428 22832 67484
rect 22832 67428 22836 67484
rect 22772 67424 22836 67428
rect 22852 67484 22916 67488
rect 22852 67428 22856 67484
rect 22856 67428 22912 67484
rect 22912 67428 22916 67484
rect 22852 67424 22916 67428
rect 27612 67484 27676 67488
rect 27612 67428 27616 67484
rect 27616 67428 27672 67484
rect 27672 67428 27676 67484
rect 27612 67424 27676 67428
rect 27692 67484 27756 67488
rect 27692 67428 27696 67484
rect 27696 67428 27752 67484
rect 27752 67428 27756 67484
rect 27692 67424 27756 67428
rect 27772 67484 27836 67488
rect 27772 67428 27776 67484
rect 27776 67428 27832 67484
rect 27832 67428 27836 67484
rect 27772 67424 27836 67428
rect 27852 67484 27916 67488
rect 27852 67428 27856 67484
rect 27856 67428 27912 67484
rect 27912 67428 27916 67484
rect 27852 67424 27916 67428
rect 32612 67484 32676 67488
rect 32612 67428 32616 67484
rect 32616 67428 32672 67484
rect 32672 67428 32676 67484
rect 32612 67424 32676 67428
rect 32692 67484 32756 67488
rect 32692 67428 32696 67484
rect 32696 67428 32752 67484
rect 32752 67428 32756 67484
rect 32692 67424 32756 67428
rect 32772 67484 32836 67488
rect 32772 67428 32776 67484
rect 32776 67428 32832 67484
rect 32832 67428 32836 67484
rect 32772 67424 32836 67428
rect 32852 67484 32916 67488
rect 32852 67428 32856 67484
rect 32856 67428 32912 67484
rect 32912 67428 32916 67484
rect 32852 67424 32916 67428
rect 37612 67484 37676 67488
rect 37612 67428 37616 67484
rect 37616 67428 37672 67484
rect 37672 67428 37676 67484
rect 37612 67424 37676 67428
rect 37692 67484 37756 67488
rect 37692 67428 37696 67484
rect 37696 67428 37752 67484
rect 37752 67428 37756 67484
rect 37692 67424 37756 67428
rect 37772 67484 37836 67488
rect 37772 67428 37776 67484
rect 37776 67428 37832 67484
rect 37832 67428 37836 67484
rect 37772 67424 37836 67428
rect 37852 67484 37916 67488
rect 37852 67428 37856 67484
rect 37856 67428 37912 67484
rect 37912 67428 37916 67484
rect 37852 67424 37916 67428
rect 1952 66940 2016 66944
rect 1952 66884 1956 66940
rect 1956 66884 2012 66940
rect 2012 66884 2016 66940
rect 1952 66880 2016 66884
rect 2032 66940 2096 66944
rect 2032 66884 2036 66940
rect 2036 66884 2092 66940
rect 2092 66884 2096 66940
rect 2032 66880 2096 66884
rect 2112 66940 2176 66944
rect 2112 66884 2116 66940
rect 2116 66884 2172 66940
rect 2172 66884 2176 66940
rect 2112 66880 2176 66884
rect 2192 66940 2256 66944
rect 2192 66884 2196 66940
rect 2196 66884 2252 66940
rect 2252 66884 2256 66940
rect 2192 66880 2256 66884
rect 6952 66940 7016 66944
rect 6952 66884 6956 66940
rect 6956 66884 7012 66940
rect 7012 66884 7016 66940
rect 6952 66880 7016 66884
rect 7032 66940 7096 66944
rect 7032 66884 7036 66940
rect 7036 66884 7092 66940
rect 7092 66884 7096 66940
rect 7032 66880 7096 66884
rect 7112 66940 7176 66944
rect 7112 66884 7116 66940
rect 7116 66884 7172 66940
rect 7172 66884 7176 66940
rect 7112 66880 7176 66884
rect 7192 66940 7256 66944
rect 7192 66884 7196 66940
rect 7196 66884 7252 66940
rect 7252 66884 7256 66940
rect 7192 66880 7256 66884
rect 11952 66940 12016 66944
rect 11952 66884 11956 66940
rect 11956 66884 12012 66940
rect 12012 66884 12016 66940
rect 11952 66880 12016 66884
rect 12032 66940 12096 66944
rect 12032 66884 12036 66940
rect 12036 66884 12092 66940
rect 12092 66884 12096 66940
rect 12032 66880 12096 66884
rect 12112 66940 12176 66944
rect 12112 66884 12116 66940
rect 12116 66884 12172 66940
rect 12172 66884 12176 66940
rect 12112 66880 12176 66884
rect 12192 66940 12256 66944
rect 12192 66884 12196 66940
rect 12196 66884 12252 66940
rect 12252 66884 12256 66940
rect 12192 66880 12256 66884
rect 16952 66940 17016 66944
rect 16952 66884 16956 66940
rect 16956 66884 17012 66940
rect 17012 66884 17016 66940
rect 16952 66880 17016 66884
rect 17032 66940 17096 66944
rect 17032 66884 17036 66940
rect 17036 66884 17092 66940
rect 17092 66884 17096 66940
rect 17032 66880 17096 66884
rect 17112 66940 17176 66944
rect 17112 66884 17116 66940
rect 17116 66884 17172 66940
rect 17172 66884 17176 66940
rect 17112 66880 17176 66884
rect 17192 66940 17256 66944
rect 17192 66884 17196 66940
rect 17196 66884 17252 66940
rect 17252 66884 17256 66940
rect 17192 66880 17256 66884
rect 21952 66940 22016 66944
rect 21952 66884 21956 66940
rect 21956 66884 22012 66940
rect 22012 66884 22016 66940
rect 21952 66880 22016 66884
rect 22032 66940 22096 66944
rect 22032 66884 22036 66940
rect 22036 66884 22092 66940
rect 22092 66884 22096 66940
rect 22032 66880 22096 66884
rect 22112 66940 22176 66944
rect 22112 66884 22116 66940
rect 22116 66884 22172 66940
rect 22172 66884 22176 66940
rect 22112 66880 22176 66884
rect 22192 66940 22256 66944
rect 22192 66884 22196 66940
rect 22196 66884 22252 66940
rect 22252 66884 22256 66940
rect 22192 66880 22256 66884
rect 26952 66940 27016 66944
rect 26952 66884 26956 66940
rect 26956 66884 27012 66940
rect 27012 66884 27016 66940
rect 26952 66880 27016 66884
rect 27032 66940 27096 66944
rect 27032 66884 27036 66940
rect 27036 66884 27092 66940
rect 27092 66884 27096 66940
rect 27032 66880 27096 66884
rect 27112 66940 27176 66944
rect 27112 66884 27116 66940
rect 27116 66884 27172 66940
rect 27172 66884 27176 66940
rect 27112 66880 27176 66884
rect 27192 66940 27256 66944
rect 27192 66884 27196 66940
rect 27196 66884 27252 66940
rect 27252 66884 27256 66940
rect 27192 66880 27256 66884
rect 31952 66940 32016 66944
rect 31952 66884 31956 66940
rect 31956 66884 32012 66940
rect 32012 66884 32016 66940
rect 31952 66880 32016 66884
rect 32032 66940 32096 66944
rect 32032 66884 32036 66940
rect 32036 66884 32092 66940
rect 32092 66884 32096 66940
rect 32032 66880 32096 66884
rect 32112 66940 32176 66944
rect 32112 66884 32116 66940
rect 32116 66884 32172 66940
rect 32172 66884 32176 66940
rect 32112 66880 32176 66884
rect 32192 66940 32256 66944
rect 32192 66884 32196 66940
rect 32196 66884 32252 66940
rect 32252 66884 32256 66940
rect 32192 66880 32256 66884
rect 36952 66940 37016 66944
rect 36952 66884 36956 66940
rect 36956 66884 37012 66940
rect 37012 66884 37016 66940
rect 36952 66880 37016 66884
rect 37032 66940 37096 66944
rect 37032 66884 37036 66940
rect 37036 66884 37092 66940
rect 37092 66884 37096 66940
rect 37032 66880 37096 66884
rect 37112 66940 37176 66944
rect 37112 66884 37116 66940
rect 37116 66884 37172 66940
rect 37172 66884 37176 66940
rect 37112 66880 37176 66884
rect 37192 66940 37256 66944
rect 37192 66884 37196 66940
rect 37196 66884 37252 66940
rect 37252 66884 37256 66940
rect 37192 66880 37256 66884
rect 2612 66396 2676 66400
rect 2612 66340 2616 66396
rect 2616 66340 2672 66396
rect 2672 66340 2676 66396
rect 2612 66336 2676 66340
rect 2692 66396 2756 66400
rect 2692 66340 2696 66396
rect 2696 66340 2752 66396
rect 2752 66340 2756 66396
rect 2692 66336 2756 66340
rect 2772 66396 2836 66400
rect 2772 66340 2776 66396
rect 2776 66340 2832 66396
rect 2832 66340 2836 66396
rect 2772 66336 2836 66340
rect 2852 66396 2916 66400
rect 2852 66340 2856 66396
rect 2856 66340 2912 66396
rect 2912 66340 2916 66396
rect 2852 66336 2916 66340
rect 7612 66396 7676 66400
rect 7612 66340 7616 66396
rect 7616 66340 7672 66396
rect 7672 66340 7676 66396
rect 7612 66336 7676 66340
rect 7692 66396 7756 66400
rect 7692 66340 7696 66396
rect 7696 66340 7752 66396
rect 7752 66340 7756 66396
rect 7692 66336 7756 66340
rect 7772 66396 7836 66400
rect 7772 66340 7776 66396
rect 7776 66340 7832 66396
rect 7832 66340 7836 66396
rect 7772 66336 7836 66340
rect 7852 66396 7916 66400
rect 7852 66340 7856 66396
rect 7856 66340 7912 66396
rect 7912 66340 7916 66396
rect 7852 66336 7916 66340
rect 12612 66396 12676 66400
rect 12612 66340 12616 66396
rect 12616 66340 12672 66396
rect 12672 66340 12676 66396
rect 12612 66336 12676 66340
rect 12692 66396 12756 66400
rect 12692 66340 12696 66396
rect 12696 66340 12752 66396
rect 12752 66340 12756 66396
rect 12692 66336 12756 66340
rect 12772 66396 12836 66400
rect 12772 66340 12776 66396
rect 12776 66340 12832 66396
rect 12832 66340 12836 66396
rect 12772 66336 12836 66340
rect 12852 66396 12916 66400
rect 12852 66340 12856 66396
rect 12856 66340 12912 66396
rect 12912 66340 12916 66396
rect 12852 66336 12916 66340
rect 17612 66396 17676 66400
rect 17612 66340 17616 66396
rect 17616 66340 17672 66396
rect 17672 66340 17676 66396
rect 17612 66336 17676 66340
rect 17692 66396 17756 66400
rect 17692 66340 17696 66396
rect 17696 66340 17752 66396
rect 17752 66340 17756 66396
rect 17692 66336 17756 66340
rect 17772 66396 17836 66400
rect 17772 66340 17776 66396
rect 17776 66340 17832 66396
rect 17832 66340 17836 66396
rect 17772 66336 17836 66340
rect 17852 66396 17916 66400
rect 17852 66340 17856 66396
rect 17856 66340 17912 66396
rect 17912 66340 17916 66396
rect 17852 66336 17916 66340
rect 22612 66396 22676 66400
rect 22612 66340 22616 66396
rect 22616 66340 22672 66396
rect 22672 66340 22676 66396
rect 22612 66336 22676 66340
rect 22692 66396 22756 66400
rect 22692 66340 22696 66396
rect 22696 66340 22752 66396
rect 22752 66340 22756 66396
rect 22692 66336 22756 66340
rect 22772 66396 22836 66400
rect 22772 66340 22776 66396
rect 22776 66340 22832 66396
rect 22832 66340 22836 66396
rect 22772 66336 22836 66340
rect 22852 66396 22916 66400
rect 22852 66340 22856 66396
rect 22856 66340 22912 66396
rect 22912 66340 22916 66396
rect 22852 66336 22916 66340
rect 27612 66396 27676 66400
rect 27612 66340 27616 66396
rect 27616 66340 27672 66396
rect 27672 66340 27676 66396
rect 27612 66336 27676 66340
rect 27692 66396 27756 66400
rect 27692 66340 27696 66396
rect 27696 66340 27752 66396
rect 27752 66340 27756 66396
rect 27692 66336 27756 66340
rect 27772 66396 27836 66400
rect 27772 66340 27776 66396
rect 27776 66340 27832 66396
rect 27832 66340 27836 66396
rect 27772 66336 27836 66340
rect 27852 66396 27916 66400
rect 27852 66340 27856 66396
rect 27856 66340 27912 66396
rect 27912 66340 27916 66396
rect 27852 66336 27916 66340
rect 32612 66396 32676 66400
rect 32612 66340 32616 66396
rect 32616 66340 32672 66396
rect 32672 66340 32676 66396
rect 32612 66336 32676 66340
rect 32692 66396 32756 66400
rect 32692 66340 32696 66396
rect 32696 66340 32752 66396
rect 32752 66340 32756 66396
rect 32692 66336 32756 66340
rect 32772 66396 32836 66400
rect 32772 66340 32776 66396
rect 32776 66340 32832 66396
rect 32832 66340 32836 66396
rect 32772 66336 32836 66340
rect 32852 66396 32916 66400
rect 32852 66340 32856 66396
rect 32856 66340 32912 66396
rect 32912 66340 32916 66396
rect 32852 66336 32916 66340
rect 37612 66396 37676 66400
rect 37612 66340 37616 66396
rect 37616 66340 37672 66396
rect 37672 66340 37676 66396
rect 37612 66336 37676 66340
rect 37692 66396 37756 66400
rect 37692 66340 37696 66396
rect 37696 66340 37752 66396
rect 37752 66340 37756 66396
rect 37692 66336 37756 66340
rect 37772 66396 37836 66400
rect 37772 66340 37776 66396
rect 37776 66340 37832 66396
rect 37832 66340 37836 66396
rect 37772 66336 37836 66340
rect 37852 66396 37916 66400
rect 37852 66340 37856 66396
rect 37856 66340 37912 66396
rect 37912 66340 37916 66396
rect 37852 66336 37916 66340
rect 1952 65852 2016 65856
rect 1952 65796 1956 65852
rect 1956 65796 2012 65852
rect 2012 65796 2016 65852
rect 1952 65792 2016 65796
rect 2032 65852 2096 65856
rect 2032 65796 2036 65852
rect 2036 65796 2092 65852
rect 2092 65796 2096 65852
rect 2032 65792 2096 65796
rect 2112 65852 2176 65856
rect 2112 65796 2116 65852
rect 2116 65796 2172 65852
rect 2172 65796 2176 65852
rect 2112 65792 2176 65796
rect 2192 65852 2256 65856
rect 2192 65796 2196 65852
rect 2196 65796 2252 65852
rect 2252 65796 2256 65852
rect 2192 65792 2256 65796
rect 6952 65852 7016 65856
rect 6952 65796 6956 65852
rect 6956 65796 7012 65852
rect 7012 65796 7016 65852
rect 6952 65792 7016 65796
rect 7032 65852 7096 65856
rect 7032 65796 7036 65852
rect 7036 65796 7092 65852
rect 7092 65796 7096 65852
rect 7032 65792 7096 65796
rect 7112 65852 7176 65856
rect 7112 65796 7116 65852
rect 7116 65796 7172 65852
rect 7172 65796 7176 65852
rect 7112 65792 7176 65796
rect 7192 65852 7256 65856
rect 7192 65796 7196 65852
rect 7196 65796 7252 65852
rect 7252 65796 7256 65852
rect 7192 65792 7256 65796
rect 11952 65852 12016 65856
rect 11952 65796 11956 65852
rect 11956 65796 12012 65852
rect 12012 65796 12016 65852
rect 11952 65792 12016 65796
rect 12032 65852 12096 65856
rect 12032 65796 12036 65852
rect 12036 65796 12092 65852
rect 12092 65796 12096 65852
rect 12032 65792 12096 65796
rect 12112 65852 12176 65856
rect 12112 65796 12116 65852
rect 12116 65796 12172 65852
rect 12172 65796 12176 65852
rect 12112 65792 12176 65796
rect 12192 65852 12256 65856
rect 12192 65796 12196 65852
rect 12196 65796 12252 65852
rect 12252 65796 12256 65852
rect 12192 65792 12256 65796
rect 16952 65852 17016 65856
rect 16952 65796 16956 65852
rect 16956 65796 17012 65852
rect 17012 65796 17016 65852
rect 16952 65792 17016 65796
rect 17032 65852 17096 65856
rect 17032 65796 17036 65852
rect 17036 65796 17092 65852
rect 17092 65796 17096 65852
rect 17032 65792 17096 65796
rect 17112 65852 17176 65856
rect 17112 65796 17116 65852
rect 17116 65796 17172 65852
rect 17172 65796 17176 65852
rect 17112 65792 17176 65796
rect 17192 65852 17256 65856
rect 17192 65796 17196 65852
rect 17196 65796 17252 65852
rect 17252 65796 17256 65852
rect 17192 65792 17256 65796
rect 21952 65852 22016 65856
rect 21952 65796 21956 65852
rect 21956 65796 22012 65852
rect 22012 65796 22016 65852
rect 21952 65792 22016 65796
rect 22032 65852 22096 65856
rect 22032 65796 22036 65852
rect 22036 65796 22092 65852
rect 22092 65796 22096 65852
rect 22032 65792 22096 65796
rect 22112 65852 22176 65856
rect 22112 65796 22116 65852
rect 22116 65796 22172 65852
rect 22172 65796 22176 65852
rect 22112 65792 22176 65796
rect 22192 65852 22256 65856
rect 22192 65796 22196 65852
rect 22196 65796 22252 65852
rect 22252 65796 22256 65852
rect 22192 65792 22256 65796
rect 26952 65852 27016 65856
rect 26952 65796 26956 65852
rect 26956 65796 27012 65852
rect 27012 65796 27016 65852
rect 26952 65792 27016 65796
rect 27032 65852 27096 65856
rect 27032 65796 27036 65852
rect 27036 65796 27092 65852
rect 27092 65796 27096 65852
rect 27032 65792 27096 65796
rect 27112 65852 27176 65856
rect 27112 65796 27116 65852
rect 27116 65796 27172 65852
rect 27172 65796 27176 65852
rect 27112 65792 27176 65796
rect 27192 65852 27256 65856
rect 27192 65796 27196 65852
rect 27196 65796 27252 65852
rect 27252 65796 27256 65852
rect 27192 65792 27256 65796
rect 31952 65852 32016 65856
rect 31952 65796 31956 65852
rect 31956 65796 32012 65852
rect 32012 65796 32016 65852
rect 31952 65792 32016 65796
rect 32032 65852 32096 65856
rect 32032 65796 32036 65852
rect 32036 65796 32092 65852
rect 32092 65796 32096 65852
rect 32032 65792 32096 65796
rect 32112 65852 32176 65856
rect 32112 65796 32116 65852
rect 32116 65796 32172 65852
rect 32172 65796 32176 65852
rect 32112 65792 32176 65796
rect 32192 65852 32256 65856
rect 32192 65796 32196 65852
rect 32196 65796 32252 65852
rect 32252 65796 32256 65852
rect 32192 65792 32256 65796
rect 36952 65852 37016 65856
rect 36952 65796 36956 65852
rect 36956 65796 37012 65852
rect 37012 65796 37016 65852
rect 36952 65792 37016 65796
rect 37032 65852 37096 65856
rect 37032 65796 37036 65852
rect 37036 65796 37092 65852
rect 37092 65796 37096 65852
rect 37032 65792 37096 65796
rect 37112 65852 37176 65856
rect 37112 65796 37116 65852
rect 37116 65796 37172 65852
rect 37172 65796 37176 65852
rect 37112 65792 37176 65796
rect 37192 65852 37256 65856
rect 37192 65796 37196 65852
rect 37196 65796 37252 65852
rect 37252 65796 37256 65852
rect 37192 65792 37256 65796
rect 2612 65308 2676 65312
rect 2612 65252 2616 65308
rect 2616 65252 2672 65308
rect 2672 65252 2676 65308
rect 2612 65248 2676 65252
rect 2692 65308 2756 65312
rect 2692 65252 2696 65308
rect 2696 65252 2752 65308
rect 2752 65252 2756 65308
rect 2692 65248 2756 65252
rect 2772 65308 2836 65312
rect 2772 65252 2776 65308
rect 2776 65252 2832 65308
rect 2832 65252 2836 65308
rect 2772 65248 2836 65252
rect 2852 65308 2916 65312
rect 2852 65252 2856 65308
rect 2856 65252 2912 65308
rect 2912 65252 2916 65308
rect 2852 65248 2916 65252
rect 7612 65308 7676 65312
rect 7612 65252 7616 65308
rect 7616 65252 7672 65308
rect 7672 65252 7676 65308
rect 7612 65248 7676 65252
rect 7692 65308 7756 65312
rect 7692 65252 7696 65308
rect 7696 65252 7752 65308
rect 7752 65252 7756 65308
rect 7692 65248 7756 65252
rect 7772 65308 7836 65312
rect 7772 65252 7776 65308
rect 7776 65252 7832 65308
rect 7832 65252 7836 65308
rect 7772 65248 7836 65252
rect 7852 65308 7916 65312
rect 7852 65252 7856 65308
rect 7856 65252 7912 65308
rect 7912 65252 7916 65308
rect 7852 65248 7916 65252
rect 12612 65308 12676 65312
rect 12612 65252 12616 65308
rect 12616 65252 12672 65308
rect 12672 65252 12676 65308
rect 12612 65248 12676 65252
rect 12692 65308 12756 65312
rect 12692 65252 12696 65308
rect 12696 65252 12752 65308
rect 12752 65252 12756 65308
rect 12692 65248 12756 65252
rect 12772 65308 12836 65312
rect 12772 65252 12776 65308
rect 12776 65252 12832 65308
rect 12832 65252 12836 65308
rect 12772 65248 12836 65252
rect 12852 65308 12916 65312
rect 12852 65252 12856 65308
rect 12856 65252 12912 65308
rect 12912 65252 12916 65308
rect 12852 65248 12916 65252
rect 17612 65308 17676 65312
rect 17612 65252 17616 65308
rect 17616 65252 17672 65308
rect 17672 65252 17676 65308
rect 17612 65248 17676 65252
rect 17692 65308 17756 65312
rect 17692 65252 17696 65308
rect 17696 65252 17752 65308
rect 17752 65252 17756 65308
rect 17692 65248 17756 65252
rect 17772 65308 17836 65312
rect 17772 65252 17776 65308
rect 17776 65252 17832 65308
rect 17832 65252 17836 65308
rect 17772 65248 17836 65252
rect 17852 65308 17916 65312
rect 17852 65252 17856 65308
rect 17856 65252 17912 65308
rect 17912 65252 17916 65308
rect 17852 65248 17916 65252
rect 22612 65308 22676 65312
rect 22612 65252 22616 65308
rect 22616 65252 22672 65308
rect 22672 65252 22676 65308
rect 22612 65248 22676 65252
rect 22692 65308 22756 65312
rect 22692 65252 22696 65308
rect 22696 65252 22752 65308
rect 22752 65252 22756 65308
rect 22692 65248 22756 65252
rect 22772 65308 22836 65312
rect 22772 65252 22776 65308
rect 22776 65252 22832 65308
rect 22832 65252 22836 65308
rect 22772 65248 22836 65252
rect 22852 65308 22916 65312
rect 22852 65252 22856 65308
rect 22856 65252 22912 65308
rect 22912 65252 22916 65308
rect 22852 65248 22916 65252
rect 27612 65308 27676 65312
rect 27612 65252 27616 65308
rect 27616 65252 27672 65308
rect 27672 65252 27676 65308
rect 27612 65248 27676 65252
rect 27692 65308 27756 65312
rect 27692 65252 27696 65308
rect 27696 65252 27752 65308
rect 27752 65252 27756 65308
rect 27692 65248 27756 65252
rect 27772 65308 27836 65312
rect 27772 65252 27776 65308
rect 27776 65252 27832 65308
rect 27832 65252 27836 65308
rect 27772 65248 27836 65252
rect 27852 65308 27916 65312
rect 27852 65252 27856 65308
rect 27856 65252 27912 65308
rect 27912 65252 27916 65308
rect 27852 65248 27916 65252
rect 32612 65308 32676 65312
rect 32612 65252 32616 65308
rect 32616 65252 32672 65308
rect 32672 65252 32676 65308
rect 32612 65248 32676 65252
rect 32692 65308 32756 65312
rect 32692 65252 32696 65308
rect 32696 65252 32752 65308
rect 32752 65252 32756 65308
rect 32692 65248 32756 65252
rect 32772 65308 32836 65312
rect 32772 65252 32776 65308
rect 32776 65252 32832 65308
rect 32832 65252 32836 65308
rect 32772 65248 32836 65252
rect 32852 65308 32916 65312
rect 32852 65252 32856 65308
rect 32856 65252 32912 65308
rect 32912 65252 32916 65308
rect 32852 65248 32916 65252
rect 37612 65308 37676 65312
rect 37612 65252 37616 65308
rect 37616 65252 37672 65308
rect 37672 65252 37676 65308
rect 37612 65248 37676 65252
rect 37692 65308 37756 65312
rect 37692 65252 37696 65308
rect 37696 65252 37752 65308
rect 37752 65252 37756 65308
rect 37692 65248 37756 65252
rect 37772 65308 37836 65312
rect 37772 65252 37776 65308
rect 37776 65252 37832 65308
rect 37832 65252 37836 65308
rect 37772 65248 37836 65252
rect 37852 65308 37916 65312
rect 37852 65252 37856 65308
rect 37856 65252 37912 65308
rect 37912 65252 37916 65308
rect 37852 65248 37916 65252
rect 1952 64764 2016 64768
rect 1952 64708 1956 64764
rect 1956 64708 2012 64764
rect 2012 64708 2016 64764
rect 1952 64704 2016 64708
rect 2032 64764 2096 64768
rect 2032 64708 2036 64764
rect 2036 64708 2092 64764
rect 2092 64708 2096 64764
rect 2032 64704 2096 64708
rect 2112 64764 2176 64768
rect 2112 64708 2116 64764
rect 2116 64708 2172 64764
rect 2172 64708 2176 64764
rect 2112 64704 2176 64708
rect 2192 64764 2256 64768
rect 2192 64708 2196 64764
rect 2196 64708 2252 64764
rect 2252 64708 2256 64764
rect 2192 64704 2256 64708
rect 6952 64764 7016 64768
rect 6952 64708 6956 64764
rect 6956 64708 7012 64764
rect 7012 64708 7016 64764
rect 6952 64704 7016 64708
rect 7032 64764 7096 64768
rect 7032 64708 7036 64764
rect 7036 64708 7092 64764
rect 7092 64708 7096 64764
rect 7032 64704 7096 64708
rect 7112 64764 7176 64768
rect 7112 64708 7116 64764
rect 7116 64708 7172 64764
rect 7172 64708 7176 64764
rect 7112 64704 7176 64708
rect 7192 64764 7256 64768
rect 7192 64708 7196 64764
rect 7196 64708 7252 64764
rect 7252 64708 7256 64764
rect 7192 64704 7256 64708
rect 11952 64764 12016 64768
rect 11952 64708 11956 64764
rect 11956 64708 12012 64764
rect 12012 64708 12016 64764
rect 11952 64704 12016 64708
rect 12032 64764 12096 64768
rect 12032 64708 12036 64764
rect 12036 64708 12092 64764
rect 12092 64708 12096 64764
rect 12032 64704 12096 64708
rect 12112 64764 12176 64768
rect 12112 64708 12116 64764
rect 12116 64708 12172 64764
rect 12172 64708 12176 64764
rect 12112 64704 12176 64708
rect 12192 64764 12256 64768
rect 12192 64708 12196 64764
rect 12196 64708 12252 64764
rect 12252 64708 12256 64764
rect 12192 64704 12256 64708
rect 16952 64764 17016 64768
rect 16952 64708 16956 64764
rect 16956 64708 17012 64764
rect 17012 64708 17016 64764
rect 16952 64704 17016 64708
rect 17032 64764 17096 64768
rect 17032 64708 17036 64764
rect 17036 64708 17092 64764
rect 17092 64708 17096 64764
rect 17032 64704 17096 64708
rect 17112 64764 17176 64768
rect 17112 64708 17116 64764
rect 17116 64708 17172 64764
rect 17172 64708 17176 64764
rect 17112 64704 17176 64708
rect 17192 64764 17256 64768
rect 17192 64708 17196 64764
rect 17196 64708 17252 64764
rect 17252 64708 17256 64764
rect 17192 64704 17256 64708
rect 21952 64764 22016 64768
rect 21952 64708 21956 64764
rect 21956 64708 22012 64764
rect 22012 64708 22016 64764
rect 21952 64704 22016 64708
rect 22032 64764 22096 64768
rect 22032 64708 22036 64764
rect 22036 64708 22092 64764
rect 22092 64708 22096 64764
rect 22032 64704 22096 64708
rect 22112 64764 22176 64768
rect 22112 64708 22116 64764
rect 22116 64708 22172 64764
rect 22172 64708 22176 64764
rect 22112 64704 22176 64708
rect 22192 64764 22256 64768
rect 22192 64708 22196 64764
rect 22196 64708 22252 64764
rect 22252 64708 22256 64764
rect 22192 64704 22256 64708
rect 26952 64764 27016 64768
rect 26952 64708 26956 64764
rect 26956 64708 27012 64764
rect 27012 64708 27016 64764
rect 26952 64704 27016 64708
rect 27032 64764 27096 64768
rect 27032 64708 27036 64764
rect 27036 64708 27092 64764
rect 27092 64708 27096 64764
rect 27032 64704 27096 64708
rect 27112 64764 27176 64768
rect 27112 64708 27116 64764
rect 27116 64708 27172 64764
rect 27172 64708 27176 64764
rect 27112 64704 27176 64708
rect 27192 64764 27256 64768
rect 27192 64708 27196 64764
rect 27196 64708 27252 64764
rect 27252 64708 27256 64764
rect 27192 64704 27256 64708
rect 31952 64764 32016 64768
rect 31952 64708 31956 64764
rect 31956 64708 32012 64764
rect 32012 64708 32016 64764
rect 31952 64704 32016 64708
rect 32032 64764 32096 64768
rect 32032 64708 32036 64764
rect 32036 64708 32092 64764
rect 32092 64708 32096 64764
rect 32032 64704 32096 64708
rect 32112 64764 32176 64768
rect 32112 64708 32116 64764
rect 32116 64708 32172 64764
rect 32172 64708 32176 64764
rect 32112 64704 32176 64708
rect 32192 64764 32256 64768
rect 32192 64708 32196 64764
rect 32196 64708 32252 64764
rect 32252 64708 32256 64764
rect 32192 64704 32256 64708
rect 36952 64764 37016 64768
rect 36952 64708 36956 64764
rect 36956 64708 37012 64764
rect 37012 64708 37016 64764
rect 36952 64704 37016 64708
rect 37032 64764 37096 64768
rect 37032 64708 37036 64764
rect 37036 64708 37092 64764
rect 37092 64708 37096 64764
rect 37032 64704 37096 64708
rect 37112 64764 37176 64768
rect 37112 64708 37116 64764
rect 37116 64708 37172 64764
rect 37172 64708 37176 64764
rect 37112 64704 37176 64708
rect 37192 64764 37256 64768
rect 37192 64708 37196 64764
rect 37196 64708 37252 64764
rect 37252 64708 37256 64764
rect 37192 64704 37256 64708
rect 2612 64220 2676 64224
rect 2612 64164 2616 64220
rect 2616 64164 2672 64220
rect 2672 64164 2676 64220
rect 2612 64160 2676 64164
rect 2692 64220 2756 64224
rect 2692 64164 2696 64220
rect 2696 64164 2752 64220
rect 2752 64164 2756 64220
rect 2692 64160 2756 64164
rect 2772 64220 2836 64224
rect 2772 64164 2776 64220
rect 2776 64164 2832 64220
rect 2832 64164 2836 64220
rect 2772 64160 2836 64164
rect 2852 64220 2916 64224
rect 2852 64164 2856 64220
rect 2856 64164 2912 64220
rect 2912 64164 2916 64220
rect 2852 64160 2916 64164
rect 7612 64220 7676 64224
rect 7612 64164 7616 64220
rect 7616 64164 7672 64220
rect 7672 64164 7676 64220
rect 7612 64160 7676 64164
rect 7692 64220 7756 64224
rect 7692 64164 7696 64220
rect 7696 64164 7752 64220
rect 7752 64164 7756 64220
rect 7692 64160 7756 64164
rect 7772 64220 7836 64224
rect 7772 64164 7776 64220
rect 7776 64164 7832 64220
rect 7832 64164 7836 64220
rect 7772 64160 7836 64164
rect 7852 64220 7916 64224
rect 7852 64164 7856 64220
rect 7856 64164 7912 64220
rect 7912 64164 7916 64220
rect 7852 64160 7916 64164
rect 12612 64220 12676 64224
rect 12612 64164 12616 64220
rect 12616 64164 12672 64220
rect 12672 64164 12676 64220
rect 12612 64160 12676 64164
rect 12692 64220 12756 64224
rect 12692 64164 12696 64220
rect 12696 64164 12752 64220
rect 12752 64164 12756 64220
rect 12692 64160 12756 64164
rect 12772 64220 12836 64224
rect 12772 64164 12776 64220
rect 12776 64164 12832 64220
rect 12832 64164 12836 64220
rect 12772 64160 12836 64164
rect 12852 64220 12916 64224
rect 12852 64164 12856 64220
rect 12856 64164 12912 64220
rect 12912 64164 12916 64220
rect 12852 64160 12916 64164
rect 17612 64220 17676 64224
rect 17612 64164 17616 64220
rect 17616 64164 17672 64220
rect 17672 64164 17676 64220
rect 17612 64160 17676 64164
rect 17692 64220 17756 64224
rect 17692 64164 17696 64220
rect 17696 64164 17752 64220
rect 17752 64164 17756 64220
rect 17692 64160 17756 64164
rect 17772 64220 17836 64224
rect 17772 64164 17776 64220
rect 17776 64164 17832 64220
rect 17832 64164 17836 64220
rect 17772 64160 17836 64164
rect 17852 64220 17916 64224
rect 17852 64164 17856 64220
rect 17856 64164 17912 64220
rect 17912 64164 17916 64220
rect 17852 64160 17916 64164
rect 22612 64220 22676 64224
rect 22612 64164 22616 64220
rect 22616 64164 22672 64220
rect 22672 64164 22676 64220
rect 22612 64160 22676 64164
rect 22692 64220 22756 64224
rect 22692 64164 22696 64220
rect 22696 64164 22752 64220
rect 22752 64164 22756 64220
rect 22692 64160 22756 64164
rect 22772 64220 22836 64224
rect 22772 64164 22776 64220
rect 22776 64164 22832 64220
rect 22832 64164 22836 64220
rect 22772 64160 22836 64164
rect 22852 64220 22916 64224
rect 22852 64164 22856 64220
rect 22856 64164 22912 64220
rect 22912 64164 22916 64220
rect 22852 64160 22916 64164
rect 27612 64220 27676 64224
rect 27612 64164 27616 64220
rect 27616 64164 27672 64220
rect 27672 64164 27676 64220
rect 27612 64160 27676 64164
rect 27692 64220 27756 64224
rect 27692 64164 27696 64220
rect 27696 64164 27752 64220
rect 27752 64164 27756 64220
rect 27692 64160 27756 64164
rect 27772 64220 27836 64224
rect 27772 64164 27776 64220
rect 27776 64164 27832 64220
rect 27832 64164 27836 64220
rect 27772 64160 27836 64164
rect 27852 64220 27916 64224
rect 27852 64164 27856 64220
rect 27856 64164 27912 64220
rect 27912 64164 27916 64220
rect 27852 64160 27916 64164
rect 32612 64220 32676 64224
rect 32612 64164 32616 64220
rect 32616 64164 32672 64220
rect 32672 64164 32676 64220
rect 32612 64160 32676 64164
rect 32692 64220 32756 64224
rect 32692 64164 32696 64220
rect 32696 64164 32752 64220
rect 32752 64164 32756 64220
rect 32692 64160 32756 64164
rect 32772 64220 32836 64224
rect 32772 64164 32776 64220
rect 32776 64164 32832 64220
rect 32832 64164 32836 64220
rect 32772 64160 32836 64164
rect 32852 64220 32916 64224
rect 32852 64164 32856 64220
rect 32856 64164 32912 64220
rect 32912 64164 32916 64220
rect 32852 64160 32916 64164
rect 37612 64220 37676 64224
rect 37612 64164 37616 64220
rect 37616 64164 37672 64220
rect 37672 64164 37676 64220
rect 37612 64160 37676 64164
rect 37692 64220 37756 64224
rect 37692 64164 37696 64220
rect 37696 64164 37752 64220
rect 37752 64164 37756 64220
rect 37692 64160 37756 64164
rect 37772 64220 37836 64224
rect 37772 64164 37776 64220
rect 37776 64164 37832 64220
rect 37832 64164 37836 64220
rect 37772 64160 37836 64164
rect 37852 64220 37916 64224
rect 37852 64164 37856 64220
rect 37856 64164 37912 64220
rect 37912 64164 37916 64220
rect 37852 64160 37916 64164
rect 1952 63676 2016 63680
rect 1952 63620 1956 63676
rect 1956 63620 2012 63676
rect 2012 63620 2016 63676
rect 1952 63616 2016 63620
rect 2032 63676 2096 63680
rect 2032 63620 2036 63676
rect 2036 63620 2092 63676
rect 2092 63620 2096 63676
rect 2032 63616 2096 63620
rect 2112 63676 2176 63680
rect 2112 63620 2116 63676
rect 2116 63620 2172 63676
rect 2172 63620 2176 63676
rect 2112 63616 2176 63620
rect 2192 63676 2256 63680
rect 2192 63620 2196 63676
rect 2196 63620 2252 63676
rect 2252 63620 2256 63676
rect 2192 63616 2256 63620
rect 6952 63676 7016 63680
rect 6952 63620 6956 63676
rect 6956 63620 7012 63676
rect 7012 63620 7016 63676
rect 6952 63616 7016 63620
rect 7032 63676 7096 63680
rect 7032 63620 7036 63676
rect 7036 63620 7092 63676
rect 7092 63620 7096 63676
rect 7032 63616 7096 63620
rect 7112 63676 7176 63680
rect 7112 63620 7116 63676
rect 7116 63620 7172 63676
rect 7172 63620 7176 63676
rect 7112 63616 7176 63620
rect 7192 63676 7256 63680
rect 7192 63620 7196 63676
rect 7196 63620 7252 63676
rect 7252 63620 7256 63676
rect 7192 63616 7256 63620
rect 11952 63676 12016 63680
rect 11952 63620 11956 63676
rect 11956 63620 12012 63676
rect 12012 63620 12016 63676
rect 11952 63616 12016 63620
rect 12032 63676 12096 63680
rect 12032 63620 12036 63676
rect 12036 63620 12092 63676
rect 12092 63620 12096 63676
rect 12032 63616 12096 63620
rect 12112 63676 12176 63680
rect 12112 63620 12116 63676
rect 12116 63620 12172 63676
rect 12172 63620 12176 63676
rect 12112 63616 12176 63620
rect 12192 63676 12256 63680
rect 12192 63620 12196 63676
rect 12196 63620 12252 63676
rect 12252 63620 12256 63676
rect 12192 63616 12256 63620
rect 16952 63676 17016 63680
rect 16952 63620 16956 63676
rect 16956 63620 17012 63676
rect 17012 63620 17016 63676
rect 16952 63616 17016 63620
rect 17032 63676 17096 63680
rect 17032 63620 17036 63676
rect 17036 63620 17092 63676
rect 17092 63620 17096 63676
rect 17032 63616 17096 63620
rect 17112 63676 17176 63680
rect 17112 63620 17116 63676
rect 17116 63620 17172 63676
rect 17172 63620 17176 63676
rect 17112 63616 17176 63620
rect 17192 63676 17256 63680
rect 17192 63620 17196 63676
rect 17196 63620 17252 63676
rect 17252 63620 17256 63676
rect 17192 63616 17256 63620
rect 21952 63676 22016 63680
rect 21952 63620 21956 63676
rect 21956 63620 22012 63676
rect 22012 63620 22016 63676
rect 21952 63616 22016 63620
rect 22032 63676 22096 63680
rect 22032 63620 22036 63676
rect 22036 63620 22092 63676
rect 22092 63620 22096 63676
rect 22032 63616 22096 63620
rect 22112 63676 22176 63680
rect 22112 63620 22116 63676
rect 22116 63620 22172 63676
rect 22172 63620 22176 63676
rect 22112 63616 22176 63620
rect 22192 63676 22256 63680
rect 22192 63620 22196 63676
rect 22196 63620 22252 63676
rect 22252 63620 22256 63676
rect 22192 63616 22256 63620
rect 26952 63676 27016 63680
rect 26952 63620 26956 63676
rect 26956 63620 27012 63676
rect 27012 63620 27016 63676
rect 26952 63616 27016 63620
rect 27032 63676 27096 63680
rect 27032 63620 27036 63676
rect 27036 63620 27092 63676
rect 27092 63620 27096 63676
rect 27032 63616 27096 63620
rect 27112 63676 27176 63680
rect 27112 63620 27116 63676
rect 27116 63620 27172 63676
rect 27172 63620 27176 63676
rect 27112 63616 27176 63620
rect 27192 63676 27256 63680
rect 27192 63620 27196 63676
rect 27196 63620 27252 63676
rect 27252 63620 27256 63676
rect 27192 63616 27256 63620
rect 31952 63676 32016 63680
rect 31952 63620 31956 63676
rect 31956 63620 32012 63676
rect 32012 63620 32016 63676
rect 31952 63616 32016 63620
rect 32032 63676 32096 63680
rect 32032 63620 32036 63676
rect 32036 63620 32092 63676
rect 32092 63620 32096 63676
rect 32032 63616 32096 63620
rect 32112 63676 32176 63680
rect 32112 63620 32116 63676
rect 32116 63620 32172 63676
rect 32172 63620 32176 63676
rect 32112 63616 32176 63620
rect 32192 63676 32256 63680
rect 32192 63620 32196 63676
rect 32196 63620 32252 63676
rect 32252 63620 32256 63676
rect 32192 63616 32256 63620
rect 36952 63676 37016 63680
rect 36952 63620 36956 63676
rect 36956 63620 37012 63676
rect 37012 63620 37016 63676
rect 36952 63616 37016 63620
rect 37032 63676 37096 63680
rect 37032 63620 37036 63676
rect 37036 63620 37092 63676
rect 37092 63620 37096 63676
rect 37032 63616 37096 63620
rect 37112 63676 37176 63680
rect 37112 63620 37116 63676
rect 37116 63620 37172 63676
rect 37172 63620 37176 63676
rect 37112 63616 37176 63620
rect 37192 63676 37256 63680
rect 37192 63620 37196 63676
rect 37196 63620 37252 63676
rect 37252 63620 37256 63676
rect 37192 63616 37256 63620
rect 2612 63132 2676 63136
rect 2612 63076 2616 63132
rect 2616 63076 2672 63132
rect 2672 63076 2676 63132
rect 2612 63072 2676 63076
rect 2692 63132 2756 63136
rect 2692 63076 2696 63132
rect 2696 63076 2752 63132
rect 2752 63076 2756 63132
rect 2692 63072 2756 63076
rect 2772 63132 2836 63136
rect 2772 63076 2776 63132
rect 2776 63076 2832 63132
rect 2832 63076 2836 63132
rect 2772 63072 2836 63076
rect 2852 63132 2916 63136
rect 2852 63076 2856 63132
rect 2856 63076 2912 63132
rect 2912 63076 2916 63132
rect 2852 63072 2916 63076
rect 7612 63132 7676 63136
rect 7612 63076 7616 63132
rect 7616 63076 7672 63132
rect 7672 63076 7676 63132
rect 7612 63072 7676 63076
rect 7692 63132 7756 63136
rect 7692 63076 7696 63132
rect 7696 63076 7752 63132
rect 7752 63076 7756 63132
rect 7692 63072 7756 63076
rect 7772 63132 7836 63136
rect 7772 63076 7776 63132
rect 7776 63076 7832 63132
rect 7832 63076 7836 63132
rect 7772 63072 7836 63076
rect 7852 63132 7916 63136
rect 7852 63076 7856 63132
rect 7856 63076 7912 63132
rect 7912 63076 7916 63132
rect 7852 63072 7916 63076
rect 12612 63132 12676 63136
rect 12612 63076 12616 63132
rect 12616 63076 12672 63132
rect 12672 63076 12676 63132
rect 12612 63072 12676 63076
rect 12692 63132 12756 63136
rect 12692 63076 12696 63132
rect 12696 63076 12752 63132
rect 12752 63076 12756 63132
rect 12692 63072 12756 63076
rect 12772 63132 12836 63136
rect 12772 63076 12776 63132
rect 12776 63076 12832 63132
rect 12832 63076 12836 63132
rect 12772 63072 12836 63076
rect 12852 63132 12916 63136
rect 12852 63076 12856 63132
rect 12856 63076 12912 63132
rect 12912 63076 12916 63132
rect 12852 63072 12916 63076
rect 17612 63132 17676 63136
rect 17612 63076 17616 63132
rect 17616 63076 17672 63132
rect 17672 63076 17676 63132
rect 17612 63072 17676 63076
rect 17692 63132 17756 63136
rect 17692 63076 17696 63132
rect 17696 63076 17752 63132
rect 17752 63076 17756 63132
rect 17692 63072 17756 63076
rect 17772 63132 17836 63136
rect 17772 63076 17776 63132
rect 17776 63076 17832 63132
rect 17832 63076 17836 63132
rect 17772 63072 17836 63076
rect 17852 63132 17916 63136
rect 17852 63076 17856 63132
rect 17856 63076 17912 63132
rect 17912 63076 17916 63132
rect 17852 63072 17916 63076
rect 22612 63132 22676 63136
rect 22612 63076 22616 63132
rect 22616 63076 22672 63132
rect 22672 63076 22676 63132
rect 22612 63072 22676 63076
rect 22692 63132 22756 63136
rect 22692 63076 22696 63132
rect 22696 63076 22752 63132
rect 22752 63076 22756 63132
rect 22692 63072 22756 63076
rect 22772 63132 22836 63136
rect 22772 63076 22776 63132
rect 22776 63076 22832 63132
rect 22832 63076 22836 63132
rect 22772 63072 22836 63076
rect 22852 63132 22916 63136
rect 22852 63076 22856 63132
rect 22856 63076 22912 63132
rect 22912 63076 22916 63132
rect 22852 63072 22916 63076
rect 27612 63132 27676 63136
rect 27612 63076 27616 63132
rect 27616 63076 27672 63132
rect 27672 63076 27676 63132
rect 27612 63072 27676 63076
rect 27692 63132 27756 63136
rect 27692 63076 27696 63132
rect 27696 63076 27752 63132
rect 27752 63076 27756 63132
rect 27692 63072 27756 63076
rect 27772 63132 27836 63136
rect 27772 63076 27776 63132
rect 27776 63076 27832 63132
rect 27832 63076 27836 63132
rect 27772 63072 27836 63076
rect 27852 63132 27916 63136
rect 27852 63076 27856 63132
rect 27856 63076 27912 63132
rect 27912 63076 27916 63132
rect 27852 63072 27916 63076
rect 32612 63132 32676 63136
rect 32612 63076 32616 63132
rect 32616 63076 32672 63132
rect 32672 63076 32676 63132
rect 32612 63072 32676 63076
rect 32692 63132 32756 63136
rect 32692 63076 32696 63132
rect 32696 63076 32752 63132
rect 32752 63076 32756 63132
rect 32692 63072 32756 63076
rect 32772 63132 32836 63136
rect 32772 63076 32776 63132
rect 32776 63076 32832 63132
rect 32832 63076 32836 63132
rect 32772 63072 32836 63076
rect 32852 63132 32916 63136
rect 32852 63076 32856 63132
rect 32856 63076 32912 63132
rect 32912 63076 32916 63132
rect 32852 63072 32916 63076
rect 37612 63132 37676 63136
rect 37612 63076 37616 63132
rect 37616 63076 37672 63132
rect 37672 63076 37676 63132
rect 37612 63072 37676 63076
rect 37692 63132 37756 63136
rect 37692 63076 37696 63132
rect 37696 63076 37752 63132
rect 37752 63076 37756 63132
rect 37692 63072 37756 63076
rect 37772 63132 37836 63136
rect 37772 63076 37776 63132
rect 37776 63076 37832 63132
rect 37832 63076 37836 63132
rect 37772 63072 37836 63076
rect 37852 63132 37916 63136
rect 37852 63076 37856 63132
rect 37856 63076 37912 63132
rect 37912 63076 37916 63132
rect 37852 63072 37916 63076
rect 1952 62588 2016 62592
rect 1952 62532 1956 62588
rect 1956 62532 2012 62588
rect 2012 62532 2016 62588
rect 1952 62528 2016 62532
rect 2032 62588 2096 62592
rect 2032 62532 2036 62588
rect 2036 62532 2092 62588
rect 2092 62532 2096 62588
rect 2032 62528 2096 62532
rect 2112 62588 2176 62592
rect 2112 62532 2116 62588
rect 2116 62532 2172 62588
rect 2172 62532 2176 62588
rect 2112 62528 2176 62532
rect 2192 62588 2256 62592
rect 2192 62532 2196 62588
rect 2196 62532 2252 62588
rect 2252 62532 2256 62588
rect 2192 62528 2256 62532
rect 6952 62588 7016 62592
rect 6952 62532 6956 62588
rect 6956 62532 7012 62588
rect 7012 62532 7016 62588
rect 6952 62528 7016 62532
rect 7032 62588 7096 62592
rect 7032 62532 7036 62588
rect 7036 62532 7092 62588
rect 7092 62532 7096 62588
rect 7032 62528 7096 62532
rect 7112 62588 7176 62592
rect 7112 62532 7116 62588
rect 7116 62532 7172 62588
rect 7172 62532 7176 62588
rect 7112 62528 7176 62532
rect 7192 62588 7256 62592
rect 7192 62532 7196 62588
rect 7196 62532 7252 62588
rect 7252 62532 7256 62588
rect 7192 62528 7256 62532
rect 11952 62588 12016 62592
rect 11952 62532 11956 62588
rect 11956 62532 12012 62588
rect 12012 62532 12016 62588
rect 11952 62528 12016 62532
rect 12032 62588 12096 62592
rect 12032 62532 12036 62588
rect 12036 62532 12092 62588
rect 12092 62532 12096 62588
rect 12032 62528 12096 62532
rect 12112 62588 12176 62592
rect 12112 62532 12116 62588
rect 12116 62532 12172 62588
rect 12172 62532 12176 62588
rect 12112 62528 12176 62532
rect 12192 62588 12256 62592
rect 12192 62532 12196 62588
rect 12196 62532 12252 62588
rect 12252 62532 12256 62588
rect 12192 62528 12256 62532
rect 16952 62588 17016 62592
rect 16952 62532 16956 62588
rect 16956 62532 17012 62588
rect 17012 62532 17016 62588
rect 16952 62528 17016 62532
rect 17032 62588 17096 62592
rect 17032 62532 17036 62588
rect 17036 62532 17092 62588
rect 17092 62532 17096 62588
rect 17032 62528 17096 62532
rect 17112 62588 17176 62592
rect 17112 62532 17116 62588
rect 17116 62532 17172 62588
rect 17172 62532 17176 62588
rect 17112 62528 17176 62532
rect 17192 62588 17256 62592
rect 17192 62532 17196 62588
rect 17196 62532 17252 62588
rect 17252 62532 17256 62588
rect 17192 62528 17256 62532
rect 21952 62588 22016 62592
rect 21952 62532 21956 62588
rect 21956 62532 22012 62588
rect 22012 62532 22016 62588
rect 21952 62528 22016 62532
rect 22032 62588 22096 62592
rect 22032 62532 22036 62588
rect 22036 62532 22092 62588
rect 22092 62532 22096 62588
rect 22032 62528 22096 62532
rect 22112 62588 22176 62592
rect 22112 62532 22116 62588
rect 22116 62532 22172 62588
rect 22172 62532 22176 62588
rect 22112 62528 22176 62532
rect 22192 62588 22256 62592
rect 22192 62532 22196 62588
rect 22196 62532 22252 62588
rect 22252 62532 22256 62588
rect 22192 62528 22256 62532
rect 26952 62588 27016 62592
rect 26952 62532 26956 62588
rect 26956 62532 27012 62588
rect 27012 62532 27016 62588
rect 26952 62528 27016 62532
rect 27032 62588 27096 62592
rect 27032 62532 27036 62588
rect 27036 62532 27092 62588
rect 27092 62532 27096 62588
rect 27032 62528 27096 62532
rect 27112 62588 27176 62592
rect 27112 62532 27116 62588
rect 27116 62532 27172 62588
rect 27172 62532 27176 62588
rect 27112 62528 27176 62532
rect 27192 62588 27256 62592
rect 27192 62532 27196 62588
rect 27196 62532 27252 62588
rect 27252 62532 27256 62588
rect 27192 62528 27256 62532
rect 31952 62588 32016 62592
rect 31952 62532 31956 62588
rect 31956 62532 32012 62588
rect 32012 62532 32016 62588
rect 31952 62528 32016 62532
rect 32032 62588 32096 62592
rect 32032 62532 32036 62588
rect 32036 62532 32092 62588
rect 32092 62532 32096 62588
rect 32032 62528 32096 62532
rect 32112 62588 32176 62592
rect 32112 62532 32116 62588
rect 32116 62532 32172 62588
rect 32172 62532 32176 62588
rect 32112 62528 32176 62532
rect 32192 62588 32256 62592
rect 32192 62532 32196 62588
rect 32196 62532 32252 62588
rect 32252 62532 32256 62588
rect 32192 62528 32256 62532
rect 36952 62588 37016 62592
rect 36952 62532 36956 62588
rect 36956 62532 37012 62588
rect 37012 62532 37016 62588
rect 36952 62528 37016 62532
rect 37032 62588 37096 62592
rect 37032 62532 37036 62588
rect 37036 62532 37092 62588
rect 37092 62532 37096 62588
rect 37032 62528 37096 62532
rect 37112 62588 37176 62592
rect 37112 62532 37116 62588
rect 37116 62532 37172 62588
rect 37172 62532 37176 62588
rect 37112 62528 37176 62532
rect 37192 62588 37256 62592
rect 37192 62532 37196 62588
rect 37196 62532 37252 62588
rect 37252 62532 37256 62588
rect 37192 62528 37256 62532
rect 2612 62044 2676 62048
rect 2612 61988 2616 62044
rect 2616 61988 2672 62044
rect 2672 61988 2676 62044
rect 2612 61984 2676 61988
rect 2692 62044 2756 62048
rect 2692 61988 2696 62044
rect 2696 61988 2752 62044
rect 2752 61988 2756 62044
rect 2692 61984 2756 61988
rect 2772 62044 2836 62048
rect 2772 61988 2776 62044
rect 2776 61988 2832 62044
rect 2832 61988 2836 62044
rect 2772 61984 2836 61988
rect 2852 62044 2916 62048
rect 2852 61988 2856 62044
rect 2856 61988 2912 62044
rect 2912 61988 2916 62044
rect 2852 61984 2916 61988
rect 7612 62044 7676 62048
rect 7612 61988 7616 62044
rect 7616 61988 7672 62044
rect 7672 61988 7676 62044
rect 7612 61984 7676 61988
rect 7692 62044 7756 62048
rect 7692 61988 7696 62044
rect 7696 61988 7752 62044
rect 7752 61988 7756 62044
rect 7692 61984 7756 61988
rect 7772 62044 7836 62048
rect 7772 61988 7776 62044
rect 7776 61988 7832 62044
rect 7832 61988 7836 62044
rect 7772 61984 7836 61988
rect 7852 62044 7916 62048
rect 7852 61988 7856 62044
rect 7856 61988 7912 62044
rect 7912 61988 7916 62044
rect 7852 61984 7916 61988
rect 12612 62044 12676 62048
rect 12612 61988 12616 62044
rect 12616 61988 12672 62044
rect 12672 61988 12676 62044
rect 12612 61984 12676 61988
rect 12692 62044 12756 62048
rect 12692 61988 12696 62044
rect 12696 61988 12752 62044
rect 12752 61988 12756 62044
rect 12692 61984 12756 61988
rect 12772 62044 12836 62048
rect 12772 61988 12776 62044
rect 12776 61988 12832 62044
rect 12832 61988 12836 62044
rect 12772 61984 12836 61988
rect 12852 62044 12916 62048
rect 12852 61988 12856 62044
rect 12856 61988 12912 62044
rect 12912 61988 12916 62044
rect 12852 61984 12916 61988
rect 17612 62044 17676 62048
rect 17612 61988 17616 62044
rect 17616 61988 17672 62044
rect 17672 61988 17676 62044
rect 17612 61984 17676 61988
rect 17692 62044 17756 62048
rect 17692 61988 17696 62044
rect 17696 61988 17752 62044
rect 17752 61988 17756 62044
rect 17692 61984 17756 61988
rect 17772 62044 17836 62048
rect 17772 61988 17776 62044
rect 17776 61988 17832 62044
rect 17832 61988 17836 62044
rect 17772 61984 17836 61988
rect 17852 62044 17916 62048
rect 17852 61988 17856 62044
rect 17856 61988 17912 62044
rect 17912 61988 17916 62044
rect 17852 61984 17916 61988
rect 22612 62044 22676 62048
rect 22612 61988 22616 62044
rect 22616 61988 22672 62044
rect 22672 61988 22676 62044
rect 22612 61984 22676 61988
rect 22692 62044 22756 62048
rect 22692 61988 22696 62044
rect 22696 61988 22752 62044
rect 22752 61988 22756 62044
rect 22692 61984 22756 61988
rect 22772 62044 22836 62048
rect 22772 61988 22776 62044
rect 22776 61988 22832 62044
rect 22832 61988 22836 62044
rect 22772 61984 22836 61988
rect 22852 62044 22916 62048
rect 22852 61988 22856 62044
rect 22856 61988 22912 62044
rect 22912 61988 22916 62044
rect 22852 61984 22916 61988
rect 27612 62044 27676 62048
rect 27612 61988 27616 62044
rect 27616 61988 27672 62044
rect 27672 61988 27676 62044
rect 27612 61984 27676 61988
rect 27692 62044 27756 62048
rect 27692 61988 27696 62044
rect 27696 61988 27752 62044
rect 27752 61988 27756 62044
rect 27692 61984 27756 61988
rect 27772 62044 27836 62048
rect 27772 61988 27776 62044
rect 27776 61988 27832 62044
rect 27832 61988 27836 62044
rect 27772 61984 27836 61988
rect 27852 62044 27916 62048
rect 27852 61988 27856 62044
rect 27856 61988 27912 62044
rect 27912 61988 27916 62044
rect 27852 61984 27916 61988
rect 32612 62044 32676 62048
rect 32612 61988 32616 62044
rect 32616 61988 32672 62044
rect 32672 61988 32676 62044
rect 32612 61984 32676 61988
rect 32692 62044 32756 62048
rect 32692 61988 32696 62044
rect 32696 61988 32752 62044
rect 32752 61988 32756 62044
rect 32692 61984 32756 61988
rect 32772 62044 32836 62048
rect 32772 61988 32776 62044
rect 32776 61988 32832 62044
rect 32832 61988 32836 62044
rect 32772 61984 32836 61988
rect 32852 62044 32916 62048
rect 32852 61988 32856 62044
rect 32856 61988 32912 62044
rect 32912 61988 32916 62044
rect 32852 61984 32916 61988
rect 37612 62044 37676 62048
rect 37612 61988 37616 62044
rect 37616 61988 37672 62044
rect 37672 61988 37676 62044
rect 37612 61984 37676 61988
rect 37692 62044 37756 62048
rect 37692 61988 37696 62044
rect 37696 61988 37752 62044
rect 37752 61988 37756 62044
rect 37692 61984 37756 61988
rect 37772 62044 37836 62048
rect 37772 61988 37776 62044
rect 37776 61988 37832 62044
rect 37832 61988 37836 62044
rect 37772 61984 37836 61988
rect 37852 62044 37916 62048
rect 37852 61988 37856 62044
rect 37856 61988 37912 62044
rect 37912 61988 37916 62044
rect 37852 61984 37916 61988
rect 1952 61500 2016 61504
rect 1952 61444 1956 61500
rect 1956 61444 2012 61500
rect 2012 61444 2016 61500
rect 1952 61440 2016 61444
rect 2032 61500 2096 61504
rect 2032 61444 2036 61500
rect 2036 61444 2092 61500
rect 2092 61444 2096 61500
rect 2032 61440 2096 61444
rect 2112 61500 2176 61504
rect 2112 61444 2116 61500
rect 2116 61444 2172 61500
rect 2172 61444 2176 61500
rect 2112 61440 2176 61444
rect 2192 61500 2256 61504
rect 2192 61444 2196 61500
rect 2196 61444 2252 61500
rect 2252 61444 2256 61500
rect 2192 61440 2256 61444
rect 6952 61500 7016 61504
rect 6952 61444 6956 61500
rect 6956 61444 7012 61500
rect 7012 61444 7016 61500
rect 6952 61440 7016 61444
rect 7032 61500 7096 61504
rect 7032 61444 7036 61500
rect 7036 61444 7092 61500
rect 7092 61444 7096 61500
rect 7032 61440 7096 61444
rect 7112 61500 7176 61504
rect 7112 61444 7116 61500
rect 7116 61444 7172 61500
rect 7172 61444 7176 61500
rect 7112 61440 7176 61444
rect 7192 61500 7256 61504
rect 7192 61444 7196 61500
rect 7196 61444 7252 61500
rect 7252 61444 7256 61500
rect 7192 61440 7256 61444
rect 11952 61500 12016 61504
rect 11952 61444 11956 61500
rect 11956 61444 12012 61500
rect 12012 61444 12016 61500
rect 11952 61440 12016 61444
rect 12032 61500 12096 61504
rect 12032 61444 12036 61500
rect 12036 61444 12092 61500
rect 12092 61444 12096 61500
rect 12032 61440 12096 61444
rect 12112 61500 12176 61504
rect 12112 61444 12116 61500
rect 12116 61444 12172 61500
rect 12172 61444 12176 61500
rect 12112 61440 12176 61444
rect 12192 61500 12256 61504
rect 12192 61444 12196 61500
rect 12196 61444 12252 61500
rect 12252 61444 12256 61500
rect 12192 61440 12256 61444
rect 16952 61500 17016 61504
rect 16952 61444 16956 61500
rect 16956 61444 17012 61500
rect 17012 61444 17016 61500
rect 16952 61440 17016 61444
rect 17032 61500 17096 61504
rect 17032 61444 17036 61500
rect 17036 61444 17092 61500
rect 17092 61444 17096 61500
rect 17032 61440 17096 61444
rect 17112 61500 17176 61504
rect 17112 61444 17116 61500
rect 17116 61444 17172 61500
rect 17172 61444 17176 61500
rect 17112 61440 17176 61444
rect 17192 61500 17256 61504
rect 17192 61444 17196 61500
rect 17196 61444 17252 61500
rect 17252 61444 17256 61500
rect 17192 61440 17256 61444
rect 21952 61500 22016 61504
rect 21952 61444 21956 61500
rect 21956 61444 22012 61500
rect 22012 61444 22016 61500
rect 21952 61440 22016 61444
rect 22032 61500 22096 61504
rect 22032 61444 22036 61500
rect 22036 61444 22092 61500
rect 22092 61444 22096 61500
rect 22032 61440 22096 61444
rect 22112 61500 22176 61504
rect 22112 61444 22116 61500
rect 22116 61444 22172 61500
rect 22172 61444 22176 61500
rect 22112 61440 22176 61444
rect 22192 61500 22256 61504
rect 22192 61444 22196 61500
rect 22196 61444 22252 61500
rect 22252 61444 22256 61500
rect 22192 61440 22256 61444
rect 26952 61500 27016 61504
rect 26952 61444 26956 61500
rect 26956 61444 27012 61500
rect 27012 61444 27016 61500
rect 26952 61440 27016 61444
rect 27032 61500 27096 61504
rect 27032 61444 27036 61500
rect 27036 61444 27092 61500
rect 27092 61444 27096 61500
rect 27032 61440 27096 61444
rect 27112 61500 27176 61504
rect 27112 61444 27116 61500
rect 27116 61444 27172 61500
rect 27172 61444 27176 61500
rect 27112 61440 27176 61444
rect 27192 61500 27256 61504
rect 27192 61444 27196 61500
rect 27196 61444 27252 61500
rect 27252 61444 27256 61500
rect 27192 61440 27256 61444
rect 31952 61500 32016 61504
rect 31952 61444 31956 61500
rect 31956 61444 32012 61500
rect 32012 61444 32016 61500
rect 31952 61440 32016 61444
rect 32032 61500 32096 61504
rect 32032 61444 32036 61500
rect 32036 61444 32092 61500
rect 32092 61444 32096 61500
rect 32032 61440 32096 61444
rect 32112 61500 32176 61504
rect 32112 61444 32116 61500
rect 32116 61444 32172 61500
rect 32172 61444 32176 61500
rect 32112 61440 32176 61444
rect 32192 61500 32256 61504
rect 32192 61444 32196 61500
rect 32196 61444 32252 61500
rect 32252 61444 32256 61500
rect 32192 61440 32256 61444
rect 36952 61500 37016 61504
rect 36952 61444 36956 61500
rect 36956 61444 37012 61500
rect 37012 61444 37016 61500
rect 36952 61440 37016 61444
rect 37032 61500 37096 61504
rect 37032 61444 37036 61500
rect 37036 61444 37092 61500
rect 37092 61444 37096 61500
rect 37032 61440 37096 61444
rect 37112 61500 37176 61504
rect 37112 61444 37116 61500
rect 37116 61444 37172 61500
rect 37172 61444 37176 61500
rect 37112 61440 37176 61444
rect 37192 61500 37256 61504
rect 37192 61444 37196 61500
rect 37196 61444 37252 61500
rect 37252 61444 37256 61500
rect 37192 61440 37256 61444
rect 2612 60956 2676 60960
rect 2612 60900 2616 60956
rect 2616 60900 2672 60956
rect 2672 60900 2676 60956
rect 2612 60896 2676 60900
rect 2692 60956 2756 60960
rect 2692 60900 2696 60956
rect 2696 60900 2752 60956
rect 2752 60900 2756 60956
rect 2692 60896 2756 60900
rect 2772 60956 2836 60960
rect 2772 60900 2776 60956
rect 2776 60900 2832 60956
rect 2832 60900 2836 60956
rect 2772 60896 2836 60900
rect 2852 60956 2916 60960
rect 2852 60900 2856 60956
rect 2856 60900 2912 60956
rect 2912 60900 2916 60956
rect 2852 60896 2916 60900
rect 7612 60956 7676 60960
rect 7612 60900 7616 60956
rect 7616 60900 7672 60956
rect 7672 60900 7676 60956
rect 7612 60896 7676 60900
rect 7692 60956 7756 60960
rect 7692 60900 7696 60956
rect 7696 60900 7752 60956
rect 7752 60900 7756 60956
rect 7692 60896 7756 60900
rect 7772 60956 7836 60960
rect 7772 60900 7776 60956
rect 7776 60900 7832 60956
rect 7832 60900 7836 60956
rect 7772 60896 7836 60900
rect 7852 60956 7916 60960
rect 7852 60900 7856 60956
rect 7856 60900 7912 60956
rect 7912 60900 7916 60956
rect 7852 60896 7916 60900
rect 12612 60956 12676 60960
rect 12612 60900 12616 60956
rect 12616 60900 12672 60956
rect 12672 60900 12676 60956
rect 12612 60896 12676 60900
rect 12692 60956 12756 60960
rect 12692 60900 12696 60956
rect 12696 60900 12752 60956
rect 12752 60900 12756 60956
rect 12692 60896 12756 60900
rect 12772 60956 12836 60960
rect 12772 60900 12776 60956
rect 12776 60900 12832 60956
rect 12832 60900 12836 60956
rect 12772 60896 12836 60900
rect 12852 60956 12916 60960
rect 12852 60900 12856 60956
rect 12856 60900 12912 60956
rect 12912 60900 12916 60956
rect 12852 60896 12916 60900
rect 17612 60956 17676 60960
rect 17612 60900 17616 60956
rect 17616 60900 17672 60956
rect 17672 60900 17676 60956
rect 17612 60896 17676 60900
rect 17692 60956 17756 60960
rect 17692 60900 17696 60956
rect 17696 60900 17752 60956
rect 17752 60900 17756 60956
rect 17692 60896 17756 60900
rect 17772 60956 17836 60960
rect 17772 60900 17776 60956
rect 17776 60900 17832 60956
rect 17832 60900 17836 60956
rect 17772 60896 17836 60900
rect 17852 60956 17916 60960
rect 17852 60900 17856 60956
rect 17856 60900 17912 60956
rect 17912 60900 17916 60956
rect 17852 60896 17916 60900
rect 22612 60956 22676 60960
rect 22612 60900 22616 60956
rect 22616 60900 22672 60956
rect 22672 60900 22676 60956
rect 22612 60896 22676 60900
rect 22692 60956 22756 60960
rect 22692 60900 22696 60956
rect 22696 60900 22752 60956
rect 22752 60900 22756 60956
rect 22692 60896 22756 60900
rect 22772 60956 22836 60960
rect 22772 60900 22776 60956
rect 22776 60900 22832 60956
rect 22832 60900 22836 60956
rect 22772 60896 22836 60900
rect 22852 60956 22916 60960
rect 22852 60900 22856 60956
rect 22856 60900 22912 60956
rect 22912 60900 22916 60956
rect 22852 60896 22916 60900
rect 27612 60956 27676 60960
rect 27612 60900 27616 60956
rect 27616 60900 27672 60956
rect 27672 60900 27676 60956
rect 27612 60896 27676 60900
rect 27692 60956 27756 60960
rect 27692 60900 27696 60956
rect 27696 60900 27752 60956
rect 27752 60900 27756 60956
rect 27692 60896 27756 60900
rect 27772 60956 27836 60960
rect 27772 60900 27776 60956
rect 27776 60900 27832 60956
rect 27832 60900 27836 60956
rect 27772 60896 27836 60900
rect 27852 60956 27916 60960
rect 27852 60900 27856 60956
rect 27856 60900 27912 60956
rect 27912 60900 27916 60956
rect 27852 60896 27916 60900
rect 32612 60956 32676 60960
rect 32612 60900 32616 60956
rect 32616 60900 32672 60956
rect 32672 60900 32676 60956
rect 32612 60896 32676 60900
rect 32692 60956 32756 60960
rect 32692 60900 32696 60956
rect 32696 60900 32752 60956
rect 32752 60900 32756 60956
rect 32692 60896 32756 60900
rect 32772 60956 32836 60960
rect 32772 60900 32776 60956
rect 32776 60900 32832 60956
rect 32832 60900 32836 60956
rect 32772 60896 32836 60900
rect 32852 60956 32916 60960
rect 32852 60900 32856 60956
rect 32856 60900 32912 60956
rect 32912 60900 32916 60956
rect 32852 60896 32916 60900
rect 37612 60956 37676 60960
rect 37612 60900 37616 60956
rect 37616 60900 37672 60956
rect 37672 60900 37676 60956
rect 37612 60896 37676 60900
rect 37692 60956 37756 60960
rect 37692 60900 37696 60956
rect 37696 60900 37752 60956
rect 37752 60900 37756 60956
rect 37692 60896 37756 60900
rect 37772 60956 37836 60960
rect 37772 60900 37776 60956
rect 37776 60900 37832 60956
rect 37832 60900 37836 60956
rect 37772 60896 37836 60900
rect 37852 60956 37916 60960
rect 37852 60900 37856 60956
rect 37856 60900 37912 60956
rect 37912 60900 37916 60956
rect 37852 60896 37916 60900
rect 1952 60412 2016 60416
rect 1952 60356 1956 60412
rect 1956 60356 2012 60412
rect 2012 60356 2016 60412
rect 1952 60352 2016 60356
rect 2032 60412 2096 60416
rect 2032 60356 2036 60412
rect 2036 60356 2092 60412
rect 2092 60356 2096 60412
rect 2032 60352 2096 60356
rect 2112 60412 2176 60416
rect 2112 60356 2116 60412
rect 2116 60356 2172 60412
rect 2172 60356 2176 60412
rect 2112 60352 2176 60356
rect 2192 60412 2256 60416
rect 2192 60356 2196 60412
rect 2196 60356 2252 60412
rect 2252 60356 2256 60412
rect 2192 60352 2256 60356
rect 6952 60412 7016 60416
rect 6952 60356 6956 60412
rect 6956 60356 7012 60412
rect 7012 60356 7016 60412
rect 6952 60352 7016 60356
rect 7032 60412 7096 60416
rect 7032 60356 7036 60412
rect 7036 60356 7092 60412
rect 7092 60356 7096 60412
rect 7032 60352 7096 60356
rect 7112 60412 7176 60416
rect 7112 60356 7116 60412
rect 7116 60356 7172 60412
rect 7172 60356 7176 60412
rect 7112 60352 7176 60356
rect 7192 60412 7256 60416
rect 7192 60356 7196 60412
rect 7196 60356 7252 60412
rect 7252 60356 7256 60412
rect 7192 60352 7256 60356
rect 11952 60412 12016 60416
rect 11952 60356 11956 60412
rect 11956 60356 12012 60412
rect 12012 60356 12016 60412
rect 11952 60352 12016 60356
rect 12032 60412 12096 60416
rect 12032 60356 12036 60412
rect 12036 60356 12092 60412
rect 12092 60356 12096 60412
rect 12032 60352 12096 60356
rect 12112 60412 12176 60416
rect 12112 60356 12116 60412
rect 12116 60356 12172 60412
rect 12172 60356 12176 60412
rect 12112 60352 12176 60356
rect 12192 60412 12256 60416
rect 12192 60356 12196 60412
rect 12196 60356 12252 60412
rect 12252 60356 12256 60412
rect 12192 60352 12256 60356
rect 16952 60412 17016 60416
rect 16952 60356 16956 60412
rect 16956 60356 17012 60412
rect 17012 60356 17016 60412
rect 16952 60352 17016 60356
rect 17032 60412 17096 60416
rect 17032 60356 17036 60412
rect 17036 60356 17092 60412
rect 17092 60356 17096 60412
rect 17032 60352 17096 60356
rect 17112 60412 17176 60416
rect 17112 60356 17116 60412
rect 17116 60356 17172 60412
rect 17172 60356 17176 60412
rect 17112 60352 17176 60356
rect 17192 60412 17256 60416
rect 17192 60356 17196 60412
rect 17196 60356 17252 60412
rect 17252 60356 17256 60412
rect 17192 60352 17256 60356
rect 21952 60412 22016 60416
rect 21952 60356 21956 60412
rect 21956 60356 22012 60412
rect 22012 60356 22016 60412
rect 21952 60352 22016 60356
rect 22032 60412 22096 60416
rect 22032 60356 22036 60412
rect 22036 60356 22092 60412
rect 22092 60356 22096 60412
rect 22032 60352 22096 60356
rect 22112 60412 22176 60416
rect 22112 60356 22116 60412
rect 22116 60356 22172 60412
rect 22172 60356 22176 60412
rect 22112 60352 22176 60356
rect 22192 60412 22256 60416
rect 22192 60356 22196 60412
rect 22196 60356 22252 60412
rect 22252 60356 22256 60412
rect 22192 60352 22256 60356
rect 26952 60412 27016 60416
rect 26952 60356 26956 60412
rect 26956 60356 27012 60412
rect 27012 60356 27016 60412
rect 26952 60352 27016 60356
rect 27032 60412 27096 60416
rect 27032 60356 27036 60412
rect 27036 60356 27092 60412
rect 27092 60356 27096 60412
rect 27032 60352 27096 60356
rect 27112 60412 27176 60416
rect 27112 60356 27116 60412
rect 27116 60356 27172 60412
rect 27172 60356 27176 60412
rect 27112 60352 27176 60356
rect 27192 60412 27256 60416
rect 27192 60356 27196 60412
rect 27196 60356 27252 60412
rect 27252 60356 27256 60412
rect 27192 60352 27256 60356
rect 31952 60412 32016 60416
rect 31952 60356 31956 60412
rect 31956 60356 32012 60412
rect 32012 60356 32016 60412
rect 31952 60352 32016 60356
rect 32032 60412 32096 60416
rect 32032 60356 32036 60412
rect 32036 60356 32092 60412
rect 32092 60356 32096 60412
rect 32032 60352 32096 60356
rect 32112 60412 32176 60416
rect 32112 60356 32116 60412
rect 32116 60356 32172 60412
rect 32172 60356 32176 60412
rect 32112 60352 32176 60356
rect 32192 60412 32256 60416
rect 32192 60356 32196 60412
rect 32196 60356 32252 60412
rect 32252 60356 32256 60412
rect 32192 60352 32256 60356
rect 36952 60412 37016 60416
rect 36952 60356 36956 60412
rect 36956 60356 37012 60412
rect 37012 60356 37016 60412
rect 36952 60352 37016 60356
rect 37032 60412 37096 60416
rect 37032 60356 37036 60412
rect 37036 60356 37092 60412
rect 37092 60356 37096 60412
rect 37032 60352 37096 60356
rect 37112 60412 37176 60416
rect 37112 60356 37116 60412
rect 37116 60356 37172 60412
rect 37172 60356 37176 60412
rect 37112 60352 37176 60356
rect 37192 60412 37256 60416
rect 37192 60356 37196 60412
rect 37196 60356 37252 60412
rect 37252 60356 37256 60412
rect 37192 60352 37256 60356
rect 2612 59868 2676 59872
rect 2612 59812 2616 59868
rect 2616 59812 2672 59868
rect 2672 59812 2676 59868
rect 2612 59808 2676 59812
rect 2692 59868 2756 59872
rect 2692 59812 2696 59868
rect 2696 59812 2752 59868
rect 2752 59812 2756 59868
rect 2692 59808 2756 59812
rect 2772 59868 2836 59872
rect 2772 59812 2776 59868
rect 2776 59812 2832 59868
rect 2832 59812 2836 59868
rect 2772 59808 2836 59812
rect 2852 59868 2916 59872
rect 2852 59812 2856 59868
rect 2856 59812 2912 59868
rect 2912 59812 2916 59868
rect 2852 59808 2916 59812
rect 7612 59868 7676 59872
rect 7612 59812 7616 59868
rect 7616 59812 7672 59868
rect 7672 59812 7676 59868
rect 7612 59808 7676 59812
rect 7692 59868 7756 59872
rect 7692 59812 7696 59868
rect 7696 59812 7752 59868
rect 7752 59812 7756 59868
rect 7692 59808 7756 59812
rect 7772 59868 7836 59872
rect 7772 59812 7776 59868
rect 7776 59812 7832 59868
rect 7832 59812 7836 59868
rect 7772 59808 7836 59812
rect 7852 59868 7916 59872
rect 7852 59812 7856 59868
rect 7856 59812 7912 59868
rect 7912 59812 7916 59868
rect 7852 59808 7916 59812
rect 12612 59868 12676 59872
rect 12612 59812 12616 59868
rect 12616 59812 12672 59868
rect 12672 59812 12676 59868
rect 12612 59808 12676 59812
rect 12692 59868 12756 59872
rect 12692 59812 12696 59868
rect 12696 59812 12752 59868
rect 12752 59812 12756 59868
rect 12692 59808 12756 59812
rect 12772 59868 12836 59872
rect 12772 59812 12776 59868
rect 12776 59812 12832 59868
rect 12832 59812 12836 59868
rect 12772 59808 12836 59812
rect 12852 59868 12916 59872
rect 12852 59812 12856 59868
rect 12856 59812 12912 59868
rect 12912 59812 12916 59868
rect 12852 59808 12916 59812
rect 17612 59868 17676 59872
rect 17612 59812 17616 59868
rect 17616 59812 17672 59868
rect 17672 59812 17676 59868
rect 17612 59808 17676 59812
rect 17692 59868 17756 59872
rect 17692 59812 17696 59868
rect 17696 59812 17752 59868
rect 17752 59812 17756 59868
rect 17692 59808 17756 59812
rect 17772 59868 17836 59872
rect 17772 59812 17776 59868
rect 17776 59812 17832 59868
rect 17832 59812 17836 59868
rect 17772 59808 17836 59812
rect 17852 59868 17916 59872
rect 17852 59812 17856 59868
rect 17856 59812 17912 59868
rect 17912 59812 17916 59868
rect 17852 59808 17916 59812
rect 22612 59868 22676 59872
rect 22612 59812 22616 59868
rect 22616 59812 22672 59868
rect 22672 59812 22676 59868
rect 22612 59808 22676 59812
rect 22692 59868 22756 59872
rect 22692 59812 22696 59868
rect 22696 59812 22752 59868
rect 22752 59812 22756 59868
rect 22692 59808 22756 59812
rect 22772 59868 22836 59872
rect 22772 59812 22776 59868
rect 22776 59812 22832 59868
rect 22832 59812 22836 59868
rect 22772 59808 22836 59812
rect 22852 59868 22916 59872
rect 22852 59812 22856 59868
rect 22856 59812 22912 59868
rect 22912 59812 22916 59868
rect 22852 59808 22916 59812
rect 27612 59868 27676 59872
rect 27612 59812 27616 59868
rect 27616 59812 27672 59868
rect 27672 59812 27676 59868
rect 27612 59808 27676 59812
rect 27692 59868 27756 59872
rect 27692 59812 27696 59868
rect 27696 59812 27752 59868
rect 27752 59812 27756 59868
rect 27692 59808 27756 59812
rect 27772 59868 27836 59872
rect 27772 59812 27776 59868
rect 27776 59812 27832 59868
rect 27832 59812 27836 59868
rect 27772 59808 27836 59812
rect 27852 59868 27916 59872
rect 27852 59812 27856 59868
rect 27856 59812 27912 59868
rect 27912 59812 27916 59868
rect 27852 59808 27916 59812
rect 32612 59868 32676 59872
rect 32612 59812 32616 59868
rect 32616 59812 32672 59868
rect 32672 59812 32676 59868
rect 32612 59808 32676 59812
rect 32692 59868 32756 59872
rect 32692 59812 32696 59868
rect 32696 59812 32752 59868
rect 32752 59812 32756 59868
rect 32692 59808 32756 59812
rect 32772 59868 32836 59872
rect 32772 59812 32776 59868
rect 32776 59812 32832 59868
rect 32832 59812 32836 59868
rect 32772 59808 32836 59812
rect 32852 59868 32916 59872
rect 32852 59812 32856 59868
rect 32856 59812 32912 59868
rect 32912 59812 32916 59868
rect 32852 59808 32916 59812
rect 37612 59868 37676 59872
rect 37612 59812 37616 59868
rect 37616 59812 37672 59868
rect 37672 59812 37676 59868
rect 37612 59808 37676 59812
rect 37692 59868 37756 59872
rect 37692 59812 37696 59868
rect 37696 59812 37752 59868
rect 37752 59812 37756 59868
rect 37692 59808 37756 59812
rect 37772 59868 37836 59872
rect 37772 59812 37776 59868
rect 37776 59812 37832 59868
rect 37832 59812 37836 59868
rect 37772 59808 37836 59812
rect 37852 59868 37916 59872
rect 37852 59812 37856 59868
rect 37856 59812 37912 59868
rect 37912 59812 37916 59868
rect 37852 59808 37916 59812
rect 1952 59324 2016 59328
rect 1952 59268 1956 59324
rect 1956 59268 2012 59324
rect 2012 59268 2016 59324
rect 1952 59264 2016 59268
rect 2032 59324 2096 59328
rect 2032 59268 2036 59324
rect 2036 59268 2092 59324
rect 2092 59268 2096 59324
rect 2032 59264 2096 59268
rect 2112 59324 2176 59328
rect 2112 59268 2116 59324
rect 2116 59268 2172 59324
rect 2172 59268 2176 59324
rect 2112 59264 2176 59268
rect 2192 59324 2256 59328
rect 2192 59268 2196 59324
rect 2196 59268 2252 59324
rect 2252 59268 2256 59324
rect 2192 59264 2256 59268
rect 6952 59324 7016 59328
rect 6952 59268 6956 59324
rect 6956 59268 7012 59324
rect 7012 59268 7016 59324
rect 6952 59264 7016 59268
rect 7032 59324 7096 59328
rect 7032 59268 7036 59324
rect 7036 59268 7092 59324
rect 7092 59268 7096 59324
rect 7032 59264 7096 59268
rect 7112 59324 7176 59328
rect 7112 59268 7116 59324
rect 7116 59268 7172 59324
rect 7172 59268 7176 59324
rect 7112 59264 7176 59268
rect 7192 59324 7256 59328
rect 7192 59268 7196 59324
rect 7196 59268 7252 59324
rect 7252 59268 7256 59324
rect 7192 59264 7256 59268
rect 11952 59324 12016 59328
rect 11952 59268 11956 59324
rect 11956 59268 12012 59324
rect 12012 59268 12016 59324
rect 11952 59264 12016 59268
rect 12032 59324 12096 59328
rect 12032 59268 12036 59324
rect 12036 59268 12092 59324
rect 12092 59268 12096 59324
rect 12032 59264 12096 59268
rect 12112 59324 12176 59328
rect 12112 59268 12116 59324
rect 12116 59268 12172 59324
rect 12172 59268 12176 59324
rect 12112 59264 12176 59268
rect 12192 59324 12256 59328
rect 12192 59268 12196 59324
rect 12196 59268 12252 59324
rect 12252 59268 12256 59324
rect 12192 59264 12256 59268
rect 16952 59324 17016 59328
rect 16952 59268 16956 59324
rect 16956 59268 17012 59324
rect 17012 59268 17016 59324
rect 16952 59264 17016 59268
rect 17032 59324 17096 59328
rect 17032 59268 17036 59324
rect 17036 59268 17092 59324
rect 17092 59268 17096 59324
rect 17032 59264 17096 59268
rect 17112 59324 17176 59328
rect 17112 59268 17116 59324
rect 17116 59268 17172 59324
rect 17172 59268 17176 59324
rect 17112 59264 17176 59268
rect 17192 59324 17256 59328
rect 17192 59268 17196 59324
rect 17196 59268 17252 59324
rect 17252 59268 17256 59324
rect 17192 59264 17256 59268
rect 21952 59324 22016 59328
rect 21952 59268 21956 59324
rect 21956 59268 22012 59324
rect 22012 59268 22016 59324
rect 21952 59264 22016 59268
rect 22032 59324 22096 59328
rect 22032 59268 22036 59324
rect 22036 59268 22092 59324
rect 22092 59268 22096 59324
rect 22032 59264 22096 59268
rect 22112 59324 22176 59328
rect 22112 59268 22116 59324
rect 22116 59268 22172 59324
rect 22172 59268 22176 59324
rect 22112 59264 22176 59268
rect 22192 59324 22256 59328
rect 22192 59268 22196 59324
rect 22196 59268 22252 59324
rect 22252 59268 22256 59324
rect 22192 59264 22256 59268
rect 26952 59324 27016 59328
rect 26952 59268 26956 59324
rect 26956 59268 27012 59324
rect 27012 59268 27016 59324
rect 26952 59264 27016 59268
rect 27032 59324 27096 59328
rect 27032 59268 27036 59324
rect 27036 59268 27092 59324
rect 27092 59268 27096 59324
rect 27032 59264 27096 59268
rect 27112 59324 27176 59328
rect 27112 59268 27116 59324
rect 27116 59268 27172 59324
rect 27172 59268 27176 59324
rect 27112 59264 27176 59268
rect 27192 59324 27256 59328
rect 27192 59268 27196 59324
rect 27196 59268 27252 59324
rect 27252 59268 27256 59324
rect 27192 59264 27256 59268
rect 31952 59324 32016 59328
rect 31952 59268 31956 59324
rect 31956 59268 32012 59324
rect 32012 59268 32016 59324
rect 31952 59264 32016 59268
rect 32032 59324 32096 59328
rect 32032 59268 32036 59324
rect 32036 59268 32092 59324
rect 32092 59268 32096 59324
rect 32032 59264 32096 59268
rect 32112 59324 32176 59328
rect 32112 59268 32116 59324
rect 32116 59268 32172 59324
rect 32172 59268 32176 59324
rect 32112 59264 32176 59268
rect 32192 59324 32256 59328
rect 32192 59268 32196 59324
rect 32196 59268 32252 59324
rect 32252 59268 32256 59324
rect 32192 59264 32256 59268
rect 36952 59324 37016 59328
rect 36952 59268 36956 59324
rect 36956 59268 37012 59324
rect 37012 59268 37016 59324
rect 36952 59264 37016 59268
rect 37032 59324 37096 59328
rect 37032 59268 37036 59324
rect 37036 59268 37092 59324
rect 37092 59268 37096 59324
rect 37032 59264 37096 59268
rect 37112 59324 37176 59328
rect 37112 59268 37116 59324
rect 37116 59268 37172 59324
rect 37172 59268 37176 59324
rect 37112 59264 37176 59268
rect 37192 59324 37256 59328
rect 37192 59268 37196 59324
rect 37196 59268 37252 59324
rect 37252 59268 37256 59324
rect 37192 59264 37256 59268
rect 2612 58780 2676 58784
rect 2612 58724 2616 58780
rect 2616 58724 2672 58780
rect 2672 58724 2676 58780
rect 2612 58720 2676 58724
rect 2692 58780 2756 58784
rect 2692 58724 2696 58780
rect 2696 58724 2752 58780
rect 2752 58724 2756 58780
rect 2692 58720 2756 58724
rect 2772 58780 2836 58784
rect 2772 58724 2776 58780
rect 2776 58724 2832 58780
rect 2832 58724 2836 58780
rect 2772 58720 2836 58724
rect 2852 58780 2916 58784
rect 2852 58724 2856 58780
rect 2856 58724 2912 58780
rect 2912 58724 2916 58780
rect 2852 58720 2916 58724
rect 7612 58780 7676 58784
rect 7612 58724 7616 58780
rect 7616 58724 7672 58780
rect 7672 58724 7676 58780
rect 7612 58720 7676 58724
rect 7692 58780 7756 58784
rect 7692 58724 7696 58780
rect 7696 58724 7752 58780
rect 7752 58724 7756 58780
rect 7692 58720 7756 58724
rect 7772 58780 7836 58784
rect 7772 58724 7776 58780
rect 7776 58724 7832 58780
rect 7832 58724 7836 58780
rect 7772 58720 7836 58724
rect 7852 58780 7916 58784
rect 7852 58724 7856 58780
rect 7856 58724 7912 58780
rect 7912 58724 7916 58780
rect 7852 58720 7916 58724
rect 12612 58780 12676 58784
rect 12612 58724 12616 58780
rect 12616 58724 12672 58780
rect 12672 58724 12676 58780
rect 12612 58720 12676 58724
rect 12692 58780 12756 58784
rect 12692 58724 12696 58780
rect 12696 58724 12752 58780
rect 12752 58724 12756 58780
rect 12692 58720 12756 58724
rect 12772 58780 12836 58784
rect 12772 58724 12776 58780
rect 12776 58724 12832 58780
rect 12832 58724 12836 58780
rect 12772 58720 12836 58724
rect 12852 58780 12916 58784
rect 12852 58724 12856 58780
rect 12856 58724 12912 58780
rect 12912 58724 12916 58780
rect 12852 58720 12916 58724
rect 17612 58780 17676 58784
rect 17612 58724 17616 58780
rect 17616 58724 17672 58780
rect 17672 58724 17676 58780
rect 17612 58720 17676 58724
rect 17692 58780 17756 58784
rect 17692 58724 17696 58780
rect 17696 58724 17752 58780
rect 17752 58724 17756 58780
rect 17692 58720 17756 58724
rect 17772 58780 17836 58784
rect 17772 58724 17776 58780
rect 17776 58724 17832 58780
rect 17832 58724 17836 58780
rect 17772 58720 17836 58724
rect 17852 58780 17916 58784
rect 17852 58724 17856 58780
rect 17856 58724 17912 58780
rect 17912 58724 17916 58780
rect 17852 58720 17916 58724
rect 22612 58780 22676 58784
rect 22612 58724 22616 58780
rect 22616 58724 22672 58780
rect 22672 58724 22676 58780
rect 22612 58720 22676 58724
rect 22692 58780 22756 58784
rect 22692 58724 22696 58780
rect 22696 58724 22752 58780
rect 22752 58724 22756 58780
rect 22692 58720 22756 58724
rect 22772 58780 22836 58784
rect 22772 58724 22776 58780
rect 22776 58724 22832 58780
rect 22832 58724 22836 58780
rect 22772 58720 22836 58724
rect 22852 58780 22916 58784
rect 22852 58724 22856 58780
rect 22856 58724 22912 58780
rect 22912 58724 22916 58780
rect 22852 58720 22916 58724
rect 27612 58780 27676 58784
rect 27612 58724 27616 58780
rect 27616 58724 27672 58780
rect 27672 58724 27676 58780
rect 27612 58720 27676 58724
rect 27692 58780 27756 58784
rect 27692 58724 27696 58780
rect 27696 58724 27752 58780
rect 27752 58724 27756 58780
rect 27692 58720 27756 58724
rect 27772 58780 27836 58784
rect 27772 58724 27776 58780
rect 27776 58724 27832 58780
rect 27832 58724 27836 58780
rect 27772 58720 27836 58724
rect 27852 58780 27916 58784
rect 27852 58724 27856 58780
rect 27856 58724 27912 58780
rect 27912 58724 27916 58780
rect 27852 58720 27916 58724
rect 32612 58780 32676 58784
rect 32612 58724 32616 58780
rect 32616 58724 32672 58780
rect 32672 58724 32676 58780
rect 32612 58720 32676 58724
rect 32692 58780 32756 58784
rect 32692 58724 32696 58780
rect 32696 58724 32752 58780
rect 32752 58724 32756 58780
rect 32692 58720 32756 58724
rect 32772 58780 32836 58784
rect 32772 58724 32776 58780
rect 32776 58724 32832 58780
rect 32832 58724 32836 58780
rect 32772 58720 32836 58724
rect 32852 58780 32916 58784
rect 32852 58724 32856 58780
rect 32856 58724 32912 58780
rect 32912 58724 32916 58780
rect 32852 58720 32916 58724
rect 37612 58780 37676 58784
rect 37612 58724 37616 58780
rect 37616 58724 37672 58780
rect 37672 58724 37676 58780
rect 37612 58720 37676 58724
rect 37692 58780 37756 58784
rect 37692 58724 37696 58780
rect 37696 58724 37752 58780
rect 37752 58724 37756 58780
rect 37692 58720 37756 58724
rect 37772 58780 37836 58784
rect 37772 58724 37776 58780
rect 37776 58724 37832 58780
rect 37832 58724 37836 58780
rect 37772 58720 37836 58724
rect 37852 58780 37916 58784
rect 37852 58724 37856 58780
rect 37856 58724 37912 58780
rect 37912 58724 37916 58780
rect 37852 58720 37916 58724
rect 33180 58304 33244 58308
rect 33180 58248 33230 58304
rect 33230 58248 33244 58304
rect 33180 58244 33244 58248
rect 1952 58236 2016 58240
rect 1952 58180 1956 58236
rect 1956 58180 2012 58236
rect 2012 58180 2016 58236
rect 1952 58176 2016 58180
rect 2032 58236 2096 58240
rect 2032 58180 2036 58236
rect 2036 58180 2092 58236
rect 2092 58180 2096 58236
rect 2032 58176 2096 58180
rect 2112 58236 2176 58240
rect 2112 58180 2116 58236
rect 2116 58180 2172 58236
rect 2172 58180 2176 58236
rect 2112 58176 2176 58180
rect 2192 58236 2256 58240
rect 2192 58180 2196 58236
rect 2196 58180 2252 58236
rect 2252 58180 2256 58236
rect 2192 58176 2256 58180
rect 6952 58236 7016 58240
rect 6952 58180 6956 58236
rect 6956 58180 7012 58236
rect 7012 58180 7016 58236
rect 6952 58176 7016 58180
rect 7032 58236 7096 58240
rect 7032 58180 7036 58236
rect 7036 58180 7092 58236
rect 7092 58180 7096 58236
rect 7032 58176 7096 58180
rect 7112 58236 7176 58240
rect 7112 58180 7116 58236
rect 7116 58180 7172 58236
rect 7172 58180 7176 58236
rect 7112 58176 7176 58180
rect 7192 58236 7256 58240
rect 7192 58180 7196 58236
rect 7196 58180 7252 58236
rect 7252 58180 7256 58236
rect 7192 58176 7256 58180
rect 11952 58236 12016 58240
rect 11952 58180 11956 58236
rect 11956 58180 12012 58236
rect 12012 58180 12016 58236
rect 11952 58176 12016 58180
rect 12032 58236 12096 58240
rect 12032 58180 12036 58236
rect 12036 58180 12092 58236
rect 12092 58180 12096 58236
rect 12032 58176 12096 58180
rect 12112 58236 12176 58240
rect 12112 58180 12116 58236
rect 12116 58180 12172 58236
rect 12172 58180 12176 58236
rect 12112 58176 12176 58180
rect 12192 58236 12256 58240
rect 12192 58180 12196 58236
rect 12196 58180 12252 58236
rect 12252 58180 12256 58236
rect 12192 58176 12256 58180
rect 16952 58236 17016 58240
rect 16952 58180 16956 58236
rect 16956 58180 17012 58236
rect 17012 58180 17016 58236
rect 16952 58176 17016 58180
rect 17032 58236 17096 58240
rect 17032 58180 17036 58236
rect 17036 58180 17092 58236
rect 17092 58180 17096 58236
rect 17032 58176 17096 58180
rect 17112 58236 17176 58240
rect 17112 58180 17116 58236
rect 17116 58180 17172 58236
rect 17172 58180 17176 58236
rect 17112 58176 17176 58180
rect 17192 58236 17256 58240
rect 17192 58180 17196 58236
rect 17196 58180 17252 58236
rect 17252 58180 17256 58236
rect 17192 58176 17256 58180
rect 21952 58236 22016 58240
rect 21952 58180 21956 58236
rect 21956 58180 22012 58236
rect 22012 58180 22016 58236
rect 21952 58176 22016 58180
rect 22032 58236 22096 58240
rect 22032 58180 22036 58236
rect 22036 58180 22092 58236
rect 22092 58180 22096 58236
rect 22032 58176 22096 58180
rect 22112 58236 22176 58240
rect 22112 58180 22116 58236
rect 22116 58180 22172 58236
rect 22172 58180 22176 58236
rect 22112 58176 22176 58180
rect 22192 58236 22256 58240
rect 22192 58180 22196 58236
rect 22196 58180 22252 58236
rect 22252 58180 22256 58236
rect 22192 58176 22256 58180
rect 26952 58236 27016 58240
rect 26952 58180 26956 58236
rect 26956 58180 27012 58236
rect 27012 58180 27016 58236
rect 26952 58176 27016 58180
rect 27032 58236 27096 58240
rect 27032 58180 27036 58236
rect 27036 58180 27092 58236
rect 27092 58180 27096 58236
rect 27032 58176 27096 58180
rect 27112 58236 27176 58240
rect 27112 58180 27116 58236
rect 27116 58180 27172 58236
rect 27172 58180 27176 58236
rect 27112 58176 27176 58180
rect 27192 58236 27256 58240
rect 27192 58180 27196 58236
rect 27196 58180 27252 58236
rect 27252 58180 27256 58236
rect 27192 58176 27256 58180
rect 31952 58236 32016 58240
rect 31952 58180 31956 58236
rect 31956 58180 32012 58236
rect 32012 58180 32016 58236
rect 31952 58176 32016 58180
rect 32032 58236 32096 58240
rect 32032 58180 32036 58236
rect 32036 58180 32092 58236
rect 32092 58180 32096 58236
rect 32032 58176 32096 58180
rect 32112 58236 32176 58240
rect 32112 58180 32116 58236
rect 32116 58180 32172 58236
rect 32172 58180 32176 58236
rect 32112 58176 32176 58180
rect 32192 58236 32256 58240
rect 32192 58180 32196 58236
rect 32196 58180 32252 58236
rect 32252 58180 32256 58236
rect 32192 58176 32256 58180
rect 36952 58236 37016 58240
rect 36952 58180 36956 58236
rect 36956 58180 37012 58236
rect 37012 58180 37016 58236
rect 36952 58176 37016 58180
rect 37032 58236 37096 58240
rect 37032 58180 37036 58236
rect 37036 58180 37092 58236
rect 37092 58180 37096 58236
rect 37032 58176 37096 58180
rect 37112 58236 37176 58240
rect 37112 58180 37116 58236
rect 37116 58180 37172 58236
rect 37172 58180 37176 58236
rect 37112 58176 37176 58180
rect 37192 58236 37256 58240
rect 37192 58180 37196 58236
rect 37196 58180 37252 58236
rect 37252 58180 37256 58236
rect 37192 58176 37256 58180
rect 2612 57692 2676 57696
rect 2612 57636 2616 57692
rect 2616 57636 2672 57692
rect 2672 57636 2676 57692
rect 2612 57632 2676 57636
rect 2692 57692 2756 57696
rect 2692 57636 2696 57692
rect 2696 57636 2752 57692
rect 2752 57636 2756 57692
rect 2692 57632 2756 57636
rect 2772 57692 2836 57696
rect 2772 57636 2776 57692
rect 2776 57636 2832 57692
rect 2832 57636 2836 57692
rect 2772 57632 2836 57636
rect 2852 57692 2916 57696
rect 2852 57636 2856 57692
rect 2856 57636 2912 57692
rect 2912 57636 2916 57692
rect 2852 57632 2916 57636
rect 7612 57692 7676 57696
rect 7612 57636 7616 57692
rect 7616 57636 7672 57692
rect 7672 57636 7676 57692
rect 7612 57632 7676 57636
rect 7692 57692 7756 57696
rect 7692 57636 7696 57692
rect 7696 57636 7752 57692
rect 7752 57636 7756 57692
rect 7692 57632 7756 57636
rect 7772 57692 7836 57696
rect 7772 57636 7776 57692
rect 7776 57636 7832 57692
rect 7832 57636 7836 57692
rect 7772 57632 7836 57636
rect 7852 57692 7916 57696
rect 7852 57636 7856 57692
rect 7856 57636 7912 57692
rect 7912 57636 7916 57692
rect 7852 57632 7916 57636
rect 12612 57692 12676 57696
rect 12612 57636 12616 57692
rect 12616 57636 12672 57692
rect 12672 57636 12676 57692
rect 12612 57632 12676 57636
rect 12692 57692 12756 57696
rect 12692 57636 12696 57692
rect 12696 57636 12752 57692
rect 12752 57636 12756 57692
rect 12692 57632 12756 57636
rect 12772 57692 12836 57696
rect 12772 57636 12776 57692
rect 12776 57636 12832 57692
rect 12832 57636 12836 57692
rect 12772 57632 12836 57636
rect 12852 57692 12916 57696
rect 12852 57636 12856 57692
rect 12856 57636 12912 57692
rect 12912 57636 12916 57692
rect 12852 57632 12916 57636
rect 17612 57692 17676 57696
rect 17612 57636 17616 57692
rect 17616 57636 17672 57692
rect 17672 57636 17676 57692
rect 17612 57632 17676 57636
rect 17692 57692 17756 57696
rect 17692 57636 17696 57692
rect 17696 57636 17752 57692
rect 17752 57636 17756 57692
rect 17692 57632 17756 57636
rect 17772 57692 17836 57696
rect 17772 57636 17776 57692
rect 17776 57636 17832 57692
rect 17832 57636 17836 57692
rect 17772 57632 17836 57636
rect 17852 57692 17916 57696
rect 17852 57636 17856 57692
rect 17856 57636 17912 57692
rect 17912 57636 17916 57692
rect 17852 57632 17916 57636
rect 22612 57692 22676 57696
rect 22612 57636 22616 57692
rect 22616 57636 22672 57692
rect 22672 57636 22676 57692
rect 22612 57632 22676 57636
rect 22692 57692 22756 57696
rect 22692 57636 22696 57692
rect 22696 57636 22752 57692
rect 22752 57636 22756 57692
rect 22692 57632 22756 57636
rect 22772 57692 22836 57696
rect 22772 57636 22776 57692
rect 22776 57636 22832 57692
rect 22832 57636 22836 57692
rect 22772 57632 22836 57636
rect 22852 57692 22916 57696
rect 22852 57636 22856 57692
rect 22856 57636 22912 57692
rect 22912 57636 22916 57692
rect 22852 57632 22916 57636
rect 27612 57692 27676 57696
rect 27612 57636 27616 57692
rect 27616 57636 27672 57692
rect 27672 57636 27676 57692
rect 27612 57632 27676 57636
rect 27692 57692 27756 57696
rect 27692 57636 27696 57692
rect 27696 57636 27752 57692
rect 27752 57636 27756 57692
rect 27692 57632 27756 57636
rect 27772 57692 27836 57696
rect 27772 57636 27776 57692
rect 27776 57636 27832 57692
rect 27832 57636 27836 57692
rect 27772 57632 27836 57636
rect 27852 57692 27916 57696
rect 27852 57636 27856 57692
rect 27856 57636 27912 57692
rect 27912 57636 27916 57692
rect 27852 57632 27916 57636
rect 32612 57692 32676 57696
rect 32612 57636 32616 57692
rect 32616 57636 32672 57692
rect 32672 57636 32676 57692
rect 32612 57632 32676 57636
rect 32692 57692 32756 57696
rect 32692 57636 32696 57692
rect 32696 57636 32752 57692
rect 32752 57636 32756 57692
rect 32692 57632 32756 57636
rect 32772 57692 32836 57696
rect 32772 57636 32776 57692
rect 32776 57636 32832 57692
rect 32832 57636 32836 57692
rect 32772 57632 32836 57636
rect 32852 57692 32916 57696
rect 32852 57636 32856 57692
rect 32856 57636 32912 57692
rect 32912 57636 32916 57692
rect 32852 57632 32916 57636
rect 37612 57692 37676 57696
rect 37612 57636 37616 57692
rect 37616 57636 37672 57692
rect 37672 57636 37676 57692
rect 37612 57632 37676 57636
rect 37692 57692 37756 57696
rect 37692 57636 37696 57692
rect 37696 57636 37752 57692
rect 37752 57636 37756 57692
rect 37692 57632 37756 57636
rect 37772 57692 37836 57696
rect 37772 57636 37776 57692
rect 37776 57636 37832 57692
rect 37832 57636 37836 57692
rect 37772 57632 37836 57636
rect 37852 57692 37916 57696
rect 37852 57636 37856 57692
rect 37856 57636 37912 57692
rect 37912 57636 37916 57692
rect 37852 57632 37916 57636
rect 1952 57148 2016 57152
rect 1952 57092 1956 57148
rect 1956 57092 2012 57148
rect 2012 57092 2016 57148
rect 1952 57088 2016 57092
rect 2032 57148 2096 57152
rect 2032 57092 2036 57148
rect 2036 57092 2092 57148
rect 2092 57092 2096 57148
rect 2032 57088 2096 57092
rect 2112 57148 2176 57152
rect 2112 57092 2116 57148
rect 2116 57092 2172 57148
rect 2172 57092 2176 57148
rect 2112 57088 2176 57092
rect 2192 57148 2256 57152
rect 2192 57092 2196 57148
rect 2196 57092 2252 57148
rect 2252 57092 2256 57148
rect 2192 57088 2256 57092
rect 6952 57148 7016 57152
rect 6952 57092 6956 57148
rect 6956 57092 7012 57148
rect 7012 57092 7016 57148
rect 6952 57088 7016 57092
rect 7032 57148 7096 57152
rect 7032 57092 7036 57148
rect 7036 57092 7092 57148
rect 7092 57092 7096 57148
rect 7032 57088 7096 57092
rect 7112 57148 7176 57152
rect 7112 57092 7116 57148
rect 7116 57092 7172 57148
rect 7172 57092 7176 57148
rect 7112 57088 7176 57092
rect 7192 57148 7256 57152
rect 7192 57092 7196 57148
rect 7196 57092 7252 57148
rect 7252 57092 7256 57148
rect 7192 57088 7256 57092
rect 11952 57148 12016 57152
rect 11952 57092 11956 57148
rect 11956 57092 12012 57148
rect 12012 57092 12016 57148
rect 11952 57088 12016 57092
rect 12032 57148 12096 57152
rect 12032 57092 12036 57148
rect 12036 57092 12092 57148
rect 12092 57092 12096 57148
rect 12032 57088 12096 57092
rect 12112 57148 12176 57152
rect 12112 57092 12116 57148
rect 12116 57092 12172 57148
rect 12172 57092 12176 57148
rect 12112 57088 12176 57092
rect 12192 57148 12256 57152
rect 12192 57092 12196 57148
rect 12196 57092 12252 57148
rect 12252 57092 12256 57148
rect 12192 57088 12256 57092
rect 16952 57148 17016 57152
rect 16952 57092 16956 57148
rect 16956 57092 17012 57148
rect 17012 57092 17016 57148
rect 16952 57088 17016 57092
rect 17032 57148 17096 57152
rect 17032 57092 17036 57148
rect 17036 57092 17092 57148
rect 17092 57092 17096 57148
rect 17032 57088 17096 57092
rect 17112 57148 17176 57152
rect 17112 57092 17116 57148
rect 17116 57092 17172 57148
rect 17172 57092 17176 57148
rect 17112 57088 17176 57092
rect 17192 57148 17256 57152
rect 17192 57092 17196 57148
rect 17196 57092 17252 57148
rect 17252 57092 17256 57148
rect 17192 57088 17256 57092
rect 21952 57148 22016 57152
rect 21952 57092 21956 57148
rect 21956 57092 22012 57148
rect 22012 57092 22016 57148
rect 21952 57088 22016 57092
rect 22032 57148 22096 57152
rect 22032 57092 22036 57148
rect 22036 57092 22092 57148
rect 22092 57092 22096 57148
rect 22032 57088 22096 57092
rect 22112 57148 22176 57152
rect 22112 57092 22116 57148
rect 22116 57092 22172 57148
rect 22172 57092 22176 57148
rect 22112 57088 22176 57092
rect 22192 57148 22256 57152
rect 22192 57092 22196 57148
rect 22196 57092 22252 57148
rect 22252 57092 22256 57148
rect 22192 57088 22256 57092
rect 26952 57148 27016 57152
rect 26952 57092 26956 57148
rect 26956 57092 27012 57148
rect 27012 57092 27016 57148
rect 26952 57088 27016 57092
rect 27032 57148 27096 57152
rect 27032 57092 27036 57148
rect 27036 57092 27092 57148
rect 27092 57092 27096 57148
rect 27032 57088 27096 57092
rect 27112 57148 27176 57152
rect 27112 57092 27116 57148
rect 27116 57092 27172 57148
rect 27172 57092 27176 57148
rect 27112 57088 27176 57092
rect 27192 57148 27256 57152
rect 27192 57092 27196 57148
rect 27196 57092 27252 57148
rect 27252 57092 27256 57148
rect 27192 57088 27256 57092
rect 31952 57148 32016 57152
rect 31952 57092 31956 57148
rect 31956 57092 32012 57148
rect 32012 57092 32016 57148
rect 31952 57088 32016 57092
rect 32032 57148 32096 57152
rect 32032 57092 32036 57148
rect 32036 57092 32092 57148
rect 32092 57092 32096 57148
rect 32032 57088 32096 57092
rect 32112 57148 32176 57152
rect 32112 57092 32116 57148
rect 32116 57092 32172 57148
rect 32172 57092 32176 57148
rect 32112 57088 32176 57092
rect 32192 57148 32256 57152
rect 32192 57092 32196 57148
rect 32196 57092 32252 57148
rect 32252 57092 32256 57148
rect 32192 57088 32256 57092
rect 36952 57148 37016 57152
rect 36952 57092 36956 57148
rect 36956 57092 37012 57148
rect 37012 57092 37016 57148
rect 36952 57088 37016 57092
rect 37032 57148 37096 57152
rect 37032 57092 37036 57148
rect 37036 57092 37092 57148
rect 37092 57092 37096 57148
rect 37032 57088 37096 57092
rect 37112 57148 37176 57152
rect 37112 57092 37116 57148
rect 37116 57092 37172 57148
rect 37172 57092 37176 57148
rect 37112 57088 37176 57092
rect 37192 57148 37256 57152
rect 37192 57092 37196 57148
rect 37196 57092 37252 57148
rect 37252 57092 37256 57148
rect 37192 57088 37256 57092
rect 2612 56604 2676 56608
rect 2612 56548 2616 56604
rect 2616 56548 2672 56604
rect 2672 56548 2676 56604
rect 2612 56544 2676 56548
rect 2692 56604 2756 56608
rect 2692 56548 2696 56604
rect 2696 56548 2752 56604
rect 2752 56548 2756 56604
rect 2692 56544 2756 56548
rect 2772 56604 2836 56608
rect 2772 56548 2776 56604
rect 2776 56548 2832 56604
rect 2832 56548 2836 56604
rect 2772 56544 2836 56548
rect 2852 56604 2916 56608
rect 2852 56548 2856 56604
rect 2856 56548 2912 56604
rect 2912 56548 2916 56604
rect 2852 56544 2916 56548
rect 7612 56604 7676 56608
rect 7612 56548 7616 56604
rect 7616 56548 7672 56604
rect 7672 56548 7676 56604
rect 7612 56544 7676 56548
rect 7692 56604 7756 56608
rect 7692 56548 7696 56604
rect 7696 56548 7752 56604
rect 7752 56548 7756 56604
rect 7692 56544 7756 56548
rect 7772 56604 7836 56608
rect 7772 56548 7776 56604
rect 7776 56548 7832 56604
rect 7832 56548 7836 56604
rect 7772 56544 7836 56548
rect 7852 56604 7916 56608
rect 7852 56548 7856 56604
rect 7856 56548 7912 56604
rect 7912 56548 7916 56604
rect 7852 56544 7916 56548
rect 12612 56604 12676 56608
rect 12612 56548 12616 56604
rect 12616 56548 12672 56604
rect 12672 56548 12676 56604
rect 12612 56544 12676 56548
rect 12692 56604 12756 56608
rect 12692 56548 12696 56604
rect 12696 56548 12752 56604
rect 12752 56548 12756 56604
rect 12692 56544 12756 56548
rect 12772 56604 12836 56608
rect 12772 56548 12776 56604
rect 12776 56548 12832 56604
rect 12832 56548 12836 56604
rect 12772 56544 12836 56548
rect 12852 56604 12916 56608
rect 12852 56548 12856 56604
rect 12856 56548 12912 56604
rect 12912 56548 12916 56604
rect 12852 56544 12916 56548
rect 17612 56604 17676 56608
rect 17612 56548 17616 56604
rect 17616 56548 17672 56604
rect 17672 56548 17676 56604
rect 17612 56544 17676 56548
rect 17692 56604 17756 56608
rect 17692 56548 17696 56604
rect 17696 56548 17752 56604
rect 17752 56548 17756 56604
rect 17692 56544 17756 56548
rect 17772 56604 17836 56608
rect 17772 56548 17776 56604
rect 17776 56548 17832 56604
rect 17832 56548 17836 56604
rect 17772 56544 17836 56548
rect 17852 56604 17916 56608
rect 17852 56548 17856 56604
rect 17856 56548 17912 56604
rect 17912 56548 17916 56604
rect 17852 56544 17916 56548
rect 22612 56604 22676 56608
rect 22612 56548 22616 56604
rect 22616 56548 22672 56604
rect 22672 56548 22676 56604
rect 22612 56544 22676 56548
rect 22692 56604 22756 56608
rect 22692 56548 22696 56604
rect 22696 56548 22752 56604
rect 22752 56548 22756 56604
rect 22692 56544 22756 56548
rect 22772 56604 22836 56608
rect 22772 56548 22776 56604
rect 22776 56548 22832 56604
rect 22832 56548 22836 56604
rect 22772 56544 22836 56548
rect 22852 56604 22916 56608
rect 22852 56548 22856 56604
rect 22856 56548 22912 56604
rect 22912 56548 22916 56604
rect 22852 56544 22916 56548
rect 27612 56604 27676 56608
rect 27612 56548 27616 56604
rect 27616 56548 27672 56604
rect 27672 56548 27676 56604
rect 27612 56544 27676 56548
rect 27692 56604 27756 56608
rect 27692 56548 27696 56604
rect 27696 56548 27752 56604
rect 27752 56548 27756 56604
rect 27692 56544 27756 56548
rect 27772 56604 27836 56608
rect 27772 56548 27776 56604
rect 27776 56548 27832 56604
rect 27832 56548 27836 56604
rect 27772 56544 27836 56548
rect 27852 56604 27916 56608
rect 27852 56548 27856 56604
rect 27856 56548 27912 56604
rect 27912 56548 27916 56604
rect 27852 56544 27916 56548
rect 32612 56604 32676 56608
rect 32612 56548 32616 56604
rect 32616 56548 32672 56604
rect 32672 56548 32676 56604
rect 32612 56544 32676 56548
rect 32692 56604 32756 56608
rect 32692 56548 32696 56604
rect 32696 56548 32752 56604
rect 32752 56548 32756 56604
rect 32692 56544 32756 56548
rect 32772 56604 32836 56608
rect 32772 56548 32776 56604
rect 32776 56548 32832 56604
rect 32832 56548 32836 56604
rect 32772 56544 32836 56548
rect 32852 56604 32916 56608
rect 32852 56548 32856 56604
rect 32856 56548 32912 56604
rect 32912 56548 32916 56604
rect 32852 56544 32916 56548
rect 37612 56604 37676 56608
rect 37612 56548 37616 56604
rect 37616 56548 37672 56604
rect 37672 56548 37676 56604
rect 37612 56544 37676 56548
rect 37692 56604 37756 56608
rect 37692 56548 37696 56604
rect 37696 56548 37752 56604
rect 37752 56548 37756 56604
rect 37692 56544 37756 56548
rect 37772 56604 37836 56608
rect 37772 56548 37776 56604
rect 37776 56548 37832 56604
rect 37832 56548 37836 56604
rect 37772 56544 37836 56548
rect 37852 56604 37916 56608
rect 37852 56548 37856 56604
rect 37856 56548 37912 56604
rect 37912 56548 37916 56604
rect 37852 56544 37916 56548
rect 1952 56060 2016 56064
rect 1952 56004 1956 56060
rect 1956 56004 2012 56060
rect 2012 56004 2016 56060
rect 1952 56000 2016 56004
rect 2032 56060 2096 56064
rect 2032 56004 2036 56060
rect 2036 56004 2092 56060
rect 2092 56004 2096 56060
rect 2032 56000 2096 56004
rect 2112 56060 2176 56064
rect 2112 56004 2116 56060
rect 2116 56004 2172 56060
rect 2172 56004 2176 56060
rect 2112 56000 2176 56004
rect 2192 56060 2256 56064
rect 2192 56004 2196 56060
rect 2196 56004 2252 56060
rect 2252 56004 2256 56060
rect 2192 56000 2256 56004
rect 6952 56060 7016 56064
rect 6952 56004 6956 56060
rect 6956 56004 7012 56060
rect 7012 56004 7016 56060
rect 6952 56000 7016 56004
rect 7032 56060 7096 56064
rect 7032 56004 7036 56060
rect 7036 56004 7092 56060
rect 7092 56004 7096 56060
rect 7032 56000 7096 56004
rect 7112 56060 7176 56064
rect 7112 56004 7116 56060
rect 7116 56004 7172 56060
rect 7172 56004 7176 56060
rect 7112 56000 7176 56004
rect 7192 56060 7256 56064
rect 7192 56004 7196 56060
rect 7196 56004 7252 56060
rect 7252 56004 7256 56060
rect 7192 56000 7256 56004
rect 11952 56060 12016 56064
rect 11952 56004 11956 56060
rect 11956 56004 12012 56060
rect 12012 56004 12016 56060
rect 11952 56000 12016 56004
rect 12032 56060 12096 56064
rect 12032 56004 12036 56060
rect 12036 56004 12092 56060
rect 12092 56004 12096 56060
rect 12032 56000 12096 56004
rect 12112 56060 12176 56064
rect 12112 56004 12116 56060
rect 12116 56004 12172 56060
rect 12172 56004 12176 56060
rect 12112 56000 12176 56004
rect 12192 56060 12256 56064
rect 12192 56004 12196 56060
rect 12196 56004 12252 56060
rect 12252 56004 12256 56060
rect 12192 56000 12256 56004
rect 16952 56060 17016 56064
rect 16952 56004 16956 56060
rect 16956 56004 17012 56060
rect 17012 56004 17016 56060
rect 16952 56000 17016 56004
rect 17032 56060 17096 56064
rect 17032 56004 17036 56060
rect 17036 56004 17092 56060
rect 17092 56004 17096 56060
rect 17032 56000 17096 56004
rect 17112 56060 17176 56064
rect 17112 56004 17116 56060
rect 17116 56004 17172 56060
rect 17172 56004 17176 56060
rect 17112 56000 17176 56004
rect 17192 56060 17256 56064
rect 17192 56004 17196 56060
rect 17196 56004 17252 56060
rect 17252 56004 17256 56060
rect 17192 56000 17256 56004
rect 21952 56060 22016 56064
rect 21952 56004 21956 56060
rect 21956 56004 22012 56060
rect 22012 56004 22016 56060
rect 21952 56000 22016 56004
rect 22032 56060 22096 56064
rect 22032 56004 22036 56060
rect 22036 56004 22092 56060
rect 22092 56004 22096 56060
rect 22032 56000 22096 56004
rect 22112 56060 22176 56064
rect 22112 56004 22116 56060
rect 22116 56004 22172 56060
rect 22172 56004 22176 56060
rect 22112 56000 22176 56004
rect 22192 56060 22256 56064
rect 22192 56004 22196 56060
rect 22196 56004 22252 56060
rect 22252 56004 22256 56060
rect 22192 56000 22256 56004
rect 26952 56060 27016 56064
rect 26952 56004 26956 56060
rect 26956 56004 27012 56060
rect 27012 56004 27016 56060
rect 26952 56000 27016 56004
rect 27032 56060 27096 56064
rect 27032 56004 27036 56060
rect 27036 56004 27092 56060
rect 27092 56004 27096 56060
rect 27032 56000 27096 56004
rect 27112 56060 27176 56064
rect 27112 56004 27116 56060
rect 27116 56004 27172 56060
rect 27172 56004 27176 56060
rect 27112 56000 27176 56004
rect 27192 56060 27256 56064
rect 27192 56004 27196 56060
rect 27196 56004 27252 56060
rect 27252 56004 27256 56060
rect 27192 56000 27256 56004
rect 31952 56060 32016 56064
rect 31952 56004 31956 56060
rect 31956 56004 32012 56060
rect 32012 56004 32016 56060
rect 31952 56000 32016 56004
rect 32032 56060 32096 56064
rect 32032 56004 32036 56060
rect 32036 56004 32092 56060
rect 32092 56004 32096 56060
rect 32032 56000 32096 56004
rect 32112 56060 32176 56064
rect 32112 56004 32116 56060
rect 32116 56004 32172 56060
rect 32172 56004 32176 56060
rect 32112 56000 32176 56004
rect 32192 56060 32256 56064
rect 32192 56004 32196 56060
rect 32196 56004 32252 56060
rect 32252 56004 32256 56060
rect 32192 56000 32256 56004
rect 36952 56060 37016 56064
rect 36952 56004 36956 56060
rect 36956 56004 37012 56060
rect 37012 56004 37016 56060
rect 36952 56000 37016 56004
rect 37032 56060 37096 56064
rect 37032 56004 37036 56060
rect 37036 56004 37092 56060
rect 37092 56004 37096 56060
rect 37032 56000 37096 56004
rect 37112 56060 37176 56064
rect 37112 56004 37116 56060
rect 37116 56004 37172 56060
rect 37172 56004 37176 56060
rect 37112 56000 37176 56004
rect 37192 56060 37256 56064
rect 37192 56004 37196 56060
rect 37196 56004 37252 56060
rect 37252 56004 37256 56060
rect 37192 56000 37256 56004
rect 33916 55856 33980 55860
rect 33916 55800 33930 55856
rect 33930 55800 33980 55856
rect 33916 55796 33980 55800
rect 33548 55720 33612 55724
rect 33548 55664 33562 55720
rect 33562 55664 33612 55720
rect 33548 55660 33612 55664
rect 2612 55516 2676 55520
rect 2612 55460 2616 55516
rect 2616 55460 2672 55516
rect 2672 55460 2676 55516
rect 2612 55456 2676 55460
rect 2692 55516 2756 55520
rect 2692 55460 2696 55516
rect 2696 55460 2752 55516
rect 2752 55460 2756 55516
rect 2692 55456 2756 55460
rect 2772 55516 2836 55520
rect 2772 55460 2776 55516
rect 2776 55460 2832 55516
rect 2832 55460 2836 55516
rect 2772 55456 2836 55460
rect 2852 55516 2916 55520
rect 2852 55460 2856 55516
rect 2856 55460 2912 55516
rect 2912 55460 2916 55516
rect 2852 55456 2916 55460
rect 7612 55516 7676 55520
rect 7612 55460 7616 55516
rect 7616 55460 7672 55516
rect 7672 55460 7676 55516
rect 7612 55456 7676 55460
rect 7692 55516 7756 55520
rect 7692 55460 7696 55516
rect 7696 55460 7752 55516
rect 7752 55460 7756 55516
rect 7692 55456 7756 55460
rect 7772 55516 7836 55520
rect 7772 55460 7776 55516
rect 7776 55460 7832 55516
rect 7832 55460 7836 55516
rect 7772 55456 7836 55460
rect 7852 55516 7916 55520
rect 7852 55460 7856 55516
rect 7856 55460 7912 55516
rect 7912 55460 7916 55516
rect 7852 55456 7916 55460
rect 12612 55516 12676 55520
rect 12612 55460 12616 55516
rect 12616 55460 12672 55516
rect 12672 55460 12676 55516
rect 12612 55456 12676 55460
rect 12692 55516 12756 55520
rect 12692 55460 12696 55516
rect 12696 55460 12752 55516
rect 12752 55460 12756 55516
rect 12692 55456 12756 55460
rect 12772 55516 12836 55520
rect 12772 55460 12776 55516
rect 12776 55460 12832 55516
rect 12832 55460 12836 55516
rect 12772 55456 12836 55460
rect 12852 55516 12916 55520
rect 12852 55460 12856 55516
rect 12856 55460 12912 55516
rect 12912 55460 12916 55516
rect 12852 55456 12916 55460
rect 17612 55516 17676 55520
rect 17612 55460 17616 55516
rect 17616 55460 17672 55516
rect 17672 55460 17676 55516
rect 17612 55456 17676 55460
rect 17692 55516 17756 55520
rect 17692 55460 17696 55516
rect 17696 55460 17752 55516
rect 17752 55460 17756 55516
rect 17692 55456 17756 55460
rect 17772 55516 17836 55520
rect 17772 55460 17776 55516
rect 17776 55460 17832 55516
rect 17832 55460 17836 55516
rect 17772 55456 17836 55460
rect 17852 55516 17916 55520
rect 17852 55460 17856 55516
rect 17856 55460 17912 55516
rect 17912 55460 17916 55516
rect 17852 55456 17916 55460
rect 22612 55516 22676 55520
rect 22612 55460 22616 55516
rect 22616 55460 22672 55516
rect 22672 55460 22676 55516
rect 22612 55456 22676 55460
rect 22692 55516 22756 55520
rect 22692 55460 22696 55516
rect 22696 55460 22752 55516
rect 22752 55460 22756 55516
rect 22692 55456 22756 55460
rect 22772 55516 22836 55520
rect 22772 55460 22776 55516
rect 22776 55460 22832 55516
rect 22832 55460 22836 55516
rect 22772 55456 22836 55460
rect 22852 55516 22916 55520
rect 22852 55460 22856 55516
rect 22856 55460 22912 55516
rect 22912 55460 22916 55516
rect 22852 55456 22916 55460
rect 27612 55516 27676 55520
rect 27612 55460 27616 55516
rect 27616 55460 27672 55516
rect 27672 55460 27676 55516
rect 27612 55456 27676 55460
rect 27692 55516 27756 55520
rect 27692 55460 27696 55516
rect 27696 55460 27752 55516
rect 27752 55460 27756 55516
rect 27692 55456 27756 55460
rect 27772 55516 27836 55520
rect 27772 55460 27776 55516
rect 27776 55460 27832 55516
rect 27832 55460 27836 55516
rect 27772 55456 27836 55460
rect 27852 55516 27916 55520
rect 27852 55460 27856 55516
rect 27856 55460 27912 55516
rect 27912 55460 27916 55516
rect 27852 55456 27916 55460
rect 32612 55516 32676 55520
rect 32612 55460 32616 55516
rect 32616 55460 32672 55516
rect 32672 55460 32676 55516
rect 32612 55456 32676 55460
rect 32692 55516 32756 55520
rect 32692 55460 32696 55516
rect 32696 55460 32752 55516
rect 32752 55460 32756 55516
rect 32692 55456 32756 55460
rect 32772 55516 32836 55520
rect 32772 55460 32776 55516
rect 32776 55460 32832 55516
rect 32832 55460 32836 55516
rect 32772 55456 32836 55460
rect 32852 55516 32916 55520
rect 32852 55460 32856 55516
rect 32856 55460 32912 55516
rect 32912 55460 32916 55516
rect 32852 55456 32916 55460
rect 37612 55516 37676 55520
rect 37612 55460 37616 55516
rect 37616 55460 37672 55516
rect 37672 55460 37676 55516
rect 37612 55456 37676 55460
rect 37692 55516 37756 55520
rect 37692 55460 37696 55516
rect 37696 55460 37752 55516
rect 37752 55460 37756 55516
rect 37692 55456 37756 55460
rect 37772 55516 37836 55520
rect 37772 55460 37776 55516
rect 37776 55460 37832 55516
rect 37832 55460 37836 55516
rect 37772 55456 37836 55460
rect 37852 55516 37916 55520
rect 37852 55460 37856 55516
rect 37856 55460 37912 55516
rect 37912 55460 37916 55516
rect 37852 55456 37916 55460
rect 1952 54972 2016 54976
rect 1952 54916 1956 54972
rect 1956 54916 2012 54972
rect 2012 54916 2016 54972
rect 1952 54912 2016 54916
rect 2032 54972 2096 54976
rect 2032 54916 2036 54972
rect 2036 54916 2092 54972
rect 2092 54916 2096 54972
rect 2032 54912 2096 54916
rect 2112 54972 2176 54976
rect 2112 54916 2116 54972
rect 2116 54916 2172 54972
rect 2172 54916 2176 54972
rect 2112 54912 2176 54916
rect 2192 54972 2256 54976
rect 2192 54916 2196 54972
rect 2196 54916 2252 54972
rect 2252 54916 2256 54972
rect 2192 54912 2256 54916
rect 6952 54972 7016 54976
rect 6952 54916 6956 54972
rect 6956 54916 7012 54972
rect 7012 54916 7016 54972
rect 6952 54912 7016 54916
rect 7032 54972 7096 54976
rect 7032 54916 7036 54972
rect 7036 54916 7092 54972
rect 7092 54916 7096 54972
rect 7032 54912 7096 54916
rect 7112 54972 7176 54976
rect 7112 54916 7116 54972
rect 7116 54916 7172 54972
rect 7172 54916 7176 54972
rect 7112 54912 7176 54916
rect 7192 54972 7256 54976
rect 7192 54916 7196 54972
rect 7196 54916 7252 54972
rect 7252 54916 7256 54972
rect 7192 54912 7256 54916
rect 11952 54972 12016 54976
rect 11952 54916 11956 54972
rect 11956 54916 12012 54972
rect 12012 54916 12016 54972
rect 11952 54912 12016 54916
rect 12032 54972 12096 54976
rect 12032 54916 12036 54972
rect 12036 54916 12092 54972
rect 12092 54916 12096 54972
rect 12032 54912 12096 54916
rect 12112 54972 12176 54976
rect 12112 54916 12116 54972
rect 12116 54916 12172 54972
rect 12172 54916 12176 54972
rect 12112 54912 12176 54916
rect 12192 54972 12256 54976
rect 12192 54916 12196 54972
rect 12196 54916 12252 54972
rect 12252 54916 12256 54972
rect 12192 54912 12256 54916
rect 16952 54972 17016 54976
rect 16952 54916 16956 54972
rect 16956 54916 17012 54972
rect 17012 54916 17016 54972
rect 16952 54912 17016 54916
rect 17032 54972 17096 54976
rect 17032 54916 17036 54972
rect 17036 54916 17092 54972
rect 17092 54916 17096 54972
rect 17032 54912 17096 54916
rect 17112 54972 17176 54976
rect 17112 54916 17116 54972
rect 17116 54916 17172 54972
rect 17172 54916 17176 54972
rect 17112 54912 17176 54916
rect 17192 54972 17256 54976
rect 17192 54916 17196 54972
rect 17196 54916 17252 54972
rect 17252 54916 17256 54972
rect 17192 54912 17256 54916
rect 21952 54972 22016 54976
rect 21952 54916 21956 54972
rect 21956 54916 22012 54972
rect 22012 54916 22016 54972
rect 21952 54912 22016 54916
rect 22032 54972 22096 54976
rect 22032 54916 22036 54972
rect 22036 54916 22092 54972
rect 22092 54916 22096 54972
rect 22032 54912 22096 54916
rect 22112 54972 22176 54976
rect 22112 54916 22116 54972
rect 22116 54916 22172 54972
rect 22172 54916 22176 54972
rect 22112 54912 22176 54916
rect 22192 54972 22256 54976
rect 22192 54916 22196 54972
rect 22196 54916 22252 54972
rect 22252 54916 22256 54972
rect 22192 54912 22256 54916
rect 26952 54972 27016 54976
rect 26952 54916 26956 54972
rect 26956 54916 27012 54972
rect 27012 54916 27016 54972
rect 26952 54912 27016 54916
rect 27032 54972 27096 54976
rect 27032 54916 27036 54972
rect 27036 54916 27092 54972
rect 27092 54916 27096 54972
rect 27032 54912 27096 54916
rect 27112 54972 27176 54976
rect 27112 54916 27116 54972
rect 27116 54916 27172 54972
rect 27172 54916 27176 54972
rect 27112 54912 27176 54916
rect 27192 54972 27256 54976
rect 27192 54916 27196 54972
rect 27196 54916 27252 54972
rect 27252 54916 27256 54972
rect 27192 54912 27256 54916
rect 31952 54972 32016 54976
rect 31952 54916 31956 54972
rect 31956 54916 32012 54972
rect 32012 54916 32016 54972
rect 31952 54912 32016 54916
rect 32032 54972 32096 54976
rect 32032 54916 32036 54972
rect 32036 54916 32092 54972
rect 32092 54916 32096 54972
rect 32032 54912 32096 54916
rect 32112 54972 32176 54976
rect 32112 54916 32116 54972
rect 32116 54916 32172 54972
rect 32172 54916 32176 54972
rect 32112 54912 32176 54916
rect 32192 54972 32256 54976
rect 32192 54916 32196 54972
rect 32196 54916 32252 54972
rect 32252 54916 32256 54972
rect 32192 54912 32256 54916
rect 36952 54972 37016 54976
rect 36952 54916 36956 54972
rect 36956 54916 37012 54972
rect 37012 54916 37016 54972
rect 36952 54912 37016 54916
rect 37032 54972 37096 54976
rect 37032 54916 37036 54972
rect 37036 54916 37092 54972
rect 37092 54916 37096 54972
rect 37032 54912 37096 54916
rect 37112 54972 37176 54976
rect 37112 54916 37116 54972
rect 37116 54916 37172 54972
rect 37172 54916 37176 54972
rect 37112 54912 37176 54916
rect 37192 54972 37256 54976
rect 37192 54916 37196 54972
rect 37196 54916 37252 54972
rect 37252 54916 37256 54972
rect 37192 54912 37256 54916
rect 2612 54428 2676 54432
rect 2612 54372 2616 54428
rect 2616 54372 2672 54428
rect 2672 54372 2676 54428
rect 2612 54368 2676 54372
rect 2692 54428 2756 54432
rect 2692 54372 2696 54428
rect 2696 54372 2752 54428
rect 2752 54372 2756 54428
rect 2692 54368 2756 54372
rect 2772 54428 2836 54432
rect 2772 54372 2776 54428
rect 2776 54372 2832 54428
rect 2832 54372 2836 54428
rect 2772 54368 2836 54372
rect 2852 54428 2916 54432
rect 2852 54372 2856 54428
rect 2856 54372 2912 54428
rect 2912 54372 2916 54428
rect 2852 54368 2916 54372
rect 7612 54428 7676 54432
rect 7612 54372 7616 54428
rect 7616 54372 7672 54428
rect 7672 54372 7676 54428
rect 7612 54368 7676 54372
rect 7692 54428 7756 54432
rect 7692 54372 7696 54428
rect 7696 54372 7752 54428
rect 7752 54372 7756 54428
rect 7692 54368 7756 54372
rect 7772 54428 7836 54432
rect 7772 54372 7776 54428
rect 7776 54372 7832 54428
rect 7832 54372 7836 54428
rect 7772 54368 7836 54372
rect 7852 54428 7916 54432
rect 7852 54372 7856 54428
rect 7856 54372 7912 54428
rect 7912 54372 7916 54428
rect 7852 54368 7916 54372
rect 12612 54428 12676 54432
rect 12612 54372 12616 54428
rect 12616 54372 12672 54428
rect 12672 54372 12676 54428
rect 12612 54368 12676 54372
rect 12692 54428 12756 54432
rect 12692 54372 12696 54428
rect 12696 54372 12752 54428
rect 12752 54372 12756 54428
rect 12692 54368 12756 54372
rect 12772 54428 12836 54432
rect 12772 54372 12776 54428
rect 12776 54372 12832 54428
rect 12832 54372 12836 54428
rect 12772 54368 12836 54372
rect 12852 54428 12916 54432
rect 12852 54372 12856 54428
rect 12856 54372 12912 54428
rect 12912 54372 12916 54428
rect 12852 54368 12916 54372
rect 17612 54428 17676 54432
rect 17612 54372 17616 54428
rect 17616 54372 17672 54428
rect 17672 54372 17676 54428
rect 17612 54368 17676 54372
rect 17692 54428 17756 54432
rect 17692 54372 17696 54428
rect 17696 54372 17752 54428
rect 17752 54372 17756 54428
rect 17692 54368 17756 54372
rect 17772 54428 17836 54432
rect 17772 54372 17776 54428
rect 17776 54372 17832 54428
rect 17832 54372 17836 54428
rect 17772 54368 17836 54372
rect 17852 54428 17916 54432
rect 17852 54372 17856 54428
rect 17856 54372 17912 54428
rect 17912 54372 17916 54428
rect 17852 54368 17916 54372
rect 22612 54428 22676 54432
rect 22612 54372 22616 54428
rect 22616 54372 22672 54428
rect 22672 54372 22676 54428
rect 22612 54368 22676 54372
rect 22692 54428 22756 54432
rect 22692 54372 22696 54428
rect 22696 54372 22752 54428
rect 22752 54372 22756 54428
rect 22692 54368 22756 54372
rect 22772 54428 22836 54432
rect 22772 54372 22776 54428
rect 22776 54372 22832 54428
rect 22832 54372 22836 54428
rect 22772 54368 22836 54372
rect 22852 54428 22916 54432
rect 22852 54372 22856 54428
rect 22856 54372 22912 54428
rect 22912 54372 22916 54428
rect 22852 54368 22916 54372
rect 27612 54428 27676 54432
rect 27612 54372 27616 54428
rect 27616 54372 27672 54428
rect 27672 54372 27676 54428
rect 27612 54368 27676 54372
rect 27692 54428 27756 54432
rect 27692 54372 27696 54428
rect 27696 54372 27752 54428
rect 27752 54372 27756 54428
rect 27692 54368 27756 54372
rect 27772 54428 27836 54432
rect 27772 54372 27776 54428
rect 27776 54372 27832 54428
rect 27832 54372 27836 54428
rect 27772 54368 27836 54372
rect 27852 54428 27916 54432
rect 27852 54372 27856 54428
rect 27856 54372 27912 54428
rect 27912 54372 27916 54428
rect 27852 54368 27916 54372
rect 32612 54428 32676 54432
rect 32612 54372 32616 54428
rect 32616 54372 32672 54428
rect 32672 54372 32676 54428
rect 32612 54368 32676 54372
rect 32692 54428 32756 54432
rect 32692 54372 32696 54428
rect 32696 54372 32752 54428
rect 32752 54372 32756 54428
rect 32692 54368 32756 54372
rect 32772 54428 32836 54432
rect 32772 54372 32776 54428
rect 32776 54372 32832 54428
rect 32832 54372 32836 54428
rect 32772 54368 32836 54372
rect 32852 54428 32916 54432
rect 32852 54372 32856 54428
rect 32856 54372 32912 54428
rect 32912 54372 32916 54428
rect 32852 54368 32916 54372
rect 37612 54428 37676 54432
rect 37612 54372 37616 54428
rect 37616 54372 37672 54428
rect 37672 54372 37676 54428
rect 37612 54368 37676 54372
rect 37692 54428 37756 54432
rect 37692 54372 37696 54428
rect 37696 54372 37752 54428
rect 37752 54372 37756 54428
rect 37692 54368 37756 54372
rect 37772 54428 37836 54432
rect 37772 54372 37776 54428
rect 37776 54372 37832 54428
rect 37832 54372 37836 54428
rect 37772 54368 37836 54372
rect 37852 54428 37916 54432
rect 37852 54372 37856 54428
rect 37856 54372 37912 54428
rect 37912 54372 37916 54428
rect 37852 54368 37916 54372
rect 1952 53884 2016 53888
rect 1952 53828 1956 53884
rect 1956 53828 2012 53884
rect 2012 53828 2016 53884
rect 1952 53824 2016 53828
rect 2032 53884 2096 53888
rect 2032 53828 2036 53884
rect 2036 53828 2092 53884
rect 2092 53828 2096 53884
rect 2032 53824 2096 53828
rect 2112 53884 2176 53888
rect 2112 53828 2116 53884
rect 2116 53828 2172 53884
rect 2172 53828 2176 53884
rect 2112 53824 2176 53828
rect 2192 53884 2256 53888
rect 2192 53828 2196 53884
rect 2196 53828 2252 53884
rect 2252 53828 2256 53884
rect 2192 53824 2256 53828
rect 6952 53884 7016 53888
rect 6952 53828 6956 53884
rect 6956 53828 7012 53884
rect 7012 53828 7016 53884
rect 6952 53824 7016 53828
rect 7032 53884 7096 53888
rect 7032 53828 7036 53884
rect 7036 53828 7092 53884
rect 7092 53828 7096 53884
rect 7032 53824 7096 53828
rect 7112 53884 7176 53888
rect 7112 53828 7116 53884
rect 7116 53828 7172 53884
rect 7172 53828 7176 53884
rect 7112 53824 7176 53828
rect 7192 53884 7256 53888
rect 7192 53828 7196 53884
rect 7196 53828 7252 53884
rect 7252 53828 7256 53884
rect 7192 53824 7256 53828
rect 11952 53884 12016 53888
rect 11952 53828 11956 53884
rect 11956 53828 12012 53884
rect 12012 53828 12016 53884
rect 11952 53824 12016 53828
rect 12032 53884 12096 53888
rect 12032 53828 12036 53884
rect 12036 53828 12092 53884
rect 12092 53828 12096 53884
rect 12032 53824 12096 53828
rect 12112 53884 12176 53888
rect 12112 53828 12116 53884
rect 12116 53828 12172 53884
rect 12172 53828 12176 53884
rect 12112 53824 12176 53828
rect 12192 53884 12256 53888
rect 12192 53828 12196 53884
rect 12196 53828 12252 53884
rect 12252 53828 12256 53884
rect 12192 53824 12256 53828
rect 16952 53884 17016 53888
rect 16952 53828 16956 53884
rect 16956 53828 17012 53884
rect 17012 53828 17016 53884
rect 16952 53824 17016 53828
rect 17032 53884 17096 53888
rect 17032 53828 17036 53884
rect 17036 53828 17092 53884
rect 17092 53828 17096 53884
rect 17032 53824 17096 53828
rect 17112 53884 17176 53888
rect 17112 53828 17116 53884
rect 17116 53828 17172 53884
rect 17172 53828 17176 53884
rect 17112 53824 17176 53828
rect 17192 53884 17256 53888
rect 17192 53828 17196 53884
rect 17196 53828 17252 53884
rect 17252 53828 17256 53884
rect 17192 53824 17256 53828
rect 21952 53884 22016 53888
rect 21952 53828 21956 53884
rect 21956 53828 22012 53884
rect 22012 53828 22016 53884
rect 21952 53824 22016 53828
rect 22032 53884 22096 53888
rect 22032 53828 22036 53884
rect 22036 53828 22092 53884
rect 22092 53828 22096 53884
rect 22032 53824 22096 53828
rect 22112 53884 22176 53888
rect 22112 53828 22116 53884
rect 22116 53828 22172 53884
rect 22172 53828 22176 53884
rect 22112 53824 22176 53828
rect 22192 53884 22256 53888
rect 22192 53828 22196 53884
rect 22196 53828 22252 53884
rect 22252 53828 22256 53884
rect 22192 53824 22256 53828
rect 26952 53884 27016 53888
rect 26952 53828 26956 53884
rect 26956 53828 27012 53884
rect 27012 53828 27016 53884
rect 26952 53824 27016 53828
rect 27032 53884 27096 53888
rect 27032 53828 27036 53884
rect 27036 53828 27092 53884
rect 27092 53828 27096 53884
rect 27032 53824 27096 53828
rect 27112 53884 27176 53888
rect 27112 53828 27116 53884
rect 27116 53828 27172 53884
rect 27172 53828 27176 53884
rect 27112 53824 27176 53828
rect 27192 53884 27256 53888
rect 27192 53828 27196 53884
rect 27196 53828 27252 53884
rect 27252 53828 27256 53884
rect 27192 53824 27256 53828
rect 31952 53884 32016 53888
rect 31952 53828 31956 53884
rect 31956 53828 32012 53884
rect 32012 53828 32016 53884
rect 31952 53824 32016 53828
rect 32032 53884 32096 53888
rect 32032 53828 32036 53884
rect 32036 53828 32092 53884
rect 32092 53828 32096 53884
rect 32032 53824 32096 53828
rect 32112 53884 32176 53888
rect 32112 53828 32116 53884
rect 32116 53828 32172 53884
rect 32172 53828 32176 53884
rect 32112 53824 32176 53828
rect 32192 53884 32256 53888
rect 32192 53828 32196 53884
rect 32196 53828 32252 53884
rect 32252 53828 32256 53884
rect 32192 53824 32256 53828
rect 36952 53884 37016 53888
rect 36952 53828 36956 53884
rect 36956 53828 37012 53884
rect 37012 53828 37016 53884
rect 36952 53824 37016 53828
rect 37032 53884 37096 53888
rect 37032 53828 37036 53884
rect 37036 53828 37092 53884
rect 37092 53828 37096 53884
rect 37032 53824 37096 53828
rect 37112 53884 37176 53888
rect 37112 53828 37116 53884
rect 37116 53828 37172 53884
rect 37172 53828 37176 53884
rect 37112 53824 37176 53828
rect 37192 53884 37256 53888
rect 37192 53828 37196 53884
rect 37196 53828 37252 53884
rect 37252 53828 37256 53884
rect 37192 53824 37256 53828
rect 2612 53340 2676 53344
rect 2612 53284 2616 53340
rect 2616 53284 2672 53340
rect 2672 53284 2676 53340
rect 2612 53280 2676 53284
rect 2692 53340 2756 53344
rect 2692 53284 2696 53340
rect 2696 53284 2752 53340
rect 2752 53284 2756 53340
rect 2692 53280 2756 53284
rect 2772 53340 2836 53344
rect 2772 53284 2776 53340
rect 2776 53284 2832 53340
rect 2832 53284 2836 53340
rect 2772 53280 2836 53284
rect 2852 53340 2916 53344
rect 2852 53284 2856 53340
rect 2856 53284 2912 53340
rect 2912 53284 2916 53340
rect 2852 53280 2916 53284
rect 7612 53340 7676 53344
rect 7612 53284 7616 53340
rect 7616 53284 7672 53340
rect 7672 53284 7676 53340
rect 7612 53280 7676 53284
rect 7692 53340 7756 53344
rect 7692 53284 7696 53340
rect 7696 53284 7752 53340
rect 7752 53284 7756 53340
rect 7692 53280 7756 53284
rect 7772 53340 7836 53344
rect 7772 53284 7776 53340
rect 7776 53284 7832 53340
rect 7832 53284 7836 53340
rect 7772 53280 7836 53284
rect 7852 53340 7916 53344
rect 7852 53284 7856 53340
rect 7856 53284 7912 53340
rect 7912 53284 7916 53340
rect 7852 53280 7916 53284
rect 12612 53340 12676 53344
rect 12612 53284 12616 53340
rect 12616 53284 12672 53340
rect 12672 53284 12676 53340
rect 12612 53280 12676 53284
rect 12692 53340 12756 53344
rect 12692 53284 12696 53340
rect 12696 53284 12752 53340
rect 12752 53284 12756 53340
rect 12692 53280 12756 53284
rect 12772 53340 12836 53344
rect 12772 53284 12776 53340
rect 12776 53284 12832 53340
rect 12832 53284 12836 53340
rect 12772 53280 12836 53284
rect 12852 53340 12916 53344
rect 12852 53284 12856 53340
rect 12856 53284 12912 53340
rect 12912 53284 12916 53340
rect 12852 53280 12916 53284
rect 17612 53340 17676 53344
rect 17612 53284 17616 53340
rect 17616 53284 17672 53340
rect 17672 53284 17676 53340
rect 17612 53280 17676 53284
rect 17692 53340 17756 53344
rect 17692 53284 17696 53340
rect 17696 53284 17752 53340
rect 17752 53284 17756 53340
rect 17692 53280 17756 53284
rect 17772 53340 17836 53344
rect 17772 53284 17776 53340
rect 17776 53284 17832 53340
rect 17832 53284 17836 53340
rect 17772 53280 17836 53284
rect 17852 53340 17916 53344
rect 17852 53284 17856 53340
rect 17856 53284 17912 53340
rect 17912 53284 17916 53340
rect 17852 53280 17916 53284
rect 22612 53340 22676 53344
rect 22612 53284 22616 53340
rect 22616 53284 22672 53340
rect 22672 53284 22676 53340
rect 22612 53280 22676 53284
rect 22692 53340 22756 53344
rect 22692 53284 22696 53340
rect 22696 53284 22752 53340
rect 22752 53284 22756 53340
rect 22692 53280 22756 53284
rect 22772 53340 22836 53344
rect 22772 53284 22776 53340
rect 22776 53284 22832 53340
rect 22832 53284 22836 53340
rect 22772 53280 22836 53284
rect 22852 53340 22916 53344
rect 22852 53284 22856 53340
rect 22856 53284 22912 53340
rect 22912 53284 22916 53340
rect 22852 53280 22916 53284
rect 27612 53340 27676 53344
rect 27612 53284 27616 53340
rect 27616 53284 27672 53340
rect 27672 53284 27676 53340
rect 27612 53280 27676 53284
rect 27692 53340 27756 53344
rect 27692 53284 27696 53340
rect 27696 53284 27752 53340
rect 27752 53284 27756 53340
rect 27692 53280 27756 53284
rect 27772 53340 27836 53344
rect 27772 53284 27776 53340
rect 27776 53284 27832 53340
rect 27832 53284 27836 53340
rect 27772 53280 27836 53284
rect 27852 53340 27916 53344
rect 27852 53284 27856 53340
rect 27856 53284 27912 53340
rect 27912 53284 27916 53340
rect 27852 53280 27916 53284
rect 32612 53340 32676 53344
rect 32612 53284 32616 53340
rect 32616 53284 32672 53340
rect 32672 53284 32676 53340
rect 32612 53280 32676 53284
rect 32692 53340 32756 53344
rect 32692 53284 32696 53340
rect 32696 53284 32752 53340
rect 32752 53284 32756 53340
rect 32692 53280 32756 53284
rect 32772 53340 32836 53344
rect 32772 53284 32776 53340
rect 32776 53284 32832 53340
rect 32832 53284 32836 53340
rect 32772 53280 32836 53284
rect 32852 53340 32916 53344
rect 32852 53284 32856 53340
rect 32856 53284 32912 53340
rect 32912 53284 32916 53340
rect 32852 53280 32916 53284
rect 37612 53340 37676 53344
rect 37612 53284 37616 53340
rect 37616 53284 37672 53340
rect 37672 53284 37676 53340
rect 37612 53280 37676 53284
rect 37692 53340 37756 53344
rect 37692 53284 37696 53340
rect 37696 53284 37752 53340
rect 37752 53284 37756 53340
rect 37692 53280 37756 53284
rect 37772 53340 37836 53344
rect 37772 53284 37776 53340
rect 37776 53284 37832 53340
rect 37832 53284 37836 53340
rect 37772 53280 37836 53284
rect 37852 53340 37916 53344
rect 37852 53284 37856 53340
rect 37856 53284 37912 53340
rect 37912 53284 37916 53340
rect 37852 53280 37916 53284
rect 1952 52796 2016 52800
rect 1952 52740 1956 52796
rect 1956 52740 2012 52796
rect 2012 52740 2016 52796
rect 1952 52736 2016 52740
rect 2032 52796 2096 52800
rect 2032 52740 2036 52796
rect 2036 52740 2092 52796
rect 2092 52740 2096 52796
rect 2032 52736 2096 52740
rect 2112 52796 2176 52800
rect 2112 52740 2116 52796
rect 2116 52740 2172 52796
rect 2172 52740 2176 52796
rect 2112 52736 2176 52740
rect 2192 52796 2256 52800
rect 2192 52740 2196 52796
rect 2196 52740 2252 52796
rect 2252 52740 2256 52796
rect 2192 52736 2256 52740
rect 6952 52796 7016 52800
rect 6952 52740 6956 52796
rect 6956 52740 7012 52796
rect 7012 52740 7016 52796
rect 6952 52736 7016 52740
rect 7032 52796 7096 52800
rect 7032 52740 7036 52796
rect 7036 52740 7092 52796
rect 7092 52740 7096 52796
rect 7032 52736 7096 52740
rect 7112 52796 7176 52800
rect 7112 52740 7116 52796
rect 7116 52740 7172 52796
rect 7172 52740 7176 52796
rect 7112 52736 7176 52740
rect 7192 52796 7256 52800
rect 7192 52740 7196 52796
rect 7196 52740 7252 52796
rect 7252 52740 7256 52796
rect 7192 52736 7256 52740
rect 11952 52796 12016 52800
rect 11952 52740 11956 52796
rect 11956 52740 12012 52796
rect 12012 52740 12016 52796
rect 11952 52736 12016 52740
rect 12032 52796 12096 52800
rect 12032 52740 12036 52796
rect 12036 52740 12092 52796
rect 12092 52740 12096 52796
rect 12032 52736 12096 52740
rect 12112 52796 12176 52800
rect 12112 52740 12116 52796
rect 12116 52740 12172 52796
rect 12172 52740 12176 52796
rect 12112 52736 12176 52740
rect 12192 52796 12256 52800
rect 12192 52740 12196 52796
rect 12196 52740 12252 52796
rect 12252 52740 12256 52796
rect 12192 52736 12256 52740
rect 16952 52796 17016 52800
rect 16952 52740 16956 52796
rect 16956 52740 17012 52796
rect 17012 52740 17016 52796
rect 16952 52736 17016 52740
rect 17032 52796 17096 52800
rect 17032 52740 17036 52796
rect 17036 52740 17092 52796
rect 17092 52740 17096 52796
rect 17032 52736 17096 52740
rect 17112 52796 17176 52800
rect 17112 52740 17116 52796
rect 17116 52740 17172 52796
rect 17172 52740 17176 52796
rect 17112 52736 17176 52740
rect 17192 52796 17256 52800
rect 17192 52740 17196 52796
rect 17196 52740 17252 52796
rect 17252 52740 17256 52796
rect 17192 52736 17256 52740
rect 21952 52796 22016 52800
rect 21952 52740 21956 52796
rect 21956 52740 22012 52796
rect 22012 52740 22016 52796
rect 21952 52736 22016 52740
rect 22032 52796 22096 52800
rect 22032 52740 22036 52796
rect 22036 52740 22092 52796
rect 22092 52740 22096 52796
rect 22032 52736 22096 52740
rect 22112 52796 22176 52800
rect 22112 52740 22116 52796
rect 22116 52740 22172 52796
rect 22172 52740 22176 52796
rect 22112 52736 22176 52740
rect 22192 52796 22256 52800
rect 22192 52740 22196 52796
rect 22196 52740 22252 52796
rect 22252 52740 22256 52796
rect 22192 52736 22256 52740
rect 26952 52796 27016 52800
rect 26952 52740 26956 52796
rect 26956 52740 27012 52796
rect 27012 52740 27016 52796
rect 26952 52736 27016 52740
rect 27032 52796 27096 52800
rect 27032 52740 27036 52796
rect 27036 52740 27092 52796
rect 27092 52740 27096 52796
rect 27032 52736 27096 52740
rect 27112 52796 27176 52800
rect 27112 52740 27116 52796
rect 27116 52740 27172 52796
rect 27172 52740 27176 52796
rect 27112 52736 27176 52740
rect 27192 52796 27256 52800
rect 27192 52740 27196 52796
rect 27196 52740 27252 52796
rect 27252 52740 27256 52796
rect 27192 52736 27256 52740
rect 31952 52796 32016 52800
rect 31952 52740 31956 52796
rect 31956 52740 32012 52796
rect 32012 52740 32016 52796
rect 31952 52736 32016 52740
rect 32032 52796 32096 52800
rect 32032 52740 32036 52796
rect 32036 52740 32092 52796
rect 32092 52740 32096 52796
rect 32032 52736 32096 52740
rect 32112 52796 32176 52800
rect 32112 52740 32116 52796
rect 32116 52740 32172 52796
rect 32172 52740 32176 52796
rect 32112 52736 32176 52740
rect 32192 52796 32256 52800
rect 32192 52740 32196 52796
rect 32196 52740 32252 52796
rect 32252 52740 32256 52796
rect 32192 52736 32256 52740
rect 36952 52796 37016 52800
rect 36952 52740 36956 52796
rect 36956 52740 37012 52796
rect 37012 52740 37016 52796
rect 36952 52736 37016 52740
rect 37032 52796 37096 52800
rect 37032 52740 37036 52796
rect 37036 52740 37092 52796
rect 37092 52740 37096 52796
rect 37032 52736 37096 52740
rect 37112 52796 37176 52800
rect 37112 52740 37116 52796
rect 37116 52740 37172 52796
rect 37172 52740 37176 52796
rect 37112 52736 37176 52740
rect 37192 52796 37256 52800
rect 37192 52740 37196 52796
rect 37196 52740 37252 52796
rect 37252 52740 37256 52796
rect 37192 52736 37256 52740
rect 2612 52252 2676 52256
rect 2612 52196 2616 52252
rect 2616 52196 2672 52252
rect 2672 52196 2676 52252
rect 2612 52192 2676 52196
rect 2692 52252 2756 52256
rect 2692 52196 2696 52252
rect 2696 52196 2752 52252
rect 2752 52196 2756 52252
rect 2692 52192 2756 52196
rect 2772 52252 2836 52256
rect 2772 52196 2776 52252
rect 2776 52196 2832 52252
rect 2832 52196 2836 52252
rect 2772 52192 2836 52196
rect 2852 52252 2916 52256
rect 2852 52196 2856 52252
rect 2856 52196 2912 52252
rect 2912 52196 2916 52252
rect 2852 52192 2916 52196
rect 7612 52252 7676 52256
rect 7612 52196 7616 52252
rect 7616 52196 7672 52252
rect 7672 52196 7676 52252
rect 7612 52192 7676 52196
rect 7692 52252 7756 52256
rect 7692 52196 7696 52252
rect 7696 52196 7752 52252
rect 7752 52196 7756 52252
rect 7692 52192 7756 52196
rect 7772 52252 7836 52256
rect 7772 52196 7776 52252
rect 7776 52196 7832 52252
rect 7832 52196 7836 52252
rect 7772 52192 7836 52196
rect 7852 52252 7916 52256
rect 7852 52196 7856 52252
rect 7856 52196 7912 52252
rect 7912 52196 7916 52252
rect 7852 52192 7916 52196
rect 12612 52252 12676 52256
rect 12612 52196 12616 52252
rect 12616 52196 12672 52252
rect 12672 52196 12676 52252
rect 12612 52192 12676 52196
rect 12692 52252 12756 52256
rect 12692 52196 12696 52252
rect 12696 52196 12752 52252
rect 12752 52196 12756 52252
rect 12692 52192 12756 52196
rect 12772 52252 12836 52256
rect 12772 52196 12776 52252
rect 12776 52196 12832 52252
rect 12832 52196 12836 52252
rect 12772 52192 12836 52196
rect 12852 52252 12916 52256
rect 12852 52196 12856 52252
rect 12856 52196 12912 52252
rect 12912 52196 12916 52252
rect 12852 52192 12916 52196
rect 17612 52252 17676 52256
rect 17612 52196 17616 52252
rect 17616 52196 17672 52252
rect 17672 52196 17676 52252
rect 17612 52192 17676 52196
rect 17692 52252 17756 52256
rect 17692 52196 17696 52252
rect 17696 52196 17752 52252
rect 17752 52196 17756 52252
rect 17692 52192 17756 52196
rect 17772 52252 17836 52256
rect 17772 52196 17776 52252
rect 17776 52196 17832 52252
rect 17832 52196 17836 52252
rect 17772 52192 17836 52196
rect 17852 52252 17916 52256
rect 17852 52196 17856 52252
rect 17856 52196 17912 52252
rect 17912 52196 17916 52252
rect 17852 52192 17916 52196
rect 22612 52252 22676 52256
rect 22612 52196 22616 52252
rect 22616 52196 22672 52252
rect 22672 52196 22676 52252
rect 22612 52192 22676 52196
rect 22692 52252 22756 52256
rect 22692 52196 22696 52252
rect 22696 52196 22752 52252
rect 22752 52196 22756 52252
rect 22692 52192 22756 52196
rect 22772 52252 22836 52256
rect 22772 52196 22776 52252
rect 22776 52196 22832 52252
rect 22832 52196 22836 52252
rect 22772 52192 22836 52196
rect 22852 52252 22916 52256
rect 22852 52196 22856 52252
rect 22856 52196 22912 52252
rect 22912 52196 22916 52252
rect 22852 52192 22916 52196
rect 27612 52252 27676 52256
rect 27612 52196 27616 52252
rect 27616 52196 27672 52252
rect 27672 52196 27676 52252
rect 27612 52192 27676 52196
rect 27692 52252 27756 52256
rect 27692 52196 27696 52252
rect 27696 52196 27752 52252
rect 27752 52196 27756 52252
rect 27692 52192 27756 52196
rect 27772 52252 27836 52256
rect 27772 52196 27776 52252
rect 27776 52196 27832 52252
rect 27832 52196 27836 52252
rect 27772 52192 27836 52196
rect 27852 52252 27916 52256
rect 27852 52196 27856 52252
rect 27856 52196 27912 52252
rect 27912 52196 27916 52252
rect 27852 52192 27916 52196
rect 32612 52252 32676 52256
rect 32612 52196 32616 52252
rect 32616 52196 32672 52252
rect 32672 52196 32676 52252
rect 32612 52192 32676 52196
rect 32692 52252 32756 52256
rect 32692 52196 32696 52252
rect 32696 52196 32752 52252
rect 32752 52196 32756 52252
rect 32692 52192 32756 52196
rect 32772 52252 32836 52256
rect 32772 52196 32776 52252
rect 32776 52196 32832 52252
rect 32832 52196 32836 52252
rect 32772 52192 32836 52196
rect 32852 52252 32916 52256
rect 32852 52196 32856 52252
rect 32856 52196 32912 52252
rect 32912 52196 32916 52252
rect 32852 52192 32916 52196
rect 37612 52252 37676 52256
rect 37612 52196 37616 52252
rect 37616 52196 37672 52252
rect 37672 52196 37676 52252
rect 37612 52192 37676 52196
rect 37692 52252 37756 52256
rect 37692 52196 37696 52252
rect 37696 52196 37752 52252
rect 37752 52196 37756 52252
rect 37692 52192 37756 52196
rect 37772 52252 37836 52256
rect 37772 52196 37776 52252
rect 37776 52196 37832 52252
rect 37832 52196 37836 52252
rect 37772 52192 37836 52196
rect 37852 52252 37916 52256
rect 37852 52196 37856 52252
rect 37856 52196 37912 52252
rect 37912 52196 37916 52252
rect 37852 52192 37916 52196
rect 1952 51708 2016 51712
rect 1952 51652 1956 51708
rect 1956 51652 2012 51708
rect 2012 51652 2016 51708
rect 1952 51648 2016 51652
rect 2032 51708 2096 51712
rect 2032 51652 2036 51708
rect 2036 51652 2092 51708
rect 2092 51652 2096 51708
rect 2032 51648 2096 51652
rect 2112 51708 2176 51712
rect 2112 51652 2116 51708
rect 2116 51652 2172 51708
rect 2172 51652 2176 51708
rect 2112 51648 2176 51652
rect 2192 51708 2256 51712
rect 2192 51652 2196 51708
rect 2196 51652 2252 51708
rect 2252 51652 2256 51708
rect 2192 51648 2256 51652
rect 6952 51708 7016 51712
rect 6952 51652 6956 51708
rect 6956 51652 7012 51708
rect 7012 51652 7016 51708
rect 6952 51648 7016 51652
rect 7032 51708 7096 51712
rect 7032 51652 7036 51708
rect 7036 51652 7092 51708
rect 7092 51652 7096 51708
rect 7032 51648 7096 51652
rect 7112 51708 7176 51712
rect 7112 51652 7116 51708
rect 7116 51652 7172 51708
rect 7172 51652 7176 51708
rect 7112 51648 7176 51652
rect 7192 51708 7256 51712
rect 7192 51652 7196 51708
rect 7196 51652 7252 51708
rect 7252 51652 7256 51708
rect 7192 51648 7256 51652
rect 11952 51708 12016 51712
rect 11952 51652 11956 51708
rect 11956 51652 12012 51708
rect 12012 51652 12016 51708
rect 11952 51648 12016 51652
rect 12032 51708 12096 51712
rect 12032 51652 12036 51708
rect 12036 51652 12092 51708
rect 12092 51652 12096 51708
rect 12032 51648 12096 51652
rect 12112 51708 12176 51712
rect 12112 51652 12116 51708
rect 12116 51652 12172 51708
rect 12172 51652 12176 51708
rect 12112 51648 12176 51652
rect 12192 51708 12256 51712
rect 12192 51652 12196 51708
rect 12196 51652 12252 51708
rect 12252 51652 12256 51708
rect 12192 51648 12256 51652
rect 16952 51708 17016 51712
rect 16952 51652 16956 51708
rect 16956 51652 17012 51708
rect 17012 51652 17016 51708
rect 16952 51648 17016 51652
rect 17032 51708 17096 51712
rect 17032 51652 17036 51708
rect 17036 51652 17092 51708
rect 17092 51652 17096 51708
rect 17032 51648 17096 51652
rect 17112 51708 17176 51712
rect 17112 51652 17116 51708
rect 17116 51652 17172 51708
rect 17172 51652 17176 51708
rect 17112 51648 17176 51652
rect 17192 51708 17256 51712
rect 17192 51652 17196 51708
rect 17196 51652 17252 51708
rect 17252 51652 17256 51708
rect 17192 51648 17256 51652
rect 21952 51708 22016 51712
rect 21952 51652 21956 51708
rect 21956 51652 22012 51708
rect 22012 51652 22016 51708
rect 21952 51648 22016 51652
rect 22032 51708 22096 51712
rect 22032 51652 22036 51708
rect 22036 51652 22092 51708
rect 22092 51652 22096 51708
rect 22032 51648 22096 51652
rect 22112 51708 22176 51712
rect 22112 51652 22116 51708
rect 22116 51652 22172 51708
rect 22172 51652 22176 51708
rect 22112 51648 22176 51652
rect 22192 51708 22256 51712
rect 22192 51652 22196 51708
rect 22196 51652 22252 51708
rect 22252 51652 22256 51708
rect 22192 51648 22256 51652
rect 26952 51708 27016 51712
rect 26952 51652 26956 51708
rect 26956 51652 27012 51708
rect 27012 51652 27016 51708
rect 26952 51648 27016 51652
rect 27032 51708 27096 51712
rect 27032 51652 27036 51708
rect 27036 51652 27092 51708
rect 27092 51652 27096 51708
rect 27032 51648 27096 51652
rect 27112 51708 27176 51712
rect 27112 51652 27116 51708
rect 27116 51652 27172 51708
rect 27172 51652 27176 51708
rect 27112 51648 27176 51652
rect 27192 51708 27256 51712
rect 27192 51652 27196 51708
rect 27196 51652 27252 51708
rect 27252 51652 27256 51708
rect 27192 51648 27256 51652
rect 31952 51708 32016 51712
rect 31952 51652 31956 51708
rect 31956 51652 32012 51708
rect 32012 51652 32016 51708
rect 31952 51648 32016 51652
rect 32032 51708 32096 51712
rect 32032 51652 32036 51708
rect 32036 51652 32092 51708
rect 32092 51652 32096 51708
rect 32032 51648 32096 51652
rect 32112 51708 32176 51712
rect 32112 51652 32116 51708
rect 32116 51652 32172 51708
rect 32172 51652 32176 51708
rect 32112 51648 32176 51652
rect 32192 51708 32256 51712
rect 32192 51652 32196 51708
rect 32196 51652 32252 51708
rect 32252 51652 32256 51708
rect 32192 51648 32256 51652
rect 36952 51708 37016 51712
rect 36952 51652 36956 51708
rect 36956 51652 37012 51708
rect 37012 51652 37016 51708
rect 36952 51648 37016 51652
rect 37032 51708 37096 51712
rect 37032 51652 37036 51708
rect 37036 51652 37092 51708
rect 37092 51652 37096 51708
rect 37032 51648 37096 51652
rect 37112 51708 37176 51712
rect 37112 51652 37116 51708
rect 37116 51652 37172 51708
rect 37172 51652 37176 51708
rect 37112 51648 37176 51652
rect 37192 51708 37256 51712
rect 37192 51652 37196 51708
rect 37196 51652 37252 51708
rect 37252 51652 37256 51708
rect 37192 51648 37256 51652
rect 33364 51172 33428 51236
rect 2612 51164 2676 51168
rect 2612 51108 2616 51164
rect 2616 51108 2672 51164
rect 2672 51108 2676 51164
rect 2612 51104 2676 51108
rect 2692 51164 2756 51168
rect 2692 51108 2696 51164
rect 2696 51108 2752 51164
rect 2752 51108 2756 51164
rect 2692 51104 2756 51108
rect 2772 51164 2836 51168
rect 2772 51108 2776 51164
rect 2776 51108 2832 51164
rect 2832 51108 2836 51164
rect 2772 51104 2836 51108
rect 2852 51164 2916 51168
rect 2852 51108 2856 51164
rect 2856 51108 2912 51164
rect 2912 51108 2916 51164
rect 2852 51104 2916 51108
rect 7612 51164 7676 51168
rect 7612 51108 7616 51164
rect 7616 51108 7672 51164
rect 7672 51108 7676 51164
rect 7612 51104 7676 51108
rect 7692 51164 7756 51168
rect 7692 51108 7696 51164
rect 7696 51108 7752 51164
rect 7752 51108 7756 51164
rect 7692 51104 7756 51108
rect 7772 51164 7836 51168
rect 7772 51108 7776 51164
rect 7776 51108 7832 51164
rect 7832 51108 7836 51164
rect 7772 51104 7836 51108
rect 7852 51164 7916 51168
rect 7852 51108 7856 51164
rect 7856 51108 7912 51164
rect 7912 51108 7916 51164
rect 7852 51104 7916 51108
rect 12612 51164 12676 51168
rect 12612 51108 12616 51164
rect 12616 51108 12672 51164
rect 12672 51108 12676 51164
rect 12612 51104 12676 51108
rect 12692 51164 12756 51168
rect 12692 51108 12696 51164
rect 12696 51108 12752 51164
rect 12752 51108 12756 51164
rect 12692 51104 12756 51108
rect 12772 51164 12836 51168
rect 12772 51108 12776 51164
rect 12776 51108 12832 51164
rect 12832 51108 12836 51164
rect 12772 51104 12836 51108
rect 12852 51164 12916 51168
rect 12852 51108 12856 51164
rect 12856 51108 12912 51164
rect 12912 51108 12916 51164
rect 12852 51104 12916 51108
rect 17612 51164 17676 51168
rect 17612 51108 17616 51164
rect 17616 51108 17672 51164
rect 17672 51108 17676 51164
rect 17612 51104 17676 51108
rect 17692 51164 17756 51168
rect 17692 51108 17696 51164
rect 17696 51108 17752 51164
rect 17752 51108 17756 51164
rect 17692 51104 17756 51108
rect 17772 51164 17836 51168
rect 17772 51108 17776 51164
rect 17776 51108 17832 51164
rect 17832 51108 17836 51164
rect 17772 51104 17836 51108
rect 17852 51164 17916 51168
rect 17852 51108 17856 51164
rect 17856 51108 17912 51164
rect 17912 51108 17916 51164
rect 17852 51104 17916 51108
rect 22612 51164 22676 51168
rect 22612 51108 22616 51164
rect 22616 51108 22672 51164
rect 22672 51108 22676 51164
rect 22612 51104 22676 51108
rect 22692 51164 22756 51168
rect 22692 51108 22696 51164
rect 22696 51108 22752 51164
rect 22752 51108 22756 51164
rect 22692 51104 22756 51108
rect 22772 51164 22836 51168
rect 22772 51108 22776 51164
rect 22776 51108 22832 51164
rect 22832 51108 22836 51164
rect 22772 51104 22836 51108
rect 22852 51164 22916 51168
rect 22852 51108 22856 51164
rect 22856 51108 22912 51164
rect 22912 51108 22916 51164
rect 22852 51104 22916 51108
rect 27612 51164 27676 51168
rect 27612 51108 27616 51164
rect 27616 51108 27672 51164
rect 27672 51108 27676 51164
rect 27612 51104 27676 51108
rect 27692 51164 27756 51168
rect 27692 51108 27696 51164
rect 27696 51108 27752 51164
rect 27752 51108 27756 51164
rect 27692 51104 27756 51108
rect 27772 51164 27836 51168
rect 27772 51108 27776 51164
rect 27776 51108 27832 51164
rect 27832 51108 27836 51164
rect 27772 51104 27836 51108
rect 27852 51164 27916 51168
rect 27852 51108 27856 51164
rect 27856 51108 27912 51164
rect 27912 51108 27916 51164
rect 27852 51104 27916 51108
rect 32612 51164 32676 51168
rect 32612 51108 32616 51164
rect 32616 51108 32672 51164
rect 32672 51108 32676 51164
rect 32612 51104 32676 51108
rect 32692 51164 32756 51168
rect 32692 51108 32696 51164
rect 32696 51108 32752 51164
rect 32752 51108 32756 51164
rect 32692 51104 32756 51108
rect 32772 51164 32836 51168
rect 32772 51108 32776 51164
rect 32776 51108 32832 51164
rect 32832 51108 32836 51164
rect 32772 51104 32836 51108
rect 32852 51164 32916 51168
rect 32852 51108 32856 51164
rect 32856 51108 32912 51164
rect 32912 51108 32916 51164
rect 32852 51104 32916 51108
rect 37612 51164 37676 51168
rect 37612 51108 37616 51164
rect 37616 51108 37672 51164
rect 37672 51108 37676 51164
rect 37612 51104 37676 51108
rect 37692 51164 37756 51168
rect 37692 51108 37696 51164
rect 37696 51108 37752 51164
rect 37752 51108 37756 51164
rect 37692 51104 37756 51108
rect 37772 51164 37836 51168
rect 37772 51108 37776 51164
rect 37776 51108 37832 51164
rect 37832 51108 37836 51164
rect 37772 51104 37836 51108
rect 37852 51164 37916 51168
rect 37852 51108 37856 51164
rect 37856 51108 37912 51164
rect 37912 51108 37916 51164
rect 37852 51104 37916 51108
rect 31708 50900 31772 50964
rect 32444 50900 32508 50964
rect 1952 50620 2016 50624
rect 1952 50564 1956 50620
rect 1956 50564 2012 50620
rect 2012 50564 2016 50620
rect 1952 50560 2016 50564
rect 2032 50620 2096 50624
rect 2032 50564 2036 50620
rect 2036 50564 2092 50620
rect 2092 50564 2096 50620
rect 2032 50560 2096 50564
rect 2112 50620 2176 50624
rect 2112 50564 2116 50620
rect 2116 50564 2172 50620
rect 2172 50564 2176 50620
rect 2112 50560 2176 50564
rect 2192 50620 2256 50624
rect 2192 50564 2196 50620
rect 2196 50564 2252 50620
rect 2252 50564 2256 50620
rect 2192 50560 2256 50564
rect 6952 50620 7016 50624
rect 6952 50564 6956 50620
rect 6956 50564 7012 50620
rect 7012 50564 7016 50620
rect 6952 50560 7016 50564
rect 7032 50620 7096 50624
rect 7032 50564 7036 50620
rect 7036 50564 7092 50620
rect 7092 50564 7096 50620
rect 7032 50560 7096 50564
rect 7112 50620 7176 50624
rect 7112 50564 7116 50620
rect 7116 50564 7172 50620
rect 7172 50564 7176 50620
rect 7112 50560 7176 50564
rect 7192 50620 7256 50624
rect 7192 50564 7196 50620
rect 7196 50564 7252 50620
rect 7252 50564 7256 50620
rect 7192 50560 7256 50564
rect 11952 50620 12016 50624
rect 11952 50564 11956 50620
rect 11956 50564 12012 50620
rect 12012 50564 12016 50620
rect 11952 50560 12016 50564
rect 12032 50620 12096 50624
rect 12032 50564 12036 50620
rect 12036 50564 12092 50620
rect 12092 50564 12096 50620
rect 12032 50560 12096 50564
rect 12112 50620 12176 50624
rect 12112 50564 12116 50620
rect 12116 50564 12172 50620
rect 12172 50564 12176 50620
rect 12112 50560 12176 50564
rect 12192 50620 12256 50624
rect 12192 50564 12196 50620
rect 12196 50564 12252 50620
rect 12252 50564 12256 50620
rect 12192 50560 12256 50564
rect 16952 50620 17016 50624
rect 16952 50564 16956 50620
rect 16956 50564 17012 50620
rect 17012 50564 17016 50620
rect 16952 50560 17016 50564
rect 17032 50620 17096 50624
rect 17032 50564 17036 50620
rect 17036 50564 17092 50620
rect 17092 50564 17096 50620
rect 17032 50560 17096 50564
rect 17112 50620 17176 50624
rect 17112 50564 17116 50620
rect 17116 50564 17172 50620
rect 17172 50564 17176 50620
rect 17112 50560 17176 50564
rect 17192 50620 17256 50624
rect 17192 50564 17196 50620
rect 17196 50564 17252 50620
rect 17252 50564 17256 50620
rect 17192 50560 17256 50564
rect 21952 50620 22016 50624
rect 21952 50564 21956 50620
rect 21956 50564 22012 50620
rect 22012 50564 22016 50620
rect 21952 50560 22016 50564
rect 22032 50620 22096 50624
rect 22032 50564 22036 50620
rect 22036 50564 22092 50620
rect 22092 50564 22096 50620
rect 22032 50560 22096 50564
rect 22112 50620 22176 50624
rect 22112 50564 22116 50620
rect 22116 50564 22172 50620
rect 22172 50564 22176 50620
rect 22112 50560 22176 50564
rect 22192 50620 22256 50624
rect 22192 50564 22196 50620
rect 22196 50564 22252 50620
rect 22252 50564 22256 50620
rect 22192 50560 22256 50564
rect 26952 50620 27016 50624
rect 26952 50564 26956 50620
rect 26956 50564 27012 50620
rect 27012 50564 27016 50620
rect 26952 50560 27016 50564
rect 27032 50620 27096 50624
rect 27032 50564 27036 50620
rect 27036 50564 27092 50620
rect 27092 50564 27096 50620
rect 27032 50560 27096 50564
rect 27112 50620 27176 50624
rect 27112 50564 27116 50620
rect 27116 50564 27172 50620
rect 27172 50564 27176 50620
rect 27112 50560 27176 50564
rect 27192 50620 27256 50624
rect 27192 50564 27196 50620
rect 27196 50564 27252 50620
rect 27252 50564 27256 50620
rect 27192 50560 27256 50564
rect 31952 50620 32016 50624
rect 31952 50564 31956 50620
rect 31956 50564 32012 50620
rect 32012 50564 32016 50620
rect 31952 50560 32016 50564
rect 32032 50620 32096 50624
rect 32032 50564 32036 50620
rect 32036 50564 32092 50620
rect 32092 50564 32096 50620
rect 32032 50560 32096 50564
rect 32112 50620 32176 50624
rect 32112 50564 32116 50620
rect 32116 50564 32172 50620
rect 32172 50564 32176 50620
rect 32112 50560 32176 50564
rect 32192 50620 32256 50624
rect 32192 50564 32196 50620
rect 32196 50564 32252 50620
rect 32252 50564 32256 50620
rect 32192 50560 32256 50564
rect 36952 50620 37016 50624
rect 36952 50564 36956 50620
rect 36956 50564 37012 50620
rect 37012 50564 37016 50620
rect 36952 50560 37016 50564
rect 37032 50620 37096 50624
rect 37032 50564 37036 50620
rect 37036 50564 37092 50620
rect 37092 50564 37096 50620
rect 37032 50560 37096 50564
rect 37112 50620 37176 50624
rect 37112 50564 37116 50620
rect 37116 50564 37172 50620
rect 37172 50564 37176 50620
rect 37112 50560 37176 50564
rect 37192 50620 37256 50624
rect 37192 50564 37196 50620
rect 37196 50564 37252 50620
rect 37252 50564 37256 50620
rect 37192 50560 37256 50564
rect 2612 50076 2676 50080
rect 2612 50020 2616 50076
rect 2616 50020 2672 50076
rect 2672 50020 2676 50076
rect 2612 50016 2676 50020
rect 2692 50076 2756 50080
rect 2692 50020 2696 50076
rect 2696 50020 2752 50076
rect 2752 50020 2756 50076
rect 2692 50016 2756 50020
rect 2772 50076 2836 50080
rect 2772 50020 2776 50076
rect 2776 50020 2832 50076
rect 2832 50020 2836 50076
rect 2772 50016 2836 50020
rect 2852 50076 2916 50080
rect 2852 50020 2856 50076
rect 2856 50020 2912 50076
rect 2912 50020 2916 50076
rect 2852 50016 2916 50020
rect 7612 50076 7676 50080
rect 7612 50020 7616 50076
rect 7616 50020 7672 50076
rect 7672 50020 7676 50076
rect 7612 50016 7676 50020
rect 7692 50076 7756 50080
rect 7692 50020 7696 50076
rect 7696 50020 7752 50076
rect 7752 50020 7756 50076
rect 7692 50016 7756 50020
rect 7772 50076 7836 50080
rect 7772 50020 7776 50076
rect 7776 50020 7832 50076
rect 7832 50020 7836 50076
rect 7772 50016 7836 50020
rect 7852 50076 7916 50080
rect 7852 50020 7856 50076
rect 7856 50020 7912 50076
rect 7912 50020 7916 50076
rect 7852 50016 7916 50020
rect 12612 50076 12676 50080
rect 12612 50020 12616 50076
rect 12616 50020 12672 50076
rect 12672 50020 12676 50076
rect 12612 50016 12676 50020
rect 12692 50076 12756 50080
rect 12692 50020 12696 50076
rect 12696 50020 12752 50076
rect 12752 50020 12756 50076
rect 12692 50016 12756 50020
rect 12772 50076 12836 50080
rect 12772 50020 12776 50076
rect 12776 50020 12832 50076
rect 12832 50020 12836 50076
rect 12772 50016 12836 50020
rect 12852 50076 12916 50080
rect 12852 50020 12856 50076
rect 12856 50020 12912 50076
rect 12912 50020 12916 50076
rect 12852 50016 12916 50020
rect 17612 50076 17676 50080
rect 17612 50020 17616 50076
rect 17616 50020 17672 50076
rect 17672 50020 17676 50076
rect 17612 50016 17676 50020
rect 17692 50076 17756 50080
rect 17692 50020 17696 50076
rect 17696 50020 17752 50076
rect 17752 50020 17756 50076
rect 17692 50016 17756 50020
rect 17772 50076 17836 50080
rect 17772 50020 17776 50076
rect 17776 50020 17832 50076
rect 17832 50020 17836 50076
rect 17772 50016 17836 50020
rect 17852 50076 17916 50080
rect 17852 50020 17856 50076
rect 17856 50020 17912 50076
rect 17912 50020 17916 50076
rect 17852 50016 17916 50020
rect 22612 50076 22676 50080
rect 22612 50020 22616 50076
rect 22616 50020 22672 50076
rect 22672 50020 22676 50076
rect 22612 50016 22676 50020
rect 22692 50076 22756 50080
rect 22692 50020 22696 50076
rect 22696 50020 22752 50076
rect 22752 50020 22756 50076
rect 22692 50016 22756 50020
rect 22772 50076 22836 50080
rect 22772 50020 22776 50076
rect 22776 50020 22832 50076
rect 22832 50020 22836 50076
rect 22772 50016 22836 50020
rect 22852 50076 22916 50080
rect 22852 50020 22856 50076
rect 22856 50020 22912 50076
rect 22912 50020 22916 50076
rect 22852 50016 22916 50020
rect 27612 50076 27676 50080
rect 27612 50020 27616 50076
rect 27616 50020 27672 50076
rect 27672 50020 27676 50076
rect 27612 50016 27676 50020
rect 27692 50076 27756 50080
rect 27692 50020 27696 50076
rect 27696 50020 27752 50076
rect 27752 50020 27756 50076
rect 27692 50016 27756 50020
rect 27772 50076 27836 50080
rect 27772 50020 27776 50076
rect 27776 50020 27832 50076
rect 27832 50020 27836 50076
rect 27772 50016 27836 50020
rect 27852 50076 27916 50080
rect 27852 50020 27856 50076
rect 27856 50020 27912 50076
rect 27912 50020 27916 50076
rect 27852 50016 27916 50020
rect 32612 50076 32676 50080
rect 32612 50020 32616 50076
rect 32616 50020 32672 50076
rect 32672 50020 32676 50076
rect 32612 50016 32676 50020
rect 32692 50076 32756 50080
rect 32692 50020 32696 50076
rect 32696 50020 32752 50076
rect 32752 50020 32756 50076
rect 32692 50016 32756 50020
rect 32772 50076 32836 50080
rect 32772 50020 32776 50076
rect 32776 50020 32832 50076
rect 32832 50020 32836 50076
rect 32772 50016 32836 50020
rect 32852 50076 32916 50080
rect 32852 50020 32856 50076
rect 32856 50020 32912 50076
rect 32912 50020 32916 50076
rect 32852 50016 32916 50020
rect 37612 50076 37676 50080
rect 37612 50020 37616 50076
rect 37616 50020 37672 50076
rect 37672 50020 37676 50076
rect 37612 50016 37676 50020
rect 37692 50076 37756 50080
rect 37692 50020 37696 50076
rect 37696 50020 37752 50076
rect 37752 50020 37756 50076
rect 37692 50016 37756 50020
rect 37772 50076 37836 50080
rect 37772 50020 37776 50076
rect 37776 50020 37832 50076
rect 37832 50020 37836 50076
rect 37772 50016 37836 50020
rect 37852 50076 37916 50080
rect 37852 50020 37856 50076
rect 37856 50020 37912 50076
rect 37912 50020 37916 50076
rect 37852 50016 37916 50020
rect 1952 49532 2016 49536
rect 1952 49476 1956 49532
rect 1956 49476 2012 49532
rect 2012 49476 2016 49532
rect 1952 49472 2016 49476
rect 2032 49532 2096 49536
rect 2032 49476 2036 49532
rect 2036 49476 2092 49532
rect 2092 49476 2096 49532
rect 2032 49472 2096 49476
rect 2112 49532 2176 49536
rect 2112 49476 2116 49532
rect 2116 49476 2172 49532
rect 2172 49476 2176 49532
rect 2112 49472 2176 49476
rect 2192 49532 2256 49536
rect 2192 49476 2196 49532
rect 2196 49476 2252 49532
rect 2252 49476 2256 49532
rect 2192 49472 2256 49476
rect 6952 49532 7016 49536
rect 6952 49476 6956 49532
rect 6956 49476 7012 49532
rect 7012 49476 7016 49532
rect 6952 49472 7016 49476
rect 7032 49532 7096 49536
rect 7032 49476 7036 49532
rect 7036 49476 7092 49532
rect 7092 49476 7096 49532
rect 7032 49472 7096 49476
rect 7112 49532 7176 49536
rect 7112 49476 7116 49532
rect 7116 49476 7172 49532
rect 7172 49476 7176 49532
rect 7112 49472 7176 49476
rect 7192 49532 7256 49536
rect 7192 49476 7196 49532
rect 7196 49476 7252 49532
rect 7252 49476 7256 49532
rect 7192 49472 7256 49476
rect 11952 49532 12016 49536
rect 11952 49476 11956 49532
rect 11956 49476 12012 49532
rect 12012 49476 12016 49532
rect 11952 49472 12016 49476
rect 12032 49532 12096 49536
rect 12032 49476 12036 49532
rect 12036 49476 12092 49532
rect 12092 49476 12096 49532
rect 12032 49472 12096 49476
rect 12112 49532 12176 49536
rect 12112 49476 12116 49532
rect 12116 49476 12172 49532
rect 12172 49476 12176 49532
rect 12112 49472 12176 49476
rect 12192 49532 12256 49536
rect 12192 49476 12196 49532
rect 12196 49476 12252 49532
rect 12252 49476 12256 49532
rect 12192 49472 12256 49476
rect 16952 49532 17016 49536
rect 16952 49476 16956 49532
rect 16956 49476 17012 49532
rect 17012 49476 17016 49532
rect 16952 49472 17016 49476
rect 17032 49532 17096 49536
rect 17032 49476 17036 49532
rect 17036 49476 17092 49532
rect 17092 49476 17096 49532
rect 17032 49472 17096 49476
rect 17112 49532 17176 49536
rect 17112 49476 17116 49532
rect 17116 49476 17172 49532
rect 17172 49476 17176 49532
rect 17112 49472 17176 49476
rect 17192 49532 17256 49536
rect 17192 49476 17196 49532
rect 17196 49476 17252 49532
rect 17252 49476 17256 49532
rect 17192 49472 17256 49476
rect 21952 49532 22016 49536
rect 21952 49476 21956 49532
rect 21956 49476 22012 49532
rect 22012 49476 22016 49532
rect 21952 49472 22016 49476
rect 22032 49532 22096 49536
rect 22032 49476 22036 49532
rect 22036 49476 22092 49532
rect 22092 49476 22096 49532
rect 22032 49472 22096 49476
rect 22112 49532 22176 49536
rect 22112 49476 22116 49532
rect 22116 49476 22172 49532
rect 22172 49476 22176 49532
rect 22112 49472 22176 49476
rect 22192 49532 22256 49536
rect 22192 49476 22196 49532
rect 22196 49476 22252 49532
rect 22252 49476 22256 49532
rect 22192 49472 22256 49476
rect 26952 49532 27016 49536
rect 26952 49476 26956 49532
rect 26956 49476 27012 49532
rect 27012 49476 27016 49532
rect 26952 49472 27016 49476
rect 27032 49532 27096 49536
rect 27032 49476 27036 49532
rect 27036 49476 27092 49532
rect 27092 49476 27096 49532
rect 27032 49472 27096 49476
rect 27112 49532 27176 49536
rect 27112 49476 27116 49532
rect 27116 49476 27172 49532
rect 27172 49476 27176 49532
rect 27112 49472 27176 49476
rect 27192 49532 27256 49536
rect 27192 49476 27196 49532
rect 27196 49476 27252 49532
rect 27252 49476 27256 49532
rect 27192 49472 27256 49476
rect 31952 49532 32016 49536
rect 31952 49476 31956 49532
rect 31956 49476 32012 49532
rect 32012 49476 32016 49532
rect 31952 49472 32016 49476
rect 32032 49532 32096 49536
rect 32032 49476 32036 49532
rect 32036 49476 32092 49532
rect 32092 49476 32096 49532
rect 32032 49472 32096 49476
rect 32112 49532 32176 49536
rect 32112 49476 32116 49532
rect 32116 49476 32172 49532
rect 32172 49476 32176 49532
rect 32112 49472 32176 49476
rect 32192 49532 32256 49536
rect 32192 49476 32196 49532
rect 32196 49476 32252 49532
rect 32252 49476 32256 49532
rect 32192 49472 32256 49476
rect 36952 49532 37016 49536
rect 36952 49476 36956 49532
rect 36956 49476 37012 49532
rect 37012 49476 37016 49532
rect 36952 49472 37016 49476
rect 37032 49532 37096 49536
rect 37032 49476 37036 49532
rect 37036 49476 37092 49532
rect 37092 49476 37096 49532
rect 37032 49472 37096 49476
rect 37112 49532 37176 49536
rect 37112 49476 37116 49532
rect 37116 49476 37172 49532
rect 37172 49476 37176 49532
rect 37112 49472 37176 49476
rect 37192 49532 37256 49536
rect 37192 49476 37196 49532
rect 37196 49476 37252 49532
rect 37252 49476 37256 49532
rect 37192 49472 37256 49476
rect 2612 48988 2676 48992
rect 2612 48932 2616 48988
rect 2616 48932 2672 48988
rect 2672 48932 2676 48988
rect 2612 48928 2676 48932
rect 2692 48988 2756 48992
rect 2692 48932 2696 48988
rect 2696 48932 2752 48988
rect 2752 48932 2756 48988
rect 2692 48928 2756 48932
rect 2772 48988 2836 48992
rect 2772 48932 2776 48988
rect 2776 48932 2832 48988
rect 2832 48932 2836 48988
rect 2772 48928 2836 48932
rect 2852 48988 2916 48992
rect 2852 48932 2856 48988
rect 2856 48932 2912 48988
rect 2912 48932 2916 48988
rect 2852 48928 2916 48932
rect 7612 48988 7676 48992
rect 7612 48932 7616 48988
rect 7616 48932 7672 48988
rect 7672 48932 7676 48988
rect 7612 48928 7676 48932
rect 7692 48988 7756 48992
rect 7692 48932 7696 48988
rect 7696 48932 7752 48988
rect 7752 48932 7756 48988
rect 7692 48928 7756 48932
rect 7772 48988 7836 48992
rect 7772 48932 7776 48988
rect 7776 48932 7832 48988
rect 7832 48932 7836 48988
rect 7772 48928 7836 48932
rect 7852 48988 7916 48992
rect 7852 48932 7856 48988
rect 7856 48932 7912 48988
rect 7912 48932 7916 48988
rect 7852 48928 7916 48932
rect 12612 48988 12676 48992
rect 12612 48932 12616 48988
rect 12616 48932 12672 48988
rect 12672 48932 12676 48988
rect 12612 48928 12676 48932
rect 12692 48988 12756 48992
rect 12692 48932 12696 48988
rect 12696 48932 12752 48988
rect 12752 48932 12756 48988
rect 12692 48928 12756 48932
rect 12772 48988 12836 48992
rect 12772 48932 12776 48988
rect 12776 48932 12832 48988
rect 12832 48932 12836 48988
rect 12772 48928 12836 48932
rect 12852 48988 12916 48992
rect 12852 48932 12856 48988
rect 12856 48932 12912 48988
rect 12912 48932 12916 48988
rect 12852 48928 12916 48932
rect 17612 48988 17676 48992
rect 17612 48932 17616 48988
rect 17616 48932 17672 48988
rect 17672 48932 17676 48988
rect 17612 48928 17676 48932
rect 17692 48988 17756 48992
rect 17692 48932 17696 48988
rect 17696 48932 17752 48988
rect 17752 48932 17756 48988
rect 17692 48928 17756 48932
rect 17772 48988 17836 48992
rect 17772 48932 17776 48988
rect 17776 48932 17832 48988
rect 17832 48932 17836 48988
rect 17772 48928 17836 48932
rect 17852 48988 17916 48992
rect 17852 48932 17856 48988
rect 17856 48932 17912 48988
rect 17912 48932 17916 48988
rect 17852 48928 17916 48932
rect 22612 48988 22676 48992
rect 22612 48932 22616 48988
rect 22616 48932 22672 48988
rect 22672 48932 22676 48988
rect 22612 48928 22676 48932
rect 22692 48988 22756 48992
rect 22692 48932 22696 48988
rect 22696 48932 22752 48988
rect 22752 48932 22756 48988
rect 22692 48928 22756 48932
rect 22772 48988 22836 48992
rect 22772 48932 22776 48988
rect 22776 48932 22832 48988
rect 22832 48932 22836 48988
rect 22772 48928 22836 48932
rect 22852 48988 22916 48992
rect 22852 48932 22856 48988
rect 22856 48932 22912 48988
rect 22912 48932 22916 48988
rect 22852 48928 22916 48932
rect 27612 48988 27676 48992
rect 27612 48932 27616 48988
rect 27616 48932 27672 48988
rect 27672 48932 27676 48988
rect 27612 48928 27676 48932
rect 27692 48988 27756 48992
rect 27692 48932 27696 48988
rect 27696 48932 27752 48988
rect 27752 48932 27756 48988
rect 27692 48928 27756 48932
rect 27772 48988 27836 48992
rect 27772 48932 27776 48988
rect 27776 48932 27832 48988
rect 27832 48932 27836 48988
rect 27772 48928 27836 48932
rect 27852 48988 27916 48992
rect 27852 48932 27856 48988
rect 27856 48932 27912 48988
rect 27912 48932 27916 48988
rect 27852 48928 27916 48932
rect 32612 48988 32676 48992
rect 32612 48932 32616 48988
rect 32616 48932 32672 48988
rect 32672 48932 32676 48988
rect 32612 48928 32676 48932
rect 32692 48988 32756 48992
rect 32692 48932 32696 48988
rect 32696 48932 32752 48988
rect 32752 48932 32756 48988
rect 32692 48928 32756 48932
rect 32772 48988 32836 48992
rect 32772 48932 32776 48988
rect 32776 48932 32832 48988
rect 32832 48932 32836 48988
rect 32772 48928 32836 48932
rect 32852 48988 32916 48992
rect 32852 48932 32856 48988
rect 32856 48932 32912 48988
rect 32912 48932 32916 48988
rect 32852 48928 32916 48932
rect 37612 48988 37676 48992
rect 37612 48932 37616 48988
rect 37616 48932 37672 48988
rect 37672 48932 37676 48988
rect 37612 48928 37676 48932
rect 37692 48988 37756 48992
rect 37692 48932 37696 48988
rect 37696 48932 37752 48988
rect 37752 48932 37756 48988
rect 37692 48928 37756 48932
rect 37772 48988 37836 48992
rect 37772 48932 37776 48988
rect 37776 48932 37832 48988
rect 37832 48932 37836 48988
rect 37772 48928 37836 48932
rect 37852 48988 37916 48992
rect 37852 48932 37856 48988
rect 37856 48932 37912 48988
rect 37912 48932 37916 48988
rect 37852 48928 37916 48932
rect 1952 48444 2016 48448
rect 1952 48388 1956 48444
rect 1956 48388 2012 48444
rect 2012 48388 2016 48444
rect 1952 48384 2016 48388
rect 2032 48444 2096 48448
rect 2032 48388 2036 48444
rect 2036 48388 2092 48444
rect 2092 48388 2096 48444
rect 2032 48384 2096 48388
rect 2112 48444 2176 48448
rect 2112 48388 2116 48444
rect 2116 48388 2172 48444
rect 2172 48388 2176 48444
rect 2112 48384 2176 48388
rect 2192 48444 2256 48448
rect 2192 48388 2196 48444
rect 2196 48388 2252 48444
rect 2252 48388 2256 48444
rect 2192 48384 2256 48388
rect 6952 48444 7016 48448
rect 6952 48388 6956 48444
rect 6956 48388 7012 48444
rect 7012 48388 7016 48444
rect 6952 48384 7016 48388
rect 7032 48444 7096 48448
rect 7032 48388 7036 48444
rect 7036 48388 7092 48444
rect 7092 48388 7096 48444
rect 7032 48384 7096 48388
rect 7112 48444 7176 48448
rect 7112 48388 7116 48444
rect 7116 48388 7172 48444
rect 7172 48388 7176 48444
rect 7112 48384 7176 48388
rect 7192 48444 7256 48448
rect 7192 48388 7196 48444
rect 7196 48388 7252 48444
rect 7252 48388 7256 48444
rect 7192 48384 7256 48388
rect 11952 48444 12016 48448
rect 11952 48388 11956 48444
rect 11956 48388 12012 48444
rect 12012 48388 12016 48444
rect 11952 48384 12016 48388
rect 12032 48444 12096 48448
rect 12032 48388 12036 48444
rect 12036 48388 12092 48444
rect 12092 48388 12096 48444
rect 12032 48384 12096 48388
rect 12112 48444 12176 48448
rect 12112 48388 12116 48444
rect 12116 48388 12172 48444
rect 12172 48388 12176 48444
rect 12112 48384 12176 48388
rect 12192 48444 12256 48448
rect 12192 48388 12196 48444
rect 12196 48388 12252 48444
rect 12252 48388 12256 48444
rect 12192 48384 12256 48388
rect 16952 48444 17016 48448
rect 16952 48388 16956 48444
rect 16956 48388 17012 48444
rect 17012 48388 17016 48444
rect 16952 48384 17016 48388
rect 17032 48444 17096 48448
rect 17032 48388 17036 48444
rect 17036 48388 17092 48444
rect 17092 48388 17096 48444
rect 17032 48384 17096 48388
rect 17112 48444 17176 48448
rect 17112 48388 17116 48444
rect 17116 48388 17172 48444
rect 17172 48388 17176 48444
rect 17112 48384 17176 48388
rect 17192 48444 17256 48448
rect 17192 48388 17196 48444
rect 17196 48388 17252 48444
rect 17252 48388 17256 48444
rect 17192 48384 17256 48388
rect 21952 48444 22016 48448
rect 21952 48388 21956 48444
rect 21956 48388 22012 48444
rect 22012 48388 22016 48444
rect 21952 48384 22016 48388
rect 22032 48444 22096 48448
rect 22032 48388 22036 48444
rect 22036 48388 22092 48444
rect 22092 48388 22096 48444
rect 22032 48384 22096 48388
rect 22112 48444 22176 48448
rect 22112 48388 22116 48444
rect 22116 48388 22172 48444
rect 22172 48388 22176 48444
rect 22112 48384 22176 48388
rect 22192 48444 22256 48448
rect 22192 48388 22196 48444
rect 22196 48388 22252 48444
rect 22252 48388 22256 48444
rect 22192 48384 22256 48388
rect 26952 48444 27016 48448
rect 26952 48388 26956 48444
rect 26956 48388 27012 48444
rect 27012 48388 27016 48444
rect 26952 48384 27016 48388
rect 27032 48444 27096 48448
rect 27032 48388 27036 48444
rect 27036 48388 27092 48444
rect 27092 48388 27096 48444
rect 27032 48384 27096 48388
rect 27112 48444 27176 48448
rect 27112 48388 27116 48444
rect 27116 48388 27172 48444
rect 27172 48388 27176 48444
rect 27112 48384 27176 48388
rect 27192 48444 27256 48448
rect 27192 48388 27196 48444
rect 27196 48388 27252 48444
rect 27252 48388 27256 48444
rect 27192 48384 27256 48388
rect 31952 48444 32016 48448
rect 31952 48388 31956 48444
rect 31956 48388 32012 48444
rect 32012 48388 32016 48444
rect 31952 48384 32016 48388
rect 32032 48444 32096 48448
rect 32032 48388 32036 48444
rect 32036 48388 32092 48444
rect 32092 48388 32096 48444
rect 32032 48384 32096 48388
rect 32112 48444 32176 48448
rect 32112 48388 32116 48444
rect 32116 48388 32172 48444
rect 32172 48388 32176 48444
rect 32112 48384 32176 48388
rect 32192 48444 32256 48448
rect 32192 48388 32196 48444
rect 32196 48388 32252 48444
rect 32252 48388 32256 48444
rect 32192 48384 32256 48388
rect 36952 48444 37016 48448
rect 36952 48388 36956 48444
rect 36956 48388 37012 48444
rect 37012 48388 37016 48444
rect 36952 48384 37016 48388
rect 37032 48444 37096 48448
rect 37032 48388 37036 48444
rect 37036 48388 37092 48444
rect 37092 48388 37096 48444
rect 37032 48384 37096 48388
rect 37112 48444 37176 48448
rect 37112 48388 37116 48444
rect 37116 48388 37172 48444
rect 37172 48388 37176 48444
rect 37112 48384 37176 48388
rect 37192 48444 37256 48448
rect 37192 48388 37196 48444
rect 37196 48388 37252 48444
rect 37252 48388 37256 48444
rect 37192 48384 37256 48388
rect 2612 47900 2676 47904
rect 2612 47844 2616 47900
rect 2616 47844 2672 47900
rect 2672 47844 2676 47900
rect 2612 47840 2676 47844
rect 2692 47900 2756 47904
rect 2692 47844 2696 47900
rect 2696 47844 2752 47900
rect 2752 47844 2756 47900
rect 2692 47840 2756 47844
rect 2772 47900 2836 47904
rect 2772 47844 2776 47900
rect 2776 47844 2832 47900
rect 2832 47844 2836 47900
rect 2772 47840 2836 47844
rect 2852 47900 2916 47904
rect 2852 47844 2856 47900
rect 2856 47844 2912 47900
rect 2912 47844 2916 47900
rect 2852 47840 2916 47844
rect 7612 47900 7676 47904
rect 7612 47844 7616 47900
rect 7616 47844 7672 47900
rect 7672 47844 7676 47900
rect 7612 47840 7676 47844
rect 7692 47900 7756 47904
rect 7692 47844 7696 47900
rect 7696 47844 7752 47900
rect 7752 47844 7756 47900
rect 7692 47840 7756 47844
rect 7772 47900 7836 47904
rect 7772 47844 7776 47900
rect 7776 47844 7832 47900
rect 7832 47844 7836 47900
rect 7772 47840 7836 47844
rect 7852 47900 7916 47904
rect 7852 47844 7856 47900
rect 7856 47844 7912 47900
rect 7912 47844 7916 47900
rect 7852 47840 7916 47844
rect 12612 47900 12676 47904
rect 12612 47844 12616 47900
rect 12616 47844 12672 47900
rect 12672 47844 12676 47900
rect 12612 47840 12676 47844
rect 12692 47900 12756 47904
rect 12692 47844 12696 47900
rect 12696 47844 12752 47900
rect 12752 47844 12756 47900
rect 12692 47840 12756 47844
rect 12772 47900 12836 47904
rect 12772 47844 12776 47900
rect 12776 47844 12832 47900
rect 12832 47844 12836 47900
rect 12772 47840 12836 47844
rect 12852 47900 12916 47904
rect 12852 47844 12856 47900
rect 12856 47844 12912 47900
rect 12912 47844 12916 47900
rect 12852 47840 12916 47844
rect 17612 47900 17676 47904
rect 17612 47844 17616 47900
rect 17616 47844 17672 47900
rect 17672 47844 17676 47900
rect 17612 47840 17676 47844
rect 17692 47900 17756 47904
rect 17692 47844 17696 47900
rect 17696 47844 17752 47900
rect 17752 47844 17756 47900
rect 17692 47840 17756 47844
rect 17772 47900 17836 47904
rect 17772 47844 17776 47900
rect 17776 47844 17832 47900
rect 17832 47844 17836 47900
rect 17772 47840 17836 47844
rect 17852 47900 17916 47904
rect 17852 47844 17856 47900
rect 17856 47844 17912 47900
rect 17912 47844 17916 47900
rect 17852 47840 17916 47844
rect 22612 47900 22676 47904
rect 22612 47844 22616 47900
rect 22616 47844 22672 47900
rect 22672 47844 22676 47900
rect 22612 47840 22676 47844
rect 22692 47900 22756 47904
rect 22692 47844 22696 47900
rect 22696 47844 22752 47900
rect 22752 47844 22756 47900
rect 22692 47840 22756 47844
rect 22772 47900 22836 47904
rect 22772 47844 22776 47900
rect 22776 47844 22832 47900
rect 22832 47844 22836 47900
rect 22772 47840 22836 47844
rect 22852 47900 22916 47904
rect 22852 47844 22856 47900
rect 22856 47844 22912 47900
rect 22912 47844 22916 47900
rect 22852 47840 22916 47844
rect 27612 47900 27676 47904
rect 27612 47844 27616 47900
rect 27616 47844 27672 47900
rect 27672 47844 27676 47900
rect 27612 47840 27676 47844
rect 27692 47900 27756 47904
rect 27692 47844 27696 47900
rect 27696 47844 27752 47900
rect 27752 47844 27756 47900
rect 27692 47840 27756 47844
rect 27772 47900 27836 47904
rect 27772 47844 27776 47900
rect 27776 47844 27832 47900
rect 27832 47844 27836 47900
rect 27772 47840 27836 47844
rect 27852 47900 27916 47904
rect 27852 47844 27856 47900
rect 27856 47844 27912 47900
rect 27912 47844 27916 47900
rect 27852 47840 27916 47844
rect 32612 47900 32676 47904
rect 32612 47844 32616 47900
rect 32616 47844 32672 47900
rect 32672 47844 32676 47900
rect 32612 47840 32676 47844
rect 32692 47900 32756 47904
rect 32692 47844 32696 47900
rect 32696 47844 32752 47900
rect 32752 47844 32756 47900
rect 32692 47840 32756 47844
rect 32772 47900 32836 47904
rect 32772 47844 32776 47900
rect 32776 47844 32832 47900
rect 32832 47844 32836 47900
rect 32772 47840 32836 47844
rect 32852 47900 32916 47904
rect 32852 47844 32856 47900
rect 32856 47844 32912 47900
rect 32912 47844 32916 47900
rect 32852 47840 32916 47844
rect 37612 47900 37676 47904
rect 37612 47844 37616 47900
rect 37616 47844 37672 47900
rect 37672 47844 37676 47900
rect 37612 47840 37676 47844
rect 37692 47900 37756 47904
rect 37692 47844 37696 47900
rect 37696 47844 37752 47900
rect 37752 47844 37756 47900
rect 37692 47840 37756 47844
rect 37772 47900 37836 47904
rect 37772 47844 37776 47900
rect 37776 47844 37832 47900
rect 37832 47844 37836 47900
rect 37772 47840 37836 47844
rect 37852 47900 37916 47904
rect 37852 47844 37856 47900
rect 37856 47844 37912 47900
rect 37912 47844 37916 47900
rect 37852 47840 37916 47844
rect 1952 47356 2016 47360
rect 1952 47300 1956 47356
rect 1956 47300 2012 47356
rect 2012 47300 2016 47356
rect 1952 47296 2016 47300
rect 2032 47356 2096 47360
rect 2032 47300 2036 47356
rect 2036 47300 2092 47356
rect 2092 47300 2096 47356
rect 2032 47296 2096 47300
rect 2112 47356 2176 47360
rect 2112 47300 2116 47356
rect 2116 47300 2172 47356
rect 2172 47300 2176 47356
rect 2112 47296 2176 47300
rect 2192 47356 2256 47360
rect 2192 47300 2196 47356
rect 2196 47300 2252 47356
rect 2252 47300 2256 47356
rect 2192 47296 2256 47300
rect 6952 47356 7016 47360
rect 6952 47300 6956 47356
rect 6956 47300 7012 47356
rect 7012 47300 7016 47356
rect 6952 47296 7016 47300
rect 7032 47356 7096 47360
rect 7032 47300 7036 47356
rect 7036 47300 7092 47356
rect 7092 47300 7096 47356
rect 7032 47296 7096 47300
rect 7112 47356 7176 47360
rect 7112 47300 7116 47356
rect 7116 47300 7172 47356
rect 7172 47300 7176 47356
rect 7112 47296 7176 47300
rect 7192 47356 7256 47360
rect 7192 47300 7196 47356
rect 7196 47300 7252 47356
rect 7252 47300 7256 47356
rect 7192 47296 7256 47300
rect 11952 47356 12016 47360
rect 11952 47300 11956 47356
rect 11956 47300 12012 47356
rect 12012 47300 12016 47356
rect 11952 47296 12016 47300
rect 12032 47356 12096 47360
rect 12032 47300 12036 47356
rect 12036 47300 12092 47356
rect 12092 47300 12096 47356
rect 12032 47296 12096 47300
rect 12112 47356 12176 47360
rect 12112 47300 12116 47356
rect 12116 47300 12172 47356
rect 12172 47300 12176 47356
rect 12112 47296 12176 47300
rect 12192 47356 12256 47360
rect 12192 47300 12196 47356
rect 12196 47300 12252 47356
rect 12252 47300 12256 47356
rect 12192 47296 12256 47300
rect 16952 47356 17016 47360
rect 16952 47300 16956 47356
rect 16956 47300 17012 47356
rect 17012 47300 17016 47356
rect 16952 47296 17016 47300
rect 17032 47356 17096 47360
rect 17032 47300 17036 47356
rect 17036 47300 17092 47356
rect 17092 47300 17096 47356
rect 17032 47296 17096 47300
rect 17112 47356 17176 47360
rect 17112 47300 17116 47356
rect 17116 47300 17172 47356
rect 17172 47300 17176 47356
rect 17112 47296 17176 47300
rect 17192 47356 17256 47360
rect 17192 47300 17196 47356
rect 17196 47300 17252 47356
rect 17252 47300 17256 47356
rect 17192 47296 17256 47300
rect 21952 47356 22016 47360
rect 21952 47300 21956 47356
rect 21956 47300 22012 47356
rect 22012 47300 22016 47356
rect 21952 47296 22016 47300
rect 22032 47356 22096 47360
rect 22032 47300 22036 47356
rect 22036 47300 22092 47356
rect 22092 47300 22096 47356
rect 22032 47296 22096 47300
rect 22112 47356 22176 47360
rect 22112 47300 22116 47356
rect 22116 47300 22172 47356
rect 22172 47300 22176 47356
rect 22112 47296 22176 47300
rect 22192 47356 22256 47360
rect 22192 47300 22196 47356
rect 22196 47300 22252 47356
rect 22252 47300 22256 47356
rect 22192 47296 22256 47300
rect 26952 47356 27016 47360
rect 26952 47300 26956 47356
rect 26956 47300 27012 47356
rect 27012 47300 27016 47356
rect 26952 47296 27016 47300
rect 27032 47356 27096 47360
rect 27032 47300 27036 47356
rect 27036 47300 27092 47356
rect 27092 47300 27096 47356
rect 27032 47296 27096 47300
rect 27112 47356 27176 47360
rect 27112 47300 27116 47356
rect 27116 47300 27172 47356
rect 27172 47300 27176 47356
rect 27112 47296 27176 47300
rect 27192 47356 27256 47360
rect 27192 47300 27196 47356
rect 27196 47300 27252 47356
rect 27252 47300 27256 47356
rect 27192 47296 27256 47300
rect 31952 47356 32016 47360
rect 31952 47300 31956 47356
rect 31956 47300 32012 47356
rect 32012 47300 32016 47356
rect 31952 47296 32016 47300
rect 32032 47356 32096 47360
rect 32032 47300 32036 47356
rect 32036 47300 32092 47356
rect 32092 47300 32096 47356
rect 32032 47296 32096 47300
rect 32112 47356 32176 47360
rect 32112 47300 32116 47356
rect 32116 47300 32172 47356
rect 32172 47300 32176 47356
rect 32112 47296 32176 47300
rect 32192 47356 32256 47360
rect 32192 47300 32196 47356
rect 32196 47300 32252 47356
rect 32252 47300 32256 47356
rect 32192 47296 32256 47300
rect 36952 47356 37016 47360
rect 36952 47300 36956 47356
rect 36956 47300 37012 47356
rect 37012 47300 37016 47356
rect 36952 47296 37016 47300
rect 37032 47356 37096 47360
rect 37032 47300 37036 47356
rect 37036 47300 37092 47356
rect 37092 47300 37096 47356
rect 37032 47296 37096 47300
rect 37112 47356 37176 47360
rect 37112 47300 37116 47356
rect 37116 47300 37172 47356
rect 37172 47300 37176 47356
rect 37112 47296 37176 47300
rect 37192 47356 37256 47360
rect 37192 47300 37196 47356
rect 37196 47300 37252 47356
rect 37252 47300 37256 47356
rect 37192 47296 37256 47300
rect 2612 46812 2676 46816
rect 2612 46756 2616 46812
rect 2616 46756 2672 46812
rect 2672 46756 2676 46812
rect 2612 46752 2676 46756
rect 2692 46812 2756 46816
rect 2692 46756 2696 46812
rect 2696 46756 2752 46812
rect 2752 46756 2756 46812
rect 2692 46752 2756 46756
rect 2772 46812 2836 46816
rect 2772 46756 2776 46812
rect 2776 46756 2832 46812
rect 2832 46756 2836 46812
rect 2772 46752 2836 46756
rect 2852 46812 2916 46816
rect 2852 46756 2856 46812
rect 2856 46756 2912 46812
rect 2912 46756 2916 46812
rect 2852 46752 2916 46756
rect 7612 46812 7676 46816
rect 7612 46756 7616 46812
rect 7616 46756 7672 46812
rect 7672 46756 7676 46812
rect 7612 46752 7676 46756
rect 7692 46812 7756 46816
rect 7692 46756 7696 46812
rect 7696 46756 7752 46812
rect 7752 46756 7756 46812
rect 7692 46752 7756 46756
rect 7772 46812 7836 46816
rect 7772 46756 7776 46812
rect 7776 46756 7832 46812
rect 7832 46756 7836 46812
rect 7772 46752 7836 46756
rect 7852 46812 7916 46816
rect 7852 46756 7856 46812
rect 7856 46756 7912 46812
rect 7912 46756 7916 46812
rect 7852 46752 7916 46756
rect 12612 46812 12676 46816
rect 12612 46756 12616 46812
rect 12616 46756 12672 46812
rect 12672 46756 12676 46812
rect 12612 46752 12676 46756
rect 12692 46812 12756 46816
rect 12692 46756 12696 46812
rect 12696 46756 12752 46812
rect 12752 46756 12756 46812
rect 12692 46752 12756 46756
rect 12772 46812 12836 46816
rect 12772 46756 12776 46812
rect 12776 46756 12832 46812
rect 12832 46756 12836 46812
rect 12772 46752 12836 46756
rect 12852 46812 12916 46816
rect 12852 46756 12856 46812
rect 12856 46756 12912 46812
rect 12912 46756 12916 46812
rect 12852 46752 12916 46756
rect 17612 46812 17676 46816
rect 17612 46756 17616 46812
rect 17616 46756 17672 46812
rect 17672 46756 17676 46812
rect 17612 46752 17676 46756
rect 17692 46812 17756 46816
rect 17692 46756 17696 46812
rect 17696 46756 17752 46812
rect 17752 46756 17756 46812
rect 17692 46752 17756 46756
rect 17772 46812 17836 46816
rect 17772 46756 17776 46812
rect 17776 46756 17832 46812
rect 17832 46756 17836 46812
rect 17772 46752 17836 46756
rect 17852 46812 17916 46816
rect 17852 46756 17856 46812
rect 17856 46756 17912 46812
rect 17912 46756 17916 46812
rect 17852 46752 17916 46756
rect 22612 46812 22676 46816
rect 22612 46756 22616 46812
rect 22616 46756 22672 46812
rect 22672 46756 22676 46812
rect 22612 46752 22676 46756
rect 22692 46812 22756 46816
rect 22692 46756 22696 46812
rect 22696 46756 22752 46812
rect 22752 46756 22756 46812
rect 22692 46752 22756 46756
rect 22772 46812 22836 46816
rect 22772 46756 22776 46812
rect 22776 46756 22832 46812
rect 22832 46756 22836 46812
rect 22772 46752 22836 46756
rect 22852 46812 22916 46816
rect 22852 46756 22856 46812
rect 22856 46756 22912 46812
rect 22912 46756 22916 46812
rect 22852 46752 22916 46756
rect 27612 46812 27676 46816
rect 27612 46756 27616 46812
rect 27616 46756 27672 46812
rect 27672 46756 27676 46812
rect 27612 46752 27676 46756
rect 27692 46812 27756 46816
rect 27692 46756 27696 46812
rect 27696 46756 27752 46812
rect 27752 46756 27756 46812
rect 27692 46752 27756 46756
rect 27772 46812 27836 46816
rect 27772 46756 27776 46812
rect 27776 46756 27832 46812
rect 27832 46756 27836 46812
rect 27772 46752 27836 46756
rect 27852 46812 27916 46816
rect 27852 46756 27856 46812
rect 27856 46756 27912 46812
rect 27912 46756 27916 46812
rect 27852 46752 27916 46756
rect 32612 46812 32676 46816
rect 32612 46756 32616 46812
rect 32616 46756 32672 46812
rect 32672 46756 32676 46812
rect 32612 46752 32676 46756
rect 32692 46812 32756 46816
rect 32692 46756 32696 46812
rect 32696 46756 32752 46812
rect 32752 46756 32756 46812
rect 32692 46752 32756 46756
rect 32772 46812 32836 46816
rect 32772 46756 32776 46812
rect 32776 46756 32832 46812
rect 32832 46756 32836 46812
rect 32772 46752 32836 46756
rect 32852 46812 32916 46816
rect 32852 46756 32856 46812
rect 32856 46756 32912 46812
rect 32912 46756 32916 46812
rect 32852 46752 32916 46756
rect 37612 46812 37676 46816
rect 37612 46756 37616 46812
rect 37616 46756 37672 46812
rect 37672 46756 37676 46812
rect 37612 46752 37676 46756
rect 37692 46812 37756 46816
rect 37692 46756 37696 46812
rect 37696 46756 37752 46812
rect 37752 46756 37756 46812
rect 37692 46752 37756 46756
rect 37772 46812 37836 46816
rect 37772 46756 37776 46812
rect 37776 46756 37832 46812
rect 37832 46756 37836 46812
rect 37772 46752 37836 46756
rect 37852 46812 37916 46816
rect 37852 46756 37856 46812
rect 37856 46756 37912 46812
rect 37912 46756 37916 46812
rect 37852 46752 37916 46756
rect 1952 46268 2016 46272
rect 1952 46212 1956 46268
rect 1956 46212 2012 46268
rect 2012 46212 2016 46268
rect 1952 46208 2016 46212
rect 2032 46268 2096 46272
rect 2032 46212 2036 46268
rect 2036 46212 2092 46268
rect 2092 46212 2096 46268
rect 2032 46208 2096 46212
rect 2112 46268 2176 46272
rect 2112 46212 2116 46268
rect 2116 46212 2172 46268
rect 2172 46212 2176 46268
rect 2112 46208 2176 46212
rect 2192 46268 2256 46272
rect 2192 46212 2196 46268
rect 2196 46212 2252 46268
rect 2252 46212 2256 46268
rect 2192 46208 2256 46212
rect 6952 46268 7016 46272
rect 6952 46212 6956 46268
rect 6956 46212 7012 46268
rect 7012 46212 7016 46268
rect 6952 46208 7016 46212
rect 7032 46268 7096 46272
rect 7032 46212 7036 46268
rect 7036 46212 7092 46268
rect 7092 46212 7096 46268
rect 7032 46208 7096 46212
rect 7112 46268 7176 46272
rect 7112 46212 7116 46268
rect 7116 46212 7172 46268
rect 7172 46212 7176 46268
rect 7112 46208 7176 46212
rect 7192 46268 7256 46272
rect 7192 46212 7196 46268
rect 7196 46212 7252 46268
rect 7252 46212 7256 46268
rect 7192 46208 7256 46212
rect 11952 46268 12016 46272
rect 11952 46212 11956 46268
rect 11956 46212 12012 46268
rect 12012 46212 12016 46268
rect 11952 46208 12016 46212
rect 12032 46268 12096 46272
rect 12032 46212 12036 46268
rect 12036 46212 12092 46268
rect 12092 46212 12096 46268
rect 12032 46208 12096 46212
rect 12112 46268 12176 46272
rect 12112 46212 12116 46268
rect 12116 46212 12172 46268
rect 12172 46212 12176 46268
rect 12112 46208 12176 46212
rect 12192 46268 12256 46272
rect 12192 46212 12196 46268
rect 12196 46212 12252 46268
rect 12252 46212 12256 46268
rect 12192 46208 12256 46212
rect 16952 46268 17016 46272
rect 16952 46212 16956 46268
rect 16956 46212 17012 46268
rect 17012 46212 17016 46268
rect 16952 46208 17016 46212
rect 17032 46268 17096 46272
rect 17032 46212 17036 46268
rect 17036 46212 17092 46268
rect 17092 46212 17096 46268
rect 17032 46208 17096 46212
rect 17112 46268 17176 46272
rect 17112 46212 17116 46268
rect 17116 46212 17172 46268
rect 17172 46212 17176 46268
rect 17112 46208 17176 46212
rect 17192 46268 17256 46272
rect 17192 46212 17196 46268
rect 17196 46212 17252 46268
rect 17252 46212 17256 46268
rect 17192 46208 17256 46212
rect 21952 46268 22016 46272
rect 21952 46212 21956 46268
rect 21956 46212 22012 46268
rect 22012 46212 22016 46268
rect 21952 46208 22016 46212
rect 22032 46268 22096 46272
rect 22032 46212 22036 46268
rect 22036 46212 22092 46268
rect 22092 46212 22096 46268
rect 22032 46208 22096 46212
rect 22112 46268 22176 46272
rect 22112 46212 22116 46268
rect 22116 46212 22172 46268
rect 22172 46212 22176 46268
rect 22112 46208 22176 46212
rect 22192 46268 22256 46272
rect 22192 46212 22196 46268
rect 22196 46212 22252 46268
rect 22252 46212 22256 46268
rect 22192 46208 22256 46212
rect 26952 46268 27016 46272
rect 26952 46212 26956 46268
rect 26956 46212 27012 46268
rect 27012 46212 27016 46268
rect 26952 46208 27016 46212
rect 27032 46268 27096 46272
rect 27032 46212 27036 46268
rect 27036 46212 27092 46268
rect 27092 46212 27096 46268
rect 27032 46208 27096 46212
rect 27112 46268 27176 46272
rect 27112 46212 27116 46268
rect 27116 46212 27172 46268
rect 27172 46212 27176 46268
rect 27112 46208 27176 46212
rect 27192 46268 27256 46272
rect 27192 46212 27196 46268
rect 27196 46212 27252 46268
rect 27252 46212 27256 46268
rect 27192 46208 27256 46212
rect 31952 46268 32016 46272
rect 31952 46212 31956 46268
rect 31956 46212 32012 46268
rect 32012 46212 32016 46268
rect 31952 46208 32016 46212
rect 32032 46268 32096 46272
rect 32032 46212 32036 46268
rect 32036 46212 32092 46268
rect 32092 46212 32096 46268
rect 32032 46208 32096 46212
rect 32112 46268 32176 46272
rect 32112 46212 32116 46268
rect 32116 46212 32172 46268
rect 32172 46212 32176 46268
rect 32112 46208 32176 46212
rect 32192 46268 32256 46272
rect 32192 46212 32196 46268
rect 32196 46212 32252 46268
rect 32252 46212 32256 46268
rect 32192 46208 32256 46212
rect 36952 46268 37016 46272
rect 36952 46212 36956 46268
rect 36956 46212 37012 46268
rect 37012 46212 37016 46268
rect 36952 46208 37016 46212
rect 37032 46268 37096 46272
rect 37032 46212 37036 46268
rect 37036 46212 37092 46268
rect 37092 46212 37096 46268
rect 37032 46208 37096 46212
rect 37112 46268 37176 46272
rect 37112 46212 37116 46268
rect 37116 46212 37172 46268
rect 37172 46212 37176 46268
rect 37112 46208 37176 46212
rect 37192 46268 37256 46272
rect 37192 46212 37196 46268
rect 37196 46212 37252 46268
rect 37252 46212 37256 46268
rect 37192 46208 37256 46212
rect 21036 45868 21100 45932
rect 2612 45724 2676 45728
rect 2612 45668 2616 45724
rect 2616 45668 2672 45724
rect 2672 45668 2676 45724
rect 2612 45664 2676 45668
rect 2692 45724 2756 45728
rect 2692 45668 2696 45724
rect 2696 45668 2752 45724
rect 2752 45668 2756 45724
rect 2692 45664 2756 45668
rect 2772 45724 2836 45728
rect 2772 45668 2776 45724
rect 2776 45668 2832 45724
rect 2832 45668 2836 45724
rect 2772 45664 2836 45668
rect 2852 45724 2916 45728
rect 2852 45668 2856 45724
rect 2856 45668 2912 45724
rect 2912 45668 2916 45724
rect 2852 45664 2916 45668
rect 7612 45724 7676 45728
rect 7612 45668 7616 45724
rect 7616 45668 7672 45724
rect 7672 45668 7676 45724
rect 7612 45664 7676 45668
rect 7692 45724 7756 45728
rect 7692 45668 7696 45724
rect 7696 45668 7752 45724
rect 7752 45668 7756 45724
rect 7692 45664 7756 45668
rect 7772 45724 7836 45728
rect 7772 45668 7776 45724
rect 7776 45668 7832 45724
rect 7832 45668 7836 45724
rect 7772 45664 7836 45668
rect 7852 45724 7916 45728
rect 7852 45668 7856 45724
rect 7856 45668 7912 45724
rect 7912 45668 7916 45724
rect 7852 45664 7916 45668
rect 12612 45724 12676 45728
rect 12612 45668 12616 45724
rect 12616 45668 12672 45724
rect 12672 45668 12676 45724
rect 12612 45664 12676 45668
rect 12692 45724 12756 45728
rect 12692 45668 12696 45724
rect 12696 45668 12752 45724
rect 12752 45668 12756 45724
rect 12692 45664 12756 45668
rect 12772 45724 12836 45728
rect 12772 45668 12776 45724
rect 12776 45668 12832 45724
rect 12832 45668 12836 45724
rect 12772 45664 12836 45668
rect 12852 45724 12916 45728
rect 12852 45668 12856 45724
rect 12856 45668 12912 45724
rect 12912 45668 12916 45724
rect 12852 45664 12916 45668
rect 17612 45724 17676 45728
rect 17612 45668 17616 45724
rect 17616 45668 17672 45724
rect 17672 45668 17676 45724
rect 17612 45664 17676 45668
rect 17692 45724 17756 45728
rect 17692 45668 17696 45724
rect 17696 45668 17752 45724
rect 17752 45668 17756 45724
rect 17692 45664 17756 45668
rect 17772 45724 17836 45728
rect 17772 45668 17776 45724
rect 17776 45668 17832 45724
rect 17832 45668 17836 45724
rect 17772 45664 17836 45668
rect 17852 45724 17916 45728
rect 17852 45668 17856 45724
rect 17856 45668 17912 45724
rect 17912 45668 17916 45724
rect 17852 45664 17916 45668
rect 22612 45724 22676 45728
rect 22612 45668 22616 45724
rect 22616 45668 22672 45724
rect 22672 45668 22676 45724
rect 22612 45664 22676 45668
rect 22692 45724 22756 45728
rect 22692 45668 22696 45724
rect 22696 45668 22752 45724
rect 22752 45668 22756 45724
rect 22692 45664 22756 45668
rect 22772 45724 22836 45728
rect 22772 45668 22776 45724
rect 22776 45668 22832 45724
rect 22832 45668 22836 45724
rect 22772 45664 22836 45668
rect 22852 45724 22916 45728
rect 22852 45668 22856 45724
rect 22856 45668 22912 45724
rect 22912 45668 22916 45724
rect 22852 45664 22916 45668
rect 27612 45724 27676 45728
rect 27612 45668 27616 45724
rect 27616 45668 27672 45724
rect 27672 45668 27676 45724
rect 27612 45664 27676 45668
rect 27692 45724 27756 45728
rect 27692 45668 27696 45724
rect 27696 45668 27752 45724
rect 27752 45668 27756 45724
rect 27692 45664 27756 45668
rect 27772 45724 27836 45728
rect 27772 45668 27776 45724
rect 27776 45668 27832 45724
rect 27832 45668 27836 45724
rect 27772 45664 27836 45668
rect 27852 45724 27916 45728
rect 27852 45668 27856 45724
rect 27856 45668 27912 45724
rect 27912 45668 27916 45724
rect 27852 45664 27916 45668
rect 32612 45724 32676 45728
rect 32612 45668 32616 45724
rect 32616 45668 32672 45724
rect 32672 45668 32676 45724
rect 32612 45664 32676 45668
rect 32692 45724 32756 45728
rect 32692 45668 32696 45724
rect 32696 45668 32752 45724
rect 32752 45668 32756 45724
rect 32692 45664 32756 45668
rect 32772 45724 32836 45728
rect 32772 45668 32776 45724
rect 32776 45668 32832 45724
rect 32832 45668 32836 45724
rect 32772 45664 32836 45668
rect 32852 45724 32916 45728
rect 32852 45668 32856 45724
rect 32856 45668 32912 45724
rect 32912 45668 32916 45724
rect 32852 45664 32916 45668
rect 37612 45724 37676 45728
rect 37612 45668 37616 45724
rect 37616 45668 37672 45724
rect 37672 45668 37676 45724
rect 37612 45664 37676 45668
rect 37692 45724 37756 45728
rect 37692 45668 37696 45724
rect 37696 45668 37752 45724
rect 37752 45668 37756 45724
rect 37692 45664 37756 45668
rect 37772 45724 37836 45728
rect 37772 45668 37776 45724
rect 37776 45668 37832 45724
rect 37832 45668 37836 45724
rect 37772 45664 37836 45668
rect 37852 45724 37916 45728
rect 37852 45668 37856 45724
rect 37856 45668 37912 45724
rect 37912 45668 37916 45724
rect 37852 45664 37916 45668
rect 1952 45180 2016 45184
rect 1952 45124 1956 45180
rect 1956 45124 2012 45180
rect 2012 45124 2016 45180
rect 1952 45120 2016 45124
rect 2032 45180 2096 45184
rect 2032 45124 2036 45180
rect 2036 45124 2092 45180
rect 2092 45124 2096 45180
rect 2032 45120 2096 45124
rect 2112 45180 2176 45184
rect 2112 45124 2116 45180
rect 2116 45124 2172 45180
rect 2172 45124 2176 45180
rect 2112 45120 2176 45124
rect 2192 45180 2256 45184
rect 2192 45124 2196 45180
rect 2196 45124 2252 45180
rect 2252 45124 2256 45180
rect 2192 45120 2256 45124
rect 6952 45180 7016 45184
rect 6952 45124 6956 45180
rect 6956 45124 7012 45180
rect 7012 45124 7016 45180
rect 6952 45120 7016 45124
rect 7032 45180 7096 45184
rect 7032 45124 7036 45180
rect 7036 45124 7092 45180
rect 7092 45124 7096 45180
rect 7032 45120 7096 45124
rect 7112 45180 7176 45184
rect 7112 45124 7116 45180
rect 7116 45124 7172 45180
rect 7172 45124 7176 45180
rect 7112 45120 7176 45124
rect 7192 45180 7256 45184
rect 7192 45124 7196 45180
rect 7196 45124 7252 45180
rect 7252 45124 7256 45180
rect 7192 45120 7256 45124
rect 11952 45180 12016 45184
rect 11952 45124 11956 45180
rect 11956 45124 12012 45180
rect 12012 45124 12016 45180
rect 11952 45120 12016 45124
rect 12032 45180 12096 45184
rect 12032 45124 12036 45180
rect 12036 45124 12092 45180
rect 12092 45124 12096 45180
rect 12032 45120 12096 45124
rect 12112 45180 12176 45184
rect 12112 45124 12116 45180
rect 12116 45124 12172 45180
rect 12172 45124 12176 45180
rect 12112 45120 12176 45124
rect 12192 45180 12256 45184
rect 12192 45124 12196 45180
rect 12196 45124 12252 45180
rect 12252 45124 12256 45180
rect 12192 45120 12256 45124
rect 16952 45180 17016 45184
rect 16952 45124 16956 45180
rect 16956 45124 17012 45180
rect 17012 45124 17016 45180
rect 16952 45120 17016 45124
rect 17032 45180 17096 45184
rect 17032 45124 17036 45180
rect 17036 45124 17092 45180
rect 17092 45124 17096 45180
rect 17032 45120 17096 45124
rect 17112 45180 17176 45184
rect 17112 45124 17116 45180
rect 17116 45124 17172 45180
rect 17172 45124 17176 45180
rect 17112 45120 17176 45124
rect 17192 45180 17256 45184
rect 17192 45124 17196 45180
rect 17196 45124 17252 45180
rect 17252 45124 17256 45180
rect 17192 45120 17256 45124
rect 21952 45180 22016 45184
rect 21952 45124 21956 45180
rect 21956 45124 22012 45180
rect 22012 45124 22016 45180
rect 21952 45120 22016 45124
rect 22032 45180 22096 45184
rect 22032 45124 22036 45180
rect 22036 45124 22092 45180
rect 22092 45124 22096 45180
rect 22032 45120 22096 45124
rect 22112 45180 22176 45184
rect 22112 45124 22116 45180
rect 22116 45124 22172 45180
rect 22172 45124 22176 45180
rect 22112 45120 22176 45124
rect 22192 45180 22256 45184
rect 22192 45124 22196 45180
rect 22196 45124 22252 45180
rect 22252 45124 22256 45180
rect 22192 45120 22256 45124
rect 26952 45180 27016 45184
rect 26952 45124 26956 45180
rect 26956 45124 27012 45180
rect 27012 45124 27016 45180
rect 26952 45120 27016 45124
rect 27032 45180 27096 45184
rect 27032 45124 27036 45180
rect 27036 45124 27092 45180
rect 27092 45124 27096 45180
rect 27032 45120 27096 45124
rect 27112 45180 27176 45184
rect 27112 45124 27116 45180
rect 27116 45124 27172 45180
rect 27172 45124 27176 45180
rect 27112 45120 27176 45124
rect 27192 45180 27256 45184
rect 27192 45124 27196 45180
rect 27196 45124 27252 45180
rect 27252 45124 27256 45180
rect 27192 45120 27256 45124
rect 31952 45180 32016 45184
rect 31952 45124 31956 45180
rect 31956 45124 32012 45180
rect 32012 45124 32016 45180
rect 31952 45120 32016 45124
rect 32032 45180 32096 45184
rect 32032 45124 32036 45180
rect 32036 45124 32092 45180
rect 32092 45124 32096 45180
rect 32032 45120 32096 45124
rect 32112 45180 32176 45184
rect 32112 45124 32116 45180
rect 32116 45124 32172 45180
rect 32172 45124 32176 45180
rect 32112 45120 32176 45124
rect 32192 45180 32256 45184
rect 32192 45124 32196 45180
rect 32196 45124 32252 45180
rect 32252 45124 32256 45180
rect 32192 45120 32256 45124
rect 36952 45180 37016 45184
rect 36952 45124 36956 45180
rect 36956 45124 37012 45180
rect 37012 45124 37016 45180
rect 36952 45120 37016 45124
rect 37032 45180 37096 45184
rect 37032 45124 37036 45180
rect 37036 45124 37092 45180
rect 37092 45124 37096 45180
rect 37032 45120 37096 45124
rect 37112 45180 37176 45184
rect 37112 45124 37116 45180
rect 37116 45124 37172 45180
rect 37172 45124 37176 45180
rect 37112 45120 37176 45124
rect 37192 45180 37256 45184
rect 37192 45124 37196 45180
rect 37196 45124 37252 45180
rect 37252 45124 37256 45180
rect 37192 45120 37256 45124
rect 2612 44636 2676 44640
rect 2612 44580 2616 44636
rect 2616 44580 2672 44636
rect 2672 44580 2676 44636
rect 2612 44576 2676 44580
rect 2692 44636 2756 44640
rect 2692 44580 2696 44636
rect 2696 44580 2752 44636
rect 2752 44580 2756 44636
rect 2692 44576 2756 44580
rect 2772 44636 2836 44640
rect 2772 44580 2776 44636
rect 2776 44580 2832 44636
rect 2832 44580 2836 44636
rect 2772 44576 2836 44580
rect 2852 44636 2916 44640
rect 2852 44580 2856 44636
rect 2856 44580 2912 44636
rect 2912 44580 2916 44636
rect 2852 44576 2916 44580
rect 7612 44636 7676 44640
rect 7612 44580 7616 44636
rect 7616 44580 7672 44636
rect 7672 44580 7676 44636
rect 7612 44576 7676 44580
rect 7692 44636 7756 44640
rect 7692 44580 7696 44636
rect 7696 44580 7752 44636
rect 7752 44580 7756 44636
rect 7692 44576 7756 44580
rect 7772 44636 7836 44640
rect 7772 44580 7776 44636
rect 7776 44580 7832 44636
rect 7832 44580 7836 44636
rect 7772 44576 7836 44580
rect 7852 44636 7916 44640
rect 7852 44580 7856 44636
rect 7856 44580 7912 44636
rect 7912 44580 7916 44636
rect 7852 44576 7916 44580
rect 12612 44636 12676 44640
rect 12612 44580 12616 44636
rect 12616 44580 12672 44636
rect 12672 44580 12676 44636
rect 12612 44576 12676 44580
rect 12692 44636 12756 44640
rect 12692 44580 12696 44636
rect 12696 44580 12752 44636
rect 12752 44580 12756 44636
rect 12692 44576 12756 44580
rect 12772 44636 12836 44640
rect 12772 44580 12776 44636
rect 12776 44580 12832 44636
rect 12832 44580 12836 44636
rect 12772 44576 12836 44580
rect 12852 44636 12916 44640
rect 12852 44580 12856 44636
rect 12856 44580 12912 44636
rect 12912 44580 12916 44636
rect 12852 44576 12916 44580
rect 17612 44636 17676 44640
rect 17612 44580 17616 44636
rect 17616 44580 17672 44636
rect 17672 44580 17676 44636
rect 17612 44576 17676 44580
rect 17692 44636 17756 44640
rect 17692 44580 17696 44636
rect 17696 44580 17752 44636
rect 17752 44580 17756 44636
rect 17692 44576 17756 44580
rect 17772 44636 17836 44640
rect 17772 44580 17776 44636
rect 17776 44580 17832 44636
rect 17832 44580 17836 44636
rect 17772 44576 17836 44580
rect 17852 44636 17916 44640
rect 17852 44580 17856 44636
rect 17856 44580 17912 44636
rect 17912 44580 17916 44636
rect 17852 44576 17916 44580
rect 22612 44636 22676 44640
rect 22612 44580 22616 44636
rect 22616 44580 22672 44636
rect 22672 44580 22676 44636
rect 22612 44576 22676 44580
rect 22692 44636 22756 44640
rect 22692 44580 22696 44636
rect 22696 44580 22752 44636
rect 22752 44580 22756 44636
rect 22692 44576 22756 44580
rect 22772 44636 22836 44640
rect 22772 44580 22776 44636
rect 22776 44580 22832 44636
rect 22832 44580 22836 44636
rect 22772 44576 22836 44580
rect 22852 44636 22916 44640
rect 22852 44580 22856 44636
rect 22856 44580 22912 44636
rect 22912 44580 22916 44636
rect 22852 44576 22916 44580
rect 27612 44636 27676 44640
rect 27612 44580 27616 44636
rect 27616 44580 27672 44636
rect 27672 44580 27676 44636
rect 27612 44576 27676 44580
rect 27692 44636 27756 44640
rect 27692 44580 27696 44636
rect 27696 44580 27752 44636
rect 27752 44580 27756 44636
rect 27692 44576 27756 44580
rect 27772 44636 27836 44640
rect 27772 44580 27776 44636
rect 27776 44580 27832 44636
rect 27832 44580 27836 44636
rect 27772 44576 27836 44580
rect 27852 44636 27916 44640
rect 27852 44580 27856 44636
rect 27856 44580 27912 44636
rect 27912 44580 27916 44636
rect 27852 44576 27916 44580
rect 32612 44636 32676 44640
rect 32612 44580 32616 44636
rect 32616 44580 32672 44636
rect 32672 44580 32676 44636
rect 32612 44576 32676 44580
rect 32692 44636 32756 44640
rect 32692 44580 32696 44636
rect 32696 44580 32752 44636
rect 32752 44580 32756 44636
rect 32692 44576 32756 44580
rect 32772 44636 32836 44640
rect 32772 44580 32776 44636
rect 32776 44580 32832 44636
rect 32832 44580 32836 44636
rect 32772 44576 32836 44580
rect 32852 44636 32916 44640
rect 32852 44580 32856 44636
rect 32856 44580 32912 44636
rect 32912 44580 32916 44636
rect 32852 44576 32916 44580
rect 37612 44636 37676 44640
rect 37612 44580 37616 44636
rect 37616 44580 37672 44636
rect 37672 44580 37676 44636
rect 37612 44576 37676 44580
rect 37692 44636 37756 44640
rect 37692 44580 37696 44636
rect 37696 44580 37752 44636
rect 37752 44580 37756 44636
rect 37692 44576 37756 44580
rect 37772 44636 37836 44640
rect 37772 44580 37776 44636
rect 37776 44580 37832 44636
rect 37832 44580 37836 44636
rect 37772 44576 37836 44580
rect 37852 44636 37916 44640
rect 37852 44580 37856 44636
rect 37856 44580 37912 44636
rect 37912 44580 37916 44636
rect 37852 44576 37916 44580
rect 1952 44092 2016 44096
rect 1952 44036 1956 44092
rect 1956 44036 2012 44092
rect 2012 44036 2016 44092
rect 1952 44032 2016 44036
rect 2032 44092 2096 44096
rect 2032 44036 2036 44092
rect 2036 44036 2092 44092
rect 2092 44036 2096 44092
rect 2032 44032 2096 44036
rect 2112 44092 2176 44096
rect 2112 44036 2116 44092
rect 2116 44036 2172 44092
rect 2172 44036 2176 44092
rect 2112 44032 2176 44036
rect 2192 44092 2256 44096
rect 2192 44036 2196 44092
rect 2196 44036 2252 44092
rect 2252 44036 2256 44092
rect 2192 44032 2256 44036
rect 6952 44092 7016 44096
rect 6952 44036 6956 44092
rect 6956 44036 7012 44092
rect 7012 44036 7016 44092
rect 6952 44032 7016 44036
rect 7032 44092 7096 44096
rect 7032 44036 7036 44092
rect 7036 44036 7092 44092
rect 7092 44036 7096 44092
rect 7032 44032 7096 44036
rect 7112 44092 7176 44096
rect 7112 44036 7116 44092
rect 7116 44036 7172 44092
rect 7172 44036 7176 44092
rect 7112 44032 7176 44036
rect 7192 44092 7256 44096
rect 7192 44036 7196 44092
rect 7196 44036 7252 44092
rect 7252 44036 7256 44092
rect 7192 44032 7256 44036
rect 11952 44092 12016 44096
rect 11952 44036 11956 44092
rect 11956 44036 12012 44092
rect 12012 44036 12016 44092
rect 11952 44032 12016 44036
rect 12032 44092 12096 44096
rect 12032 44036 12036 44092
rect 12036 44036 12092 44092
rect 12092 44036 12096 44092
rect 12032 44032 12096 44036
rect 12112 44092 12176 44096
rect 12112 44036 12116 44092
rect 12116 44036 12172 44092
rect 12172 44036 12176 44092
rect 12112 44032 12176 44036
rect 12192 44092 12256 44096
rect 12192 44036 12196 44092
rect 12196 44036 12252 44092
rect 12252 44036 12256 44092
rect 12192 44032 12256 44036
rect 16952 44092 17016 44096
rect 16952 44036 16956 44092
rect 16956 44036 17012 44092
rect 17012 44036 17016 44092
rect 16952 44032 17016 44036
rect 17032 44092 17096 44096
rect 17032 44036 17036 44092
rect 17036 44036 17092 44092
rect 17092 44036 17096 44092
rect 17032 44032 17096 44036
rect 17112 44092 17176 44096
rect 17112 44036 17116 44092
rect 17116 44036 17172 44092
rect 17172 44036 17176 44092
rect 17112 44032 17176 44036
rect 17192 44092 17256 44096
rect 17192 44036 17196 44092
rect 17196 44036 17252 44092
rect 17252 44036 17256 44092
rect 17192 44032 17256 44036
rect 21952 44092 22016 44096
rect 21952 44036 21956 44092
rect 21956 44036 22012 44092
rect 22012 44036 22016 44092
rect 21952 44032 22016 44036
rect 22032 44092 22096 44096
rect 22032 44036 22036 44092
rect 22036 44036 22092 44092
rect 22092 44036 22096 44092
rect 22032 44032 22096 44036
rect 22112 44092 22176 44096
rect 22112 44036 22116 44092
rect 22116 44036 22172 44092
rect 22172 44036 22176 44092
rect 22112 44032 22176 44036
rect 22192 44092 22256 44096
rect 22192 44036 22196 44092
rect 22196 44036 22252 44092
rect 22252 44036 22256 44092
rect 22192 44032 22256 44036
rect 26952 44092 27016 44096
rect 26952 44036 26956 44092
rect 26956 44036 27012 44092
rect 27012 44036 27016 44092
rect 26952 44032 27016 44036
rect 27032 44092 27096 44096
rect 27032 44036 27036 44092
rect 27036 44036 27092 44092
rect 27092 44036 27096 44092
rect 27032 44032 27096 44036
rect 27112 44092 27176 44096
rect 27112 44036 27116 44092
rect 27116 44036 27172 44092
rect 27172 44036 27176 44092
rect 27112 44032 27176 44036
rect 27192 44092 27256 44096
rect 27192 44036 27196 44092
rect 27196 44036 27252 44092
rect 27252 44036 27256 44092
rect 27192 44032 27256 44036
rect 31952 44092 32016 44096
rect 31952 44036 31956 44092
rect 31956 44036 32012 44092
rect 32012 44036 32016 44092
rect 31952 44032 32016 44036
rect 32032 44092 32096 44096
rect 32032 44036 32036 44092
rect 32036 44036 32092 44092
rect 32092 44036 32096 44092
rect 32032 44032 32096 44036
rect 32112 44092 32176 44096
rect 32112 44036 32116 44092
rect 32116 44036 32172 44092
rect 32172 44036 32176 44092
rect 32112 44032 32176 44036
rect 32192 44092 32256 44096
rect 32192 44036 32196 44092
rect 32196 44036 32252 44092
rect 32252 44036 32256 44092
rect 32192 44032 32256 44036
rect 36952 44092 37016 44096
rect 36952 44036 36956 44092
rect 36956 44036 37012 44092
rect 37012 44036 37016 44092
rect 36952 44032 37016 44036
rect 37032 44092 37096 44096
rect 37032 44036 37036 44092
rect 37036 44036 37092 44092
rect 37092 44036 37096 44092
rect 37032 44032 37096 44036
rect 37112 44092 37176 44096
rect 37112 44036 37116 44092
rect 37116 44036 37172 44092
rect 37172 44036 37176 44092
rect 37112 44032 37176 44036
rect 37192 44092 37256 44096
rect 37192 44036 37196 44092
rect 37196 44036 37252 44092
rect 37252 44036 37256 44092
rect 37192 44032 37256 44036
rect 2612 43548 2676 43552
rect 2612 43492 2616 43548
rect 2616 43492 2672 43548
rect 2672 43492 2676 43548
rect 2612 43488 2676 43492
rect 2692 43548 2756 43552
rect 2692 43492 2696 43548
rect 2696 43492 2752 43548
rect 2752 43492 2756 43548
rect 2692 43488 2756 43492
rect 2772 43548 2836 43552
rect 2772 43492 2776 43548
rect 2776 43492 2832 43548
rect 2832 43492 2836 43548
rect 2772 43488 2836 43492
rect 2852 43548 2916 43552
rect 2852 43492 2856 43548
rect 2856 43492 2912 43548
rect 2912 43492 2916 43548
rect 2852 43488 2916 43492
rect 7612 43548 7676 43552
rect 7612 43492 7616 43548
rect 7616 43492 7672 43548
rect 7672 43492 7676 43548
rect 7612 43488 7676 43492
rect 7692 43548 7756 43552
rect 7692 43492 7696 43548
rect 7696 43492 7752 43548
rect 7752 43492 7756 43548
rect 7692 43488 7756 43492
rect 7772 43548 7836 43552
rect 7772 43492 7776 43548
rect 7776 43492 7832 43548
rect 7832 43492 7836 43548
rect 7772 43488 7836 43492
rect 7852 43548 7916 43552
rect 7852 43492 7856 43548
rect 7856 43492 7912 43548
rect 7912 43492 7916 43548
rect 7852 43488 7916 43492
rect 12612 43548 12676 43552
rect 12612 43492 12616 43548
rect 12616 43492 12672 43548
rect 12672 43492 12676 43548
rect 12612 43488 12676 43492
rect 12692 43548 12756 43552
rect 12692 43492 12696 43548
rect 12696 43492 12752 43548
rect 12752 43492 12756 43548
rect 12692 43488 12756 43492
rect 12772 43548 12836 43552
rect 12772 43492 12776 43548
rect 12776 43492 12832 43548
rect 12832 43492 12836 43548
rect 12772 43488 12836 43492
rect 12852 43548 12916 43552
rect 12852 43492 12856 43548
rect 12856 43492 12912 43548
rect 12912 43492 12916 43548
rect 12852 43488 12916 43492
rect 17612 43548 17676 43552
rect 17612 43492 17616 43548
rect 17616 43492 17672 43548
rect 17672 43492 17676 43548
rect 17612 43488 17676 43492
rect 17692 43548 17756 43552
rect 17692 43492 17696 43548
rect 17696 43492 17752 43548
rect 17752 43492 17756 43548
rect 17692 43488 17756 43492
rect 17772 43548 17836 43552
rect 17772 43492 17776 43548
rect 17776 43492 17832 43548
rect 17832 43492 17836 43548
rect 17772 43488 17836 43492
rect 17852 43548 17916 43552
rect 17852 43492 17856 43548
rect 17856 43492 17912 43548
rect 17912 43492 17916 43548
rect 17852 43488 17916 43492
rect 22612 43548 22676 43552
rect 22612 43492 22616 43548
rect 22616 43492 22672 43548
rect 22672 43492 22676 43548
rect 22612 43488 22676 43492
rect 22692 43548 22756 43552
rect 22692 43492 22696 43548
rect 22696 43492 22752 43548
rect 22752 43492 22756 43548
rect 22692 43488 22756 43492
rect 22772 43548 22836 43552
rect 22772 43492 22776 43548
rect 22776 43492 22832 43548
rect 22832 43492 22836 43548
rect 22772 43488 22836 43492
rect 22852 43548 22916 43552
rect 22852 43492 22856 43548
rect 22856 43492 22912 43548
rect 22912 43492 22916 43548
rect 22852 43488 22916 43492
rect 27612 43548 27676 43552
rect 27612 43492 27616 43548
rect 27616 43492 27672 43548
rect 27672 43492 27676 43548
rect 27612 43488 27676 43492
rect 27692 43548 27756 43552
rect 27692 43492 27696 43548
rect 27696 43492 27752 43548
rect 27752 43492 27756 43548
rect 27692 43488 27756 43492
rect 27772 43548 27836 43552
rect 27772 43492 27776 43548
rect 27776 43492 27832 43548
rect 27832 43492 27836 43548
rect 27772 43488 27836 43492
rect 27852 43548 27916 43552
rect 27852 43492 27856 43548
rect 27856 43492 27912 43548
rect 27912 43492 27916 43548
rect 27852 43488 27916 43492
rect 32612 43548 32676 43552
rect 32612 43492 32616 43548
rect 32616 43492 32672 43548
rect 32672 43492 32676 43548
rect 32612 43488 32676 43492
rect 32692 43548 32756 43552
rect 32692 43492 32696 43548
rect 32696 43492 32752 43548
rect 32752 43492 32756 43548
rect 32692 43488 32756 43492
rect 32772 43548 32836 43552
rect 32772 43492 32776 43548
rect 32776 43492 32832 43548
rect 32832 43492 32836 43548
rect 32772 43488 32836 43492
rect 32852 43548 32916 43552
rect 32852 43492 32856 43548
rect 32856 43492 32912 43548
rect 32912 43492 32916 43548
rect 32852 43488 32916 43492
rect 37612 43548 37676 43552
rect 37612 43492 37616 43548
rect 37616 43492 37672 43548
rect 37672 43492 37676 43548
rect 37612 43488 37676 43492
rect 37692 43548 37756 43552
rect 37692 43492 37696 43548
rect 37696 43492 37752 43548
rect 37752 43492 37756 43548
rect 37692 43488 37756 43492
rect 37772 43548 37836 43552
rect 37772 43492 37776 43548
rect 37776 43492 37832 43548
rect 37832 43492 37836 43548
rect 37772 43488 37836 43492
rect 37852 43548 37916 43552
rect 37852 43492 37856 43548
rect 37856 43492 37912 43548
rect 37912 43492 37916 43548
rect 37852 43488 37916 43492
rect 1952 43004 2016 43008
rect 1952 42948 1956 43004
rect 1956 42948 2012 43004
rect 2012 42948 2016 43004
rect 1952 42944 2016 42948
rect 2032 43004 2096 43008
rect 2032 42948 2036 43004
rect 2036 42948 2092 43004
rect 2092 42948 2096 43004
rect 2032 42944 2096 42948
rect 2112 43004 2176 43008
rect 2112 42948 2116 43004
rect 2116 42948 2172 43004
rect 2172 42948 2176 43004
rect 2112 42944 2176 42948
rect 2192 43004 2256 43008
rect 2192 42948 2196 43004
rect 2196 42948 2252 43004
rect 2252 42948 2256 43004
rect 2192 42944 2256 42948
rect 6952 43004 7016 43008
rect 6952 42948 6956 43004
rect 6956 42948 7012 43004
rect 7012 42948 7016 43004
rect 6952 42944 7016 42948
rect 7032 43004 7096 43008
rect 7032 42948 7036 43004
rect 7036 42948 7092 43004
rect 7092 42948 7096 43004
rect 7032 42944 7096 42948
rect 7112 43004 7176 43008
rect 7112 42948 7116 43004
rect 7116 42948 7172 43004
rect 7172 42948 7176 43004
rect 7112 42944 7176 42948
rect 7192 43004 7256 43008
rect 7192 42948 7196 43004
rect 7196 42948 7252 43004
rect 7252 42948 7256 43004
rect 7192 42944 7256 42948
rect 11952 43004 12016 43008
rect 11952 42948 11956 43004
rect 11956 42948 12012 43004
rect 12012 42948 12016 43004
rect 11952 42944 12016 42948
rect 12032 43004 12096 43008
rect 12032 42948 12036 43004
rect 12036 42948 12092 43004
rect 12092 42948 12096 43004
rect 12032 42944 12096 42948
rect 12112 43004 12176 43008
rect 12112 42948 12116 43004
rect 12116 42948 12172 43004
rect 12172 42948 12176 43004
rect 12112 42944 12176 42948
rect 12192 43004 12256 43008
rect 12192 42948 12196 43004
rect 12196 42948 12252 43004
rect 12252 42948 12256 43004
rect 12192 42944 12256 42948
rect 16952 43004 17016 43008
rect 16952 42948 16956 43004
rect 16956 42948 17012 43004
rect 17012 42948 17016 43004
rect 16952 42944 17016 42948
rect 17032 43004 17096 43008
rect 17032 42948 17036 43004
rect 17036 42948 17092 43004
rect 17092 42948 17096 43004
rect 17032 42944 17096 42948
rect 17112 43004 17176 43008
rect 17112 42948 17116 43004
rect 17116 42948 17172 43004
rect 17172 42948 17176 43004
rect 17112 42944 17176 42948
rect 17192 43004 17256 43008
rect 17192 42948 17196 43004
rect 17196 42948 17252 43004
rect 17252 42948 17256 43004
rect 17192 42944 17256 42948
rect 21952 43004 22016 43008
rect 21952 42948 21956 43004
rect 21956 42948 22012 43004
rect 22012 42948 22016 43004
rect 21952 42944 22016 42948
rect 22032 43004 22096 43008
rect 22032 42948 22036 43004
rect 22036 42948 22092 43004
rect 22092 42948 22096 43004
rect 22032 42944 22096 42948
rect 22112 43004 22176 43008
rect 22112 42948 22116 43004
rect 22116 42948 22172 43004
rect 22172 42948 22176 43004
rect 22112 42944 22176 42948
rect 22192 43004 22256 43008
rect 22192 42948 22196 43004
rect 22196 42948 22252 43004
rect 22252 42948 22256 43004
rect 22192 42944 22256 42948
rect 26952 43004 27016 43008
rect 26952 42948 26956 43004
rect 26956 42948 27012 43004
rect 27012 42948 27016 43004
rect 26952 42944 27016 42948
rect 27032 43004 27096 43008
rect 27032 42948 27036 43004
rect 27036 42948 27092 43004
rect 27092 42948 27096 43004
rect 27032 42944 27096 42948
rect 27112 43004 27176 43008
rect 27112 42948 27116 43004
rect 27116 42948 27172 43004
rect 27172 42948 27176 43004
rect 27112 42944 27176 42948
rect 27192 43004 27256 43008
rect 27192 42948 27196 43004
rect 27196 42948 27252 43004
rect 27252 42948 27256 43004
rect 27192 42944 27256 42948
rect 31952 43004 32016 43008
rect 31952 42948 31956 43004
rect 31956 42948 32012 43004
rect 32012 42948 32016 43004
rect 31952 42944 32016 42948
rect 32032 43004 32096 43008
rect 32032 42948 32036 43004
rect 32036 42948 32092 43004
rect 32092 42948 32096 43004
rect 32032 42944 32096 42948
rect 32112 43004 32176 43008
rect 32112 42948 32116 43004
rect 32116 42948 32172 43004
rect 32172 42948 32176 43004
rect 32112 42944 32176 42948
rect 32192 43004 32256 43008
rect 32192 42948 32196 43004
rect 32196 42948 32252 43004
rect 32252 42948 32256 43004
rect 32192 42944 32256 42948
rect 36952 43004 37016 43008
rect 36952 42948 36956 43004
rect 36956 42948 37012 43004
rect 37012 42948 37016 43004
rect 36952 42944 37016 42948
rect 37032 43004 37096 43008
rect 37032 42948 37036 43004
rect 37036 42948 37092 43004
rect 37092 42948 37096 43004
rect 37032 42944 37096 42948
rect 37112 43004 37176 43008
rect 37112 42948 37116 43004
rect 37116 42948 37172 43004
rect 37172 42948 37176 43004
rect 37112 42944 37176 42948
rect 37192 43004 37256 43008
rect 37192 42948 37196 43004
rect 37196 42948 37252 43004
rect 37252 42948 37256 43004
rect 37192 42944 37256 42948
rect 2612 42460 2676 42464
rect 2612 42404 2616 42460
rect 2616 42404 2672 42460
rect 2672 42404 2676 42460
rect 2612 42400 2676 42404
rect 2692 42460 2756 42464
rect 2692 42404 2696 42460
rect 2696 42404 2752 42460
rect 2752 42404 2756 42460
rect 2692 42400 2756 42404
rect 2772 42460 2836 42464
rect 2772 42404 2776 42460
rect 2776 42404 2832 42460
rect 2832 42404 2836 42460
rect 2772 42400 2836 42404
rect 2852 42460 2916 42464
rect 2852 42404 2856 42460
rect 2856 42404 2912 42460
rect 2912 42404 2916 42460
rect 2852 42400 2916 42404
rect 7612 42460 7676 42464
rect 7612 42404 7616 42460
rect 7616 42404 7672 42460
rect 7672 42404 7676 42460
rect 7612 42400 7676 42404
rect 7692 42460 7756 42464
rect 7692 42404 7696 42460
rect 7696 42404 7752 42460
rect 7752 42404 7756 42460
rect 7692 42400 7756 42404
rect 7772 42460 7836 42464
rect 7772 42404 7776 42460
rect 7776 42404 7832 42460
rect 7832 42404 7836 42460
rect 7772 42400 7836 42404
rect 7852 42460 7916 42464
rect 7852 42404 7856 42460
rect 7856 42404 7912 42460
rect 7912 42404 7916 42460
rect 7852 42400 7916 42404
rect 12612 42460 12676 42464
rect 12612 42404 12616 42460
rect 12616 42404 12672 42460
rect 12672 42404 12676 42460
rect 12612 42400 12676 42404
rect 12692 42460 12756 42464
rect 12692 42404 12696 42460
rect 12696 42404 12752 42460
rect 12752 42404 12756 42460
rect 12692 42400 12756 42404
rect 12772 42460 12836 42464
rect 12772 42404 12776 42460
rect 12776 42404 12832 42460
rect 12832 42404 12836 42460
rect 12772 42400 12836 42404
rect 12852 42460 12916 42464
rect 12852 42404 12856 42460
rect 12856 42404 12912 42460
rect 12912 42404 12916 42460
rect 12852 42400 12916 42404
rect 17612 42460 17676 42464
rect 17612 42404 17616 42460
rect 17616 42404 17672 42460
rect 17672 42404 17676 42460
rect 17612 42400 17676 42404
rect 17692 42460 17756 42464
rect 17692 42404 17696 42460
rect 17696 42404 17752 42460
rect 17752 42404 17756 42460
rect 17692 42400 17756 42404
rect 17772 42460 17836 42464
rect 17772 42404 17776 42460
rect 17776 42404 17832 42460
rect 17832 42404 17836 42460
rect 17772 42400 17836 42404
rect 17852 42460 17916 42464
rect 17852 42404 17856 42460
rect 17856 42404 17912 42460
rect 17912 42404 17916 42460
rect 17852 42400 17916 42404
rect 22612 42460 22676 42464
rect 22612 42404 22616 42460
rect 22616 42404 22672 42460
rect 22672 42404 22676 42460
rect 22612 42400 22676 42404
rect 22692 42460 22756 42464
rect 22692 42404 22696 42460
rect 22696 42404 22752 42460
rect 22752 42404 22756 42460
rect 22692 42400 22756 42404
rect 22772 42460 22836 42464
rect 22772 42404 22776 42460
rect 22776 42404 22832 42460
rect 22832 42404 22836 42460
rect 22772 42400 22836 42404
rect 22852 42460 22916 42464
rect 22852 42404 22856 42460
rect 22856 42404 22912 42460
rect 22912 42404 22916 42460
rect 22852 42400 22916 42404
rect 27612 42460 27676 42464
rect 27612 42404 27616 42460
rect 27616 42404 27672 42460
rect 27672 42404 27676 42460
rect 27612 42400 27676 42404
rect 27692 42460 27756 42464
rect 27692 42404 27696 42460
rect 27696 42404 27752 42460
rect 27752 42404 27756 42460
rect 27692 42400 27756 42404
rect 27772 42460 27836 42464
rect 27772 42404 27776 42460
rect 27776 42404 27832 42460
rect 27832 42404 27836 42460
rect 27772 42400 27836 42404
rect 27852 42460 27916 42464
rect 27852 42404 27856 42460
rect 27856 42404 27912 42460
rect 27912 42404 27916 42460
rect 27852 42400 27916 42404
rect 32612 42460 32676 42464
rect 32612 42404 32616 42460
rect 32616 42404 32672 42460
rect 32672 42404 32676 42460
rect 32612 42400 32676 42404
rect 32692 42460 32756 42464
rect 32692 42404 32696 42460
rect 32696 42404 32752 42460
rect 32752 42404 32756 42460
rect 32692 42400 32756 42404
rect 32772 42460 32836 42464
rect 32772 42404 32776 42460
rect 32776 42404 32832 42460
rect 32832 42404 32836 42460
rect 32772 42400 32836 42404
rect 32852 42460 32916 42464
rect 32852 42404 32856 42460
rect 32856 42404 32912 42460
rect 32912 42404 32916 42460
rect 32852 42400 32916 42404
rect 37612 42460 37676 42464
rect 37612 42404 37616 42460
rect 37616 42404 37672 42460
rect 37672 42404 37676 42460
rect 37612 42400 37676 42404
rect 37692 42460 37756 42464
rect 37692 42404 37696 42460
rect 37696 42404 37752 42460
rect 37752 42404 37756 42460
rect 37692 42400 37756 42404
rect 37772 42460 37836 42464
rect 37772 42404 37776 42460
rect 37776 42404 37832 42460
rect 37832 42404 37836 42460
rect 37772 42400 37836 42404
rect 37852 42460 37916 42464
rect 37852 42404 37856 42460
rect 37856 42404 37912 42460
rect 37912 42404 37916 42460
rect 37852 42400 37916 42404
rect 1952 41916 2016 41920
rect 1952 41860 1956 41916
rect 1956 41860 2012 41916
rect 2012 41860 2016 41916
rect 1952 41856 2016 41860
rect 2032 41916 2096 41920
rect 2032 41860 2036 41916
rect 2036 41860 2092 41916
rect 2092 41860 2096 41916
rect 2032 41856 2096 41860
rect 2112 41916 2176 41920
rect 2112 41860 2116 41916
rect 2116 41860 2172 41916
rect 2172 41860 2176 41916
rect 2112 41856 2176 41860
rect 2192 41916 2256 41920
rect 2192 41860 2196 41916
rect 2196 41860 2252 41916
rect 2252 41860 2256 41916
rect 2192 41856 2256 41860
rect 6952 41916 7016 41920
rect 6952 41860 6956 41916
rect 6956 41860 7012 41916
rect 7012 41860 7016 41916
rect 6952 41856 7016 41860
rect 7032 41916 7096 41920
rect 7032 41860 7036 41916
rect 7036 41860 7092 41916
rect 7092 41860 7096 41916
rect 7032 41856 7096 41860
rect 7112 41916 7176 41920
rect 7112 41860 7116 41916
rect 7116 41860 7172 41916
rect 7172 41860 7176 41916
rect 7112 41856 7176 41860
rect 7192 41916 7256 41920
rect 7192 41860 7196 41916
rect 7196 41860 7252 41916
rect 7252 41860 7256 41916
rect 7192 41856 7256 41860
rect 11952 41916 12016 41920
rect 11952 41860 11956 41916
rect 11956 41860 12012 41916
rect 12012 41860 12016 41916
rect 11952 41856 12016 41860
rect 12032 41916 12096 41920
rect 12032 41860 12036 41916
rect 12036 41860 12092 41916
rect 12092 41860 12096 41916
rect 12032 41856 12096 41860
rect 12112 41916 12176 41920
rect 12112 41860 12116 41916
rect 12116 41860 12172 41916
rect 12172 41860 12176 41916
rect 12112 41856 12176 41860
rect 12192 41916 12256 41920
rect 12192 41860 12196 41916
rect 12196 41860 12252 41916
rect 12252 41860 12256 41916
rect 12192 41856 12256 41860
rect 16952 41916 17016 41920
rect 16952 41860 16956 41916
rect 16956 41860 17012 41916
rect 17012 41860 17016 41916
rect 16952 41856 17016 41860
rect 17032 41916 17096 41920
rect 17032 41860 17036 41916
rect 17036 41860 17092 41916
rect 17092 41860 17096 41916
rect 17032 41856 17096 41860
rect 17112 41916 17176 41920
rect 17112 41860 17116 41916
rect 17116 41860 17172 41916
rect 17172 41860 17176 41916
rect 17112 41856 17176 41860
rect 17192 41916 17256 41920
rect 17192 41860 17196 41916
rect 17196 41860 17252 41916
rect 17252 41860 17256 41916
rect 17192 41856 17256 41860
rect 21952 41916 22016 41920
rect 21952 41860 21956 41916
rect 21956 41860 22012 41916
rect 22012 41860 22016 41916
rect 21952 41856 22016 41860
rect 22032 41916 22096 41920
rect 22032 41860 22036 41916
rect 22036 41860 22092 41916
rect 22092 41860 22096 41916
rect 22032 41856 22096 41860
rect 22112 41916 22176 41920
rect 22112 41860 22116 41916
rect 22116 41860 22172 41916
rect 22172 41860 22176 41916
rect 22112 41856 22176 41860
rect 22192 41916 22256 41920
rect 22192 41860 22196 41916
rect 22196 41860 22252 41916
rect 22252 41860 22256 41916
rect 22192 41856 22256 41860
rect 26952 41916 27016 41920
rect 26952 41860 26956 41916
rect 26956 41860 27012 41916
rect 27012 41860 27016 41916
rect 26952 41856 27016 41860
rect 27032 41916 27096 41920
rect 27032 41860 27036 41916
rect 27036 41860 27092 41916
rect 27092 41860 27096 41916
rect 27032 41856 27096 41860
rect 27112 41916 27176 41920
rect 27112 41860 27116 41916
rect 27116 41860 27172 41916
rect 27172 41860 27176 41916
rect 27112 41856 27176 41860
rect 27192 41916 27256 41920
rect 27192 41860 27196 41916
rect 27196 41860 27252 41916
rect 27252 41860 27256 41916
rect 27192 41856 27256 41860
rect 31952 41916 32016 41920
rect 31952 41860 31956 41916
rect 31956 41860 32012 41916
rect 32012 41860 32016 41916
rect 31952 41856 32016 41860
rect 32032 41916 32096 41920
rect 32032 41860 32036 41916
rect 32036 41860 32092 41916
rect 32092 41860 32096 41916
rect 32032 41856 32096 41860
rect 32112 41916 32176 41920
rect 32112 41860 32116 41916
rect 32116 41860 32172 41916
rect 32172 41860 32176 41916
rect 32112 41856 32176 41860
rect 32192 41916 32256 41920
rect 32192 41860 32196 41916
rect 32196 41860 32252 41916
rect 32252 41860 32256 41916
rect 32192 41856 32256 41860
rect 36952 41916 37016 41920
rect 36952 41860 36956 41916
rect 36956 41860 37012 41916
rect 37012 41860 37016 41916
rect 36952 41856 37016 41860
rect 37032 41916 37096 41920
rect 37032 41860 37036 41916
rect 37036 41860 37092 41916
rect 37092 41860 37096 41916
rect 37032 41856 37096 41860
rect 37112 41916 37176 41920
rect 37112 41860 37116 41916
rect 37116 41860 37172 41916
rect 37172 41860 37176 41916
rect 37112 41856 37176 41860
rect 37192 41916 37256 41920
rect 37192 41860 37196 41916
rect 37196 41860 37252 41916
rect 37252 41860 37256 41916
rect 37192 41856 37256 41860
rect 31708 41380 31772 41444
rect 32444 41380 32508 41444
rect 2612 41372 2676 41376
rect 2612 41316 2616 41372
rect 2616 41316 2672 41372
rect 2672 41316 2676 41372
rect 2612 41312 2676 41316
rect 2692 41372 2756 41376
rect 2692 41316 2696 41372
rect 2696 41316 2752 41372
rect 2752 41316 2756 41372
rect 2692 41312 2756 41316
rect 2772 41372 2836 41376
rect 2772 41316 2776 41372
rect 2776 41316 2832 41372
rect 2832 41316 2836 41372
rect 2772 41312 2836 41316
rect 2852 41372 2916 41376
rect 2852 41316 2856 41372
rect 2856 41316 2912 41372
rect 2912 41316 2916 41372
rect 2852 41312 2916 41316
rect 7612 41372 7676 41376
rect 7612 41316 7616 41372
rect 7616 41316 7672 41372
rect 7672 41316 7676 41372
rect 7612 41312 7676 41316
rect 7692 41372 7756 41376
rect 7692 41316 7696 41372
rect 7696 41316 7752 41372
rect 7752 41316 7756 41372
rect 7692 41312 7756 41316
rect 7772 41372 7836 41376
rect 7772 41316 7776 41372
rect 7776 41316 7832 41372
rect 7832 41316 7836 41372
rect 7772 41312 7836 41316
rect 7852 41372 7916 41376
rect 7852 41316 7856 41372
rect 7856 41316 7912 41372
rect 7912 41316 7916 41372
rect 7852 41312 7916 41316
rect 12612 41372 12676 41376
rect 12612 41316 12616 41372
rect 12616 41316 12672 41372
rect 12672 41316 12676 41372
rect 12612 41312 12676 41316
rect 12692 41372 12756 41376
rect 12692 41316 12696 41372
rect 12696 41316 12752 41372
rect 12752 41316 12756 41372
rect 12692 41312 12756 41316
rect 12772 41372 12836 41376
rect 12772 41316 12776 41372
rect 12776 41316 12832 41372
rect 12832 41316 12836 41372
rect 12772 41312 12836 41316
rect 12852 41372 12916 41376
rect 12852 41316 12856 41372
rect 12856 41316 12912 41372
rect 12912 41316 12916 41372
rect 12852 41312 12916 41316
rect 17612 41372 17676 41376
rect 17612 41316 17616 41372
rect 17616 41316 17672 41372
rect 17672 41316 17676 41372
rect 17612 41312 17676 41316
rect 17692 41372 17756 41376
rect 17692 41316 17696 41372
rect 17696 41316 17752 41372
rect 17752 41316 17756 41372
rect 17692 41312 17756 41316
rect 17772 41372 17836 41376
rect 17772 41316 17776 41372
rect 17776 41316 17832 41372
rect 17832 41316 17836 41372
rect 17772 41312 17836 41316
rect 17852 41372 17916 41376
rect 17852 41316 17856 41372
rect 17856 41316 17912 41372
rect 17912 41316 17916 41372
rect 17852 41312 17916 41316
rect 22612 41372 22676 41376
rect 22612 41316 22616 41372
rect 22616 41316 22672 41372
rect 22672 41316 22676 41372
rect 22612 41312 22676 41316
rect 22692 41372 22756 41376
rect 22692 41316 22696 41372
rect 22696 41316 22752 41372
rect 22752 41316 22756 41372
rect 22692 41312 22756 41316
rect 22772 41372 22836 41376
rect 22772 41316 22776 41372
rect 22776 41316 22832 41372
rect 22832 41316 22836 41372
rect 22772 41312 22836 41316
rect 22852 41372 22916 41376
rect 22852 41316 22856 41372
rect 22856 41316 22912 41372
rect 22912 41316 22916 41372
rect 22852 41312 22916 41316
rect 27612 41372 27676 41376
rect 27612 41316 27616 41372
rect 27616 41316 27672 41372
rect 27672 41316 27676 41372
rect 27612 41312 27676 41316
rect 27692 41372 27756 41376
rect 27692 41316 27696 41372
rect 27696 41316 27752 41372
rect 27752 41316 27756 41372
rect 27692 41312 27756 41316
rect 27772 41372 27836 41376
rect 27772 41316 27776 41372
rect 27776 41316 27832 41372
rect 27832 41316 27836 41372
rect 27772 41312 27836 41316
rect 27852 41372 27916 41376
rect 27852 41316 27856 41372
rect 27856 41316 27912 41372
rect 27912 41316 27916 41372
rect 27852 41312 27916 41316
rect 32612 41372 32676 41376
rect 32612 41316 32616 41372
rect 32616 41316 32672 41372
rect 32672 41316 32676 41372
rect 32612 41312 32676 41316
rect 32692 41372 32756 41376
rect 32692 41316 32696 41372
rect 32696 41316 32752 41372
rect 32752 41316 32756 41372
rect 32692 41312 32756 41316
rect 32772 41372 32836 41376
rect 32772 41316 32776 41372
rect 32776 41316 32832 41372
rect 32832 41316 32836 41372
rect 32772 41312 32836 41316
rect 32852 41372 32916 41376
rect 32852 41316 32856 41372
rect 32856 41316 32912 41372
rect 32912 41316 32916 41372
rect 32852 41312 32916 41316
rect 37612 41372 37676 41376
rect 37612 41316 37616 41372
rect 37616 41316 37672 41372
rect 37672 41316 37676 41372
rect 37612 41312 37676 41316
rect 37692 41372 37756 41376
rect 37692 41316 37696 41372
rect 37696 41316 37752 41372
rect 37752 41316 37756 41372
rect 37692 41312 37756 41316
rect 37772 41372 37836 41376
rect 37772 41316 37776 41372
rect 37776 41316 37832 41372
rect 37832 41316 37836 41372
rect 37772 41312 37836 41316
rect 37852 41372 37916 41376
rect 37852 41316 37856 41372
rect 37856 41316 37912 41372
rect 37912 41316 37916 41372
rect 37852 41312 37916 41316
rect 1952 40828 2016 40832
rect 1952 40772 1956 40828
rect 1956 40772 2012 40828
rect 2012 40772 2016 40828
rect 1952 40768 2016 40772
rect 2032 40828 2096 40832
rect 2032 40772 2036 40828
rect 2036 40772 2092 40828
rect 2092 40772 2096 40828
rect 2032 40768 2096 40772
rect 2112 40828 2176 40832
rect 2112 40772 2116 40828
rect 2116 40772 2172 40828
rect 2172 40772 2176 40828
rect 2112 40768 2176 40772
rect 2192 40828 2256 40832
rect 2192 40772 2196 40828
rect 2196 40772 2252 40828
rect 2252 40772 2256 40828
rect 2192 40768 2256 40772
rect 6952 40828 7016 40832
rect 6952 40772 6956 40828
rect 6956 40772 7012 40828
rect 7012 40772 7016 40828
rect 6952 40768 7016 40772
rect 7032 40828 7096 40832
rect 7032 40772 7036 40828
rect 7036 40772 7092 40828
rect 7092 40772 7096 40828
rect 7032 40768 7096 40772
rect 7112 40828 7176 40832
rect 7112 40772 7116 40828
rect 7116 40772 7172 40828
rect 7172 40772 7176 40828
rect 7112 40768 7176 40772
rect 7192 40828 7256 40832
rect 7192 40772 7196 40828
rect 7196 40772 7252 40828
rect 7252 40772 7256 40828
rect 7192 40768 7256 40772
rect 11952 40828 12016 40832
rect 11952 40772 11956 40828
rect 11956 40772 12012 40828
rect 12012 40772 12016 40828
rect 11952 40768 12016 40772
rect 12032 40828 12096 40832
rect 12032 40772 12036 40828
rect 12036 40772 12092 40828
rect 12092 40772 12096 40828
rect 12032 40768 12096 40772
rect 12112 40828 12176 40832
rect 12112 40772 12116 40828
rect 12116 40772 12172 40828
rect 12172 40772 12176 40828
rect 12112 40768 12176 40772
rect 12192 40828 12256 40832
rect 12192 40772 12196 40828
rect 12196 40772 12252 40828
rect 12252 40772 12256 40828
rect 12192 40768 12256 40772
rect 16952 40828 17016 40832
rect 16952 40772 16956 40828
rect 16956 40772 17012 40828
rect 17012 40772 17016 40828
rect 16952 40768 17016 40772
rect 17032 40828 17096 40832
rect 17032 40772 17036 40828
rect 17036 40772 17092 40828
rect 17092 40772 17096 40828
rect 17032 40768 17096 40772
rect 17112 40828 17176 40832
rect 17112 40772 17116 40828
rect 17116 40772 17172 40828
rect 17172 40772 17176 40828
rect 17112 40768 17176 40772
rect 17192 40828 17256 40832
rect 17192 40772 17196 40828
rect 17196 40772 17252 40828
rect 17252 40772 17256 40828
rect 17192 40768 17256 40772
rect 21952 40828 22016 40832
rect 21952 40772 21956 40828
rect 21956 40772 22012 40828
rect 22012 40772 22016 40828
rect 21952 40768 22016 40772
rect 22032 40828 22096 40832
rect 22032 40772 22036 40828
rect 22036 40772 22092 40828
rect 22092 40772 22096 40828
rect 22032 40768 22096 40772
rect 22112 40828 22176 40832
rect 22112 40772 22116 40828
rect 22116 40772 22172 40828
rect 22172 40772 22176 40828
rect 22112 40768 22176 40772
rect 22192 40828 22256 40832
rect 22192 40772 22196 40828
rect 22196 40772 22252 40828
rect 22252 40772 22256 40828
rect 22192 40768 22256 40772
rect 26952 40828 27016 40832
rect 26952 40772 26956 40828
rect 26956 40772 27012 40828
rect 27012 40772 27016 40828
rect 26952 40768 27016 40772
rect 27032 40828 27096 40832
rect 27032 40772 27036 40828
rect 27036 40772 27092 40828
rect 27092 40772 27096 40828
rect 27032 40768 27096 40772
rect 27112 40828 27176 40832
rect 27112 40772 27116 40828
rect 27116 40772 27172 40828
rect 27172 40772 27176 40828
rect 27112 40768 27176 40772
rect 27192 40828 27256 40832
rect 27192 40772 27196 40828
rect 27196 40772 27252 40828
rect 27252 40772 27256 40828
rect 27192 40768 27256 40772
rect 31952 40828 32016 40832
rect 31952 40772 31956 40828
rect 31956 40772 32012 40828
rect 32012 40772 32016 40828
rect 31952 40768 32016 40772
rect 32032 40828 32096 40832
rect 32032 40772 32036 40828
rect 32036 40772 32092 40828
rect 32092 40772 32096 40828
rect 32032 40768 32096 40772
rect 32112 40828 32176 40832
rect 32112 40772 32116 40828
rect 32116 40772 32172 40828
rect 32172 40772 32176 40828
rect 32112 40768 32176 40772
rect 32192 40828 32256 40832
rect 32192 40772 32196 40828
rect 32196 40772 32252 40828
rect 32252 40772 32256 40828
rect 32192 40768 32256 40772
rect 36952 40828 37016 40832
rect 36952 40772 36956 40828
rect 36956 40772 37012 40828
rect 37012 40772 37016 40828
rect 36952 40768 37016 40772
rect 37032 40828 37096 40832
rect 37032 40772 37036 40828
rect 37036 40772 37092 40828
rect 37092 40772 37096 40828
rect 37032 40768 37096 40772
rect 37112 40828 37176 40832
rect 37112 40772 37116 40828
rect 37116 40772 37172 40828
rect 37172 40772 37176 40828
rect 37112 40768 37176 40772
rect 37192 40828 37256 40832
rect 37192 40772 37196 40828
rect 37196 40772 37252 40828
rect 37252 40772 37256 40828
rect 37192 40768 37256 40772
rect 2612 40284 2676 40288
rect 2612 40228 2616 40284
rect 2616 40228 2672 40284
rect 2672 40228 2676 40284
rect 2612 40224 2676 40228
rect 2692 40284 2756 40288
rect 2692 40228 2696 40284
rect 2696 40228 2752 40284
rect 2752 40228 2756 40284
rect 2692 40224 2756 40228
rect 2772 40284 2836 40288
rect 2772 40228 2776 40284
rect 2776 40228 2832 40284
rect 2832 40228 2836 40284
rect 2772 40224 2836 40228
rect 2852 40284 2916 40288
rect 2852 40228 2856 40284
rect 2856 40228 2912 40284
rect 2912 40228 2916 40284
rect 2852 40224 2916 40228
rect 7612 40284 7676 40288
rect 7612 40228 7616 40284
rect 7616 40228 7672 40284
rect 7672 40228 7676 40284
rect 7612 40224 7676 40228
rect 7692 40284 7756 40288
rect 7692 40228 7696 40284
rect 7696 40228 7752 40284
rect 7752 40228 7756 40284
rect 7692 40224 7756 40228
rect 7772 40284 7836 40288
rect 7772 40228 7776 40284
rect 7776 40228 7832 40284
rect 7832 40228 7836 40284
rect 7772 40224 7836 40228
rect 7852 40284 7916 40288
rect 7852 40228 7856 40284
rect 7856 40228 7912 40284
rect 7912 40228 7916 40284
rect 7852 40224 7916 40228
rect 12612 40284 12676 40288
rect 12612 40228 12616 40284
rect 12616 40228 12672 40284
rect 12672 40228 12676 40284
rect 12612 40224 12676 40228
rect 12692 40284 12756 40288
rect 12692 40228 12696 40284
rect 12696 40228 12752 40284
rect 12752 40228 12756 40284
rect 12692 40224 12756 40228
rect 12772 40284 12836 40288
rect 12772 40228 12776 40284
rect 12776 40228 12832 40284
rect 12832 40228 12836 40284
rect 12772 40224 12836 40228
rect 12852 40284 12916 40288
rect 12852 40228 12856 40284
rect 12856 40228 12912 40284
rect 12912 40228 12916 40284
rect 12852 40224 12916 40228
rect 17612 40284 17676 40288
rect 17612 40228 17616 40284
rect 17616 40228 17672 40284
rect 17672 40228 17676 40284
rect 17612 40224 17676 40228
rect 17692 40284 17756 40288
rect 17692 40228 17696 40284
rect 17696 40228 17752 40284
rect 17752 40228 17756 40284
rect 17692 40224 17756 40228
rect 17772 40284 17836 40288
rect 17772 40228 17776 40284
rect 17776 40228 17832 40284
rect 17832 40228 17836 40284
rect 17772 40224 17836 40228
rect 17852 40284 17916 40288
rect 17852 40228 17856 40284
rect 17856 40228 17912 40284
rect 17912 40228 17916 40284
rect 17852 40224 17916 40228
rect 22612 40284 22676 40288
rect 22612 40228 22616 40284
rect 22616 40228 22672 40284
rect 22672 40228 22676 40284
rect 22612 40224 22676 40228
rect 22692 40284 22756 40288
rect 22692 40228 22696 40284
rect 22696 40228 22752 40284
rect 22752 40228 22756 40284
rect 22692 40224 22756 40228
rect 22772 40284 22836 40288
rect 22772 40228 22776 40284
rect 22776 40228 22832 40284
rect 22832 40228 22836 40284
rect 22772 40224 22836 40228
rect 22852 40284 22916 40288
rect 22852 40228 22856 40284
rect 22856 40228 22912 40284
rect 22912 40228 22916 40284
rect 22852 40224 22916 40228
rect 27612 40284 27676 40288
rect 27612 40228 27616 40284
rect 27616 40228 27672 40284
rect 27672 40228 27676 40284
rect 27612 40224 27676 40228
rect 27692 40284 27756 40288
rect 27692 40228 27696 40284
rect 27696 40228 27752 40284
rect 27752 40228 27756 40284
rect 27692 40224 27756 40228
rect 27772 40284 27836 40288
rect 27772 40228 27776 40284
rect 27776 40228 27832 40284
rect 27832 40228 27836 40284
rect 27772 40224 27836 40228
rect 27852 40284 27916 40288
rect 27852 40228 27856 40284
rect 27856 40228 27912 40284
rect 27912 40228 27916 40284
rect 27852 40224 27916 40228
rect 32612 40284 32676 40288
rect 32612 40228 32616 40284
rect 32616 40228 32672 40284
rect 32672 40228 32676 40284
rect 32612 40224 32676 40228
rect 32692 40284 32756 40288
rect 32692 40228 32696 40284
rect 32696 40228 32752 40284
rect 32752 40228 32756 40284
rect 32692 40224 32756 40228
rect 32772 40284 32836 40288
rect 32772 40228 32776 40284
rect 32776 40228 32832 40284
rect 32832 40228 32836 40284
rect 32772 40224 32836 40228
rect 32852 40284 32916 40288
rect 32852 40228 32856 40284
rect 32856 40228 32912 40284
rect 32912 40228 32916 40284
rect 32852 40224 32916 40228
rect 37612 40284 37676 40288
rect 37612 40228 37616 40284
rect 37616 40228 37672 40284
rect 37672 40228 37676 40284
rect 37612 40224 37676 40228
rect 37692 40284 37756 40288
rect 37692 40228 37696 40284
rect 37696 40228 37752 40284
rect 37752 40228 37756 40284
rect 37692 40224 37756 40228
rect 37772 40284 37836 40288
rect 37772 40228 37776 40284
rect 37776 40228 37832 40284
rect 37832 40228 37836 40284
rect 37772 40224 37836 40228
rect 37852 40284 37916 40288
rect 37852 40228 37856 40284
rect 37856 40228 37912 40284
rect 37912 40228 37916 40284
rect 37852 40224 37916 40228
rect 1952 39740 2016 39744
rect 1952 39684 1956 39740
rect 1956 39684 2012 39740
rect 2012 39684 2016 39740
rect 1952 39680 2016 39684
rect 2032 39740 2096 39744
rect 2032 39684 2036 39740
rect 2036 39684 2092 39740
rect 2092 39684 2096 39740
rect 2032 39680 2096 39684
rect 2112 39740 2176 39744
rect 2112 39684 2116 39740
rect 2116 39684 2172 39740
rect 2172 39684 2176 39740
rect 2112 39680 2176 39684
rect 2192 39740 2256 39744
rect 2192 39684 2196 39740
rect 2196 39684 2252 39740
rect 2252 39684 2256 39740
rect 2192 39680 2256 39684
rect 6952 39740 7016 39744
rect 6952 39684 6956 39740
rect 6956 39684 7012 39740
rect 7012 39684 7016 39740
rect 6952 39680 7016 39684
rect 7032 39740 7096 39744
rect 7032 39684 7036 39740
rect 7036 39684 7092 39740
rect 7092 39684 7096 39740
rect 7032 39680 7096 39684
rect 7112 39740 7176 39744
rect 7112 39684 7116 39740
rect 7116 39684 7172 39740
rect 7172 39684 7176 39740
rect 7112 39680 7176 39684
rect 7192 39740 7256 39744
rect 7192 39684 7196 39740
rect 7196 39684 7252 39740
rect 7252 39684 7256 39740
rect 7192 39680 7256 39684
rect 11952 39740 12016 39744
rect 11952 39684 11956 39740
rect 11956 39684 12012 39740
rect 12012 39684 12016 39740
rect 11952 39680 12016 39684
rect 12032 39740 12096 39744
rect 12032 39684 12036 39740
rect 12036 39684 12092 39740
rect 12092 39684 12096 39740
rect 12032 39680 12096 39684
rect 12112 39740 12176 39744
rect 12112 39684 12116 39740
rect 12116 39684 12172 39740
rect 12172 39684 12176 39740
rect 12112 39680 12176 39684
rect 12192 39740 12256 39744
rect 12192 39684 12196 39740
rect 12196 39684 12252 39740
rect 12252 39684 12256 39740
rect 12192 39680 12256 39684
rect 16952 39740 17016 39744
rect 16952 39684 16956 39740
rect 16956 39684 17012 39740
rect 17012 39684 17016 39740
rect 16952 39680 17016 39684
rect 17032 39740 17096 39744
rect 17032 39684 17036 39740
rect 17036 39684 17092 39740
rect 17092 39684 17096 39740
rect 17032 39680 17096 39684
rect 17112 39740 17176 39744
rect 17112 39684 17116 39740
rect 17116 39684 17172 39740
rect 17172 39684 17176 39740
rect 17112 39680 17176 39684
rect 17192 39740 17256 39744
rect 17192 39684 17196 39740
rect 17196 39684 17252 39740
rect 17252 39684 17256 39740
rect 17192 39680 17256 39684
rect 21952 39740 22016 39744
rect 21952 39684 21956 39740
rect 21956 39684 22012 39740
rect 22012 39684 22016 39740
rect 21952 39680 22016 39684
rect 22032 39740 22096 39744
rect 22032 39684 22036 39740
rect 22036 39684 22092 39740
rect 22092 39684 22096 39740
rect 22032 39680 22096 39684
rect 22112 39740 22176 39744
rect 22112 39684 22116 39740
rect 22116 39684 22172 39740
rect 22172 39684 22176 39740
rect 22112 39680 22176 39684
rect 22192 39740 22256 39744
rect 22192 39684 22196 39740
rect 22196 39684 22252 39740
rect 22252 39684 22256 39740
rect 22192 39680 22256 39684
rect 26952 39740 27016 39744
rect 26952 39684 26956 39740
rect 26956 39684 27012 39740
rect 27012 39684 27016 39740
rect 26952 39680 27016 39684
rect 27032 39740 27096 39744
rect 27032 39684 27036 39740
rect 27036 39684 27092 39740
rect 27092 39684 27096 39740
rect 27032 39680 27096 39684
rect 27112 39740 27176 39744
rect 27112 39684 27116 39740
rect 27116 39684 27172 39740
rect 27172 39684 27176 39740
rect 27112 39680 27176 39684
rect 27192 39740 27256 39744
rect 27192 39684 27196 39740
rect 27196 39684 27252 39740
rect 27252 39684 27256 39740
rect 27192 39680 27256 39684
rect 31952 39740 32016 39744
rect 31952 39684 31956 39740
rect 31956 39684 32012 39740
rect 32012 39684 32016 39740
rect 31952 39680 32016 39684
rect 32032 39740 32096 39744
rect 32032 39684 32036 39740
rect 32036 39684 32092 39740
rect 32092 39684 32096 39740
rect 32032 39680 32096 39684
rect 32112 39740 32176 39744
rect 32112 39684 32116 39740
rect 32116 39684 32172 39740
rect 32172 39684 32176 39740
rect 32112 39680 32176 39684
rect 32192 39740 32256 39744
rect 32192 39684 32196 39740
rect 32196 39684 32252 39740
rect 32252 39684 32256 39740
rect 32192 39680 32256 39684
rect 36952 39740 37016 39744
rect 36952 39684 36956 39740
rect 36956 39684 37012 39740
rect 37012 39684 37016 39740
rect 36952 39680 37016 39684
rect 37032 39740 37096 39744
rect 37032 39684 37036 39740
rect 37036 39684 37092 39740
rect 37092 39684 37096 39740
rect 37032 39680 37096 39684
rect 37112 39740 37176 39744
rect 37112 39684 37116 39740
rect 37116 39684 37172 39740
rect 37172 39684 37176 39740
rect 37112 39680 37176 39684
rect 37192 39740 37256 39744
rect 37192 39684 37196 39740
rect 37196 39684 37252 39740
rect 37252 39684 37256 39740
rect 37192 39680 37256 39684
rect 2612 39196 2676 39200
rect 2612 39140 2616 39196
rect 2616 39140 2672 39196
rect 2672 39140 2676 39196
rect 2612 39136 2676 39140
rect 2692 39196 2756 39200
rect 2692 39140 2696 39196
rect 2696 39140 2752 39196
rect 2752 39140 2756 39196
rect 2692 39136 2756 39140
rect 2772 39196 2836 39200
rect 2772 39140 2776 39196
rect 2776 39140 2832 39196
rect 2832 39140 2836 39196
rect 2772 39136 2836 39140
rect 2852 39196 2916 39200
rect 2852 39140 2856 39196
rect 2856 39140 2912 39196
rect 2912 39140 2916 39196
rect 2852 39136 2916 39140
rect 7612 39196 7676 39200
rect 7612 39140 7616 39196
rect 7616 39140 7672 39196
rect 7672 39140 7676 39196
rect 7612 39136 7676 39140
rect 7692 39196 7756 39200
rect 7692 39140 7696 39196
rect 7696 39140 7752 39196
rect 7752 39140 7756 39196
rect 7692 39136 7756 39140
rect 7772 39196 7836 39200
rect 7772 39140 7776 39196
rect 7776 39140 7832 39196
rect 7832 39140 7836 39196
rect 7772 39136 7836 39140
rect 7852 39196 7916 39200
rect 7852 39140 7856 39196
rect 7856 39140 7912 39196
rect 7912 39140 7916 39196
rect 7852 39136 7916 39140
rect 12612 39196 12676 39200
rect 12612 39140 12616 39196
rect 12616 39140 12672 39196
rect 12672 39140 12676 39196
rect 12612 39136 12676 39140
rect 12692 39196 12756 39200
rect 12692 39140 12696 39196
rect 12696 39140 12752 39196
rect 12752 39140 12756 39196
rect 12692 39136 12756 39140
rect 12772 39196 12836 39200
rect 12772 39140 12776 39196
rect 12776 39140 12832 39196
rect 12832 39140 12836 39196
rect 12772 39136 12836 39140
rect 12852 39196 12916 39200
rect 12852 39140 12856 39196
rect 12856 39140 12912 39196
rect 12912 39140 12916 39196
rect 12852 39136 12916 39140
rect 17612 39196 17676 39200
rect 17612 39140 17616 39196
rect 17616 39140 17672 39196
rect 17672 39140 17676 39196
rect 17612 39136 17676 39140
rect 17692 39196 17756 39200
rect 17692 39140 17696 39196
rect 17696 39140 17752 39196
rect 17752 39140 17756 39196
rect 17692 39136 17756 39140
rect 17772 39196 17836 39200
rect 17772 39140 17776 39196
rect 17776 39140 17832 39196
rect 17832 39140 17836 39196
rect 17772 39136 17836 39140
rect 17852 39196 17916 39200
rect 17852 39140 17856 39196
rect 17856 39140 17912 39196
rect 17912 39140 17916 39196
rect 17852 39136 17916 39140
rect 22612 39196 22676 39200
rect 22612 39140 22616 39196
rect 22616 39140 22672 39196
rect 22672 39140 22676 39196
rect 22612 39136 22676 39140
rect 22692 39196 22756 39200
rect 22692 39140 22696 39196
rect 22696 39140 22752 39196
rect 22752 39140 22756 39196
rect 22692 39136 22756 39140
rect 22772 39196 22836 39200
rect 22772 39140 22776 39196
rect 22776 39140 22832 39196
rect 22832 39140 22836 39196
rect 22772 39136 22836 39140
rect 22852 39196 22916 39200
rect 22852 39140 22856 39196
rect 22856 39140 22912 39196
rect 22912 39140 22916 39196
rect 22852 39136 22916 39140
rect 27612 39196 27676 39200
rect 27612 39140 27616 39196
rect 27616 39140 27672 39196
rect 27672 39140 27676 39196
rect 27612 39136 27676 39140
rect 27692 39196 27756 39200
rect 27692 39140 27696 39196
rect 27696 39140 27752 39196
rect 27752 39140 27756 39196
rect 27692 39136 27756 39140
rect 27772 39196 27836 39200
rect 27772 39140 27776 39196
rect 27776 39140 27832 39196
rect 27832 39140 27836 39196
rect 27772 39136 27836 39140
rect 27852 39196 27916 39200
rect 27852 39140 27856 39196
rect 27856 39140 27912 39196
rect 27912 39140 27916 39196
rect 27852 39136 27916 39140
rect 32612 39196 32676 39200
rect 32612 39140 32616 39196
rect 32616 39140 32672 39196
rect 32672 39140 32676 39196
rect 32612 39136 32676 39140
rect 32692 39196 32756 39200
rect 32692 39140 32696 39196
rect 32696 39140 32752 39196
rect 32752 39140 32756 39196
rect 32692 39136 32756 39140
rect 32772 39196 32836 39200
rect 32772 39140 32776 39196
rect 32776 39140 32832 39196
rect 32832 39140 32836 39196
rect 32772 39136 32836 39140
rect 32852 39196 32916 39200
rect 32852 39140 32856 39196
rect 32856 39140 32912 39196
rect 32912 39140 32916 39196
rect 32852 39136 32916 39140
rect 37612 39196 37676 39200
rect 37612 39140 37616 39196
rect 37616 39140 37672 39196
rect 37672 39140 37676 39196
rect 37612 39136 37676 39140
rect 37692 39196 37756 39200
rect 37692 39140 37696 39196
rect 37696 39140 37752 39196
rect 37752 39140 37756 39196
rect 37692 39136 37756 39140
rect 37772 39196 37836 39200
rect 37772 39140 37776 39196
rect 37776 39140 37832 39196
rect 37832 39140 37836 39196
rect 37772 39136 37836 39140
rect 37852 39196 37916 39200
rect 37852 39140 37856 39196
rect 37856 39140 37912 39196
rect 37912 39140 37916 39196
rect 37852 39136 37916 39140
rect 1952 38652 2016 38656
rect 1952 38596 1956 38652
rect 1956 38596 2012 38652
rect 2012 38596 2016 38652
rect 1952 38592 2016 38596
rect 2032 38652 2096 38656
rect 2032 38596 2036 38652
rect 2036 38596 2092 38652
rect 2092 38596 2096 38652
rect 2032 38592 2096 38596
rect 2112 38652 2176 38656
rect 2112 38596 2116 38652
rect 2116 38596 2172 38652
rect 2172 38596 2176 38652
rect 2112 38592 2176 38596
rect 2192 38652 2256 38656
rect 2192 38596 2196 38652
rect 2196 38596 2252 38652
rect 2252 38596 2256 38652
rect 2192 38592 2256 38596
rect 6952 38652 7016 38656
rect 6952 38596 6956 38652
rect 6956 38596 7012 38652
rect 7012 38596 7016 38652
rect 6952 38592 7016 38596
rect 7032 38652 7096 38656
rect 7032 38596 7036 38652
rect 7036 38596 7092 38652
rect 7092 38596 7096 38652
rect 7032 38592 7096 38596
rect 7112 38652 7176 38656
rect 7112 38596 7116 38652
rect 7116 38596 7172 38652
rect 7172 38596 7176 38652
rect 7112 38592 7176 38596
rect 7192 38652 7256 38656
rect 7192 38596 7196 38652
rect 7196 38596 7252 38652
rect 7252 38596 7256 38652
rect 7192 38592 7256 38596
rect 11952 38652 12016 38656
rect 11952 38596 11956 38652
rect 11956 38596 12012 38652
rect 12012 38596 12016 38652
rect 11952 38592 12016 38596
rect 12032 38652 12096 38656
rect 12032 38596 12036 38652
rect 12036 38596 12092 38652
rect 12092 38596 12096 38652
rect 12032 38592 12096 38596
rect 12112 38652 12176 38656
rect 12112 38596 12116 38652
rect 12116 38596 12172 38652
rect 12172 38596 12176 38652
rect 12112 38592 12176 38596
rect 12192 38652 12256 38656
rect 12192 38596 12196 38652
rect 12196 38596 12252 38652
rect 12252 38596 12256 38652
rect 12192 38592 12256 38596
rect 16952 38652 17016 38656
rect 16952 38596 16956 38652
rect 16956 38596 17012 38652
rect 17012 38596 17016 38652
rect 16952 38592 17016 38596
rect 17032 38652 17096 38656
rect 17032 38596 17036 38652
rect 17036 38596 17092 38652
rect 17092 38596 17096 38652
rect 17032 38592 17096 38596
rect 17112 38652 17176 38656
rect 17112 38596 17116 38652
rect 17116 38596 17172 38652
rect 17172 38596 17176 38652
rect 17112 38592 17176 38596
rect 17192 38652 17256 38656
rect 17192 38596 17196 38652
rect 17196 38596 17252 38652
rect 17252 38596 17256 38652
rect 17192 38592 17256 38596
rect 21952 38652 22016 38656
rect 21952 38596 21956 38652
rect 21956 38596 22012 38652
rect 22012 38596 22016 38652
rect 21952 38592 22016 38596
rect 22032 38652 22096 38656
rect 22032 38596 22036 38652
rect 22036 38596 22092 38652
rect 22092 38596 22096 38652
rect 22032 38592 22096 38596
rect 22112 38652 22176 38656
rect 22112 38596 22116 38652
rect 22116 38596 22172 38652
rect 22172 38596 22176 38652
rect 22112 38592 22176 38596
rect 22192 38652 22256 38656
rect 22192 38596 22196 38652
rect 22196 38596 22252 38652
rect 22252 38596 22256 38652
rect 22192 38592 22256 38596
rect 26952 38652 27016 38656
rect 26952 38596 26956 38652
rect 26956 38596 27012 38652
rect 27012 38596 27016 38652
rect 26952 38592 27016 38596
rect 27032 38652 27096 38656
rect 27032 38596 27036 38652
rect 27036 38596 27092 38652
rect 27092 38596 27096 38652
rect 27032 38592 27096 38596
rect 27112 38652 27176 38656
rect 27112 38596 27116 38652
rect 27116 38596 27172 38652
rect 27172 38596 27176 38652
rect 27112 38592 27176 38596
rect 27192 38652 27256 38656
rect 27192 38596 27196 38652
rect 27196 38596 27252 38652
rect 27252 38596 27256 38652
rect 27192 38592 27256 38596
rect 31952 38652 32016 38656
rect 31952 38596 31956 38652
rect 31956 38596 32012 38652
rect 32012 38596 32016 38652
rect 31952 38592 32016 38596
rect 32032 38652 32096 38656
rect 32032 38596 32036 38652
rect 32036 38596 32092 38652
rect 32092 38596 32096 38652
rect 32032 38592 32096 38596
rect 32112 38652 32176 38656
rect 32112 38596 32116 38652
rect 32116 38596 32172 38652
rect 32172 38596 32176 38652
rect 32112 38592 32176 38596
rect 32192 38652 32256 38656
rect 32192 38596 32196 38652
rect 32196 38596 32252 38652
rect 32252 38596 32256 38652
rect 32192 38592 32256 38596
rect 36952 38652 37016 38656
rect 36952 38596 36956 38652
rect 36956 38596 37012 38652
rect 37012 38596 37016 38652
rect 36952 38592 37016 38596
rect 37032 38652 37096 38656
rect 37032 38596 37036 38652
rect 37036 38596 37092 38652
rect 37092 38596 37096 38652
rect 37032 38592 37096 38596
rect 37112 38652 37176 38656
rect 37112 38596 37116 38652
rect 37116 38596 37172 38652
rect 37172 38596 37176 38652
rect 37112 38592 37176 38596
rect 37192 38652 37256 38656
rect 37192 38596 37196 38652
rect 37196 38596 37252 38652
rect 37252 38596 37256 38652
rect 37192 38592 37256 38596
rect 2612 38108 2676 38112
rect 2612 38052 2616 38108
rect 2616 38052 2672 38108
rect 2672 38052 2676 38108
rect 2612 38048 2676 38052
rect 2692 38108 2756 38112
rect 2692 38052 2696 38108
rect 2696 38052 2752 38108
rect 2752 38052 2756 38108
rect 2692 38048 2756 38052
rect 2772 38108 2836 38112
rect 2772 38052 2776 38108
rect 2776 38052 2832 38108
rect 2832 38052 2836 38108
rect 2772 38048 2836 38052
rect 2852 38108 2916 38112
rect 2852 38052 2856 38108
rect 2856 38052 2912 38108
rect 2912 38052 2916 38108
rect 2852 38048 2916 38052
rect 7612 38108 7676 38112
rect 7612 38052 7616 38108
rect 7616 38052 7672 38108
rect 7672 38052 7676 38108
rect 7612 38048 7676 38052
rect 7692 38108 7756 38112
rect 7692 38052 7696 38108
rect 7696 38052 7752 38108
rect 7752 38052 7756 38108
rect 7692 38048 7756 38052
rect 7772 38108 7836 38112
rect 7772 38052 7776 38108
rect 7776 38052 7832 38108
rect 7832 38052 7836 38108
rect 7772 38048 7836 38052
rect 7852 38108 7916 38112
rect 7852 38052 7856 38108
rect 7856 38052 7912 38108
rect 7912 38052 7916 38108
rect 7852 38048 7916 38052
rect 12612 38108 12676 38112
rect 12612 38052 12616 38108
rect 12616 38052 12672 38108
rect 12672 38052 12676 38108
rect 12612 38048 12676 38052
rect 12692 38108 12756 38112
rect 12692 38052 12696 38108
rect 12696 38052 12752 38108
rect 12752 38052 12756 38108
rect 12692 38048 12756 38052
rect 12772 38108 12836 38112
rect 12772 38052 12776 38108
rect 12776 38052 12832 38108
rect 12832 38052 12836 38108
rect 12772 38048 12836 38052
rect 12852 38108 12916 38112
rect 12852 38052 12856 38108
rect 12856 38052 12912 38108
rect 12912 38052 12916 38108
rect 12852 38048 12916 38052
rect 17612 38108 17676 38112
rect 17612 38052 17616 38108
rect 17616 38052 17672 38108
rect 17672 38052 17676 38108
rect 17612 38048 17676 38052
rect 17692 38108 17756 38112
rect 17692 38052 17696 38108
rect 17696 38052 17752 38108
rect 17752 38052 17756 38108
rect 17692 38048 17756 38052
rect 17772 38108 17836 38112
rect 17772 38052 17776 38108
rect 17776 38052 17832 38108
rect 17832 38052 17836 38108
rect 17772 38048 17836 38052
rect 17852 38108 17916 38112
rect 17852 38052 17856 38108
rect 17856 38052 17912 38108
rect 17912 38052 17916 38108
rect 17852 38048 17916 38052
rect 22612 38108 22676 38112
rect 22612 38052 22616 38108
rect 22616 38052 22672 38108
rect 22672 38052 22676 38108
rect 22612 38048 22676 38052
rect 22692 38108 22756 38112
rect 22692 38052 22696 38108
rect 22696 38052 22752 38108
rect 22752 38052 22756 38108
rect 22692 38048 22756 38052
rect 22772 38108 22836 38112
rect 22772 38052 22776 38108
rect 22776 38052 22832 38108
rect 22832 38052 22836 38108
rect 22772 38048 22836 38052
rect 22852 38108 22916 38112
rect 22852 38052 22856 38108
rect 22856 38052 22912 38108
rect 22912 38052 22916 38108
rect 22852 38048 22916 38052
rect 27612 38108 27676 38112
rect 27612 38052 27616 38108
rect 27616 38052 27672 38108
rect 27672 38052 27676 38108
rect 27612 38048 27676 38052
rect 27692 38108 27756 38112
rect 27692 38052 27696 38108
rect 27696 38052 27752 38108
rect 27752 38052 27756 38108
rect 27692 38048 27756 38052
rect 27772 38108 27836 38112
rect 27772 38052 27776 38108
rect 27776 38052 27832 38108
rect 27832 38052 27836 38108
rect 27772 38048 27836 38052
rect 27852 38108 27916 38112
rect 27852 38052 27856 38108
rect 27856 38052 27912 38108
rect 27912 38052 27916 38108
rect 27852 38048 27916 38052
rect 32612 38108 32676 38112
rect 32612 38052 32616 38108
rect 32616 38052 32672 38108
rect 32672 38052 32676 38108
rect 32612 38048 32676 38052
rect 32692 38108 32756 38112
rect 32692 38052 32696 38108
rect 32696 38052 32752 38108
rect 32752 38052 32756 38108
rect 32692 38048 32756 38052
rect 32772 38108 32836 38112
rect 32772 38052 32776 38108
rect 32776 38052 32832 38108
rect 32832 38052 32836 38108
rect 32772 38048 32836 38052
rect 32852 38108 32916 38112
rect 32852 38052 32856 38108
rect 32856 38052 32912 38108
rect 32912 38052 32916 38108
rect 32852 38048 32916 38052
rect 37612 38108 37676 38112
rect 37612 38052 37616 38108
rect 37616 38052 37672 38108
rect 37672 38052 37676 38108
rect 37612 38048 37676 38052
rect 37692 38108 37756 38112
rect 37692 38052 37696 38108
rect 37696 38052 37752 38108
rect 37752 38052 37756 38108
rect 37692 38048 37756 38052
rect 37772 38108 37836 38112
rect 37772 38052 37776 38108
rect 37776 38052 37832 38108
rect 37832 38052 37836 38108
rect 37772 38048 37836 38052
rect 37852 38108 37916 38112
rect 37852 38052 37856 38108
rect 37856 38052 37912 38108
rect 37912 38052 37916 38108
rect 37852 38048 37916 38052
rect 1952 37564 2016 37568
rect 1952 37508 1956 37564
rect 1956 37508 2012 37564
rect 2012 37508 2016 37564
rect 1952 37504 2016 37508
rect 2032 37564 2096 37568
rect 2032 37508 2036 37564
rect 2036 37508 2092 37564
rect 2092 37508 2096 37564
rect 2032 37504 2096 37508
rect 2112 37564 2176 37568
rect 2112 37508 2116 37564
rect 2116 37508 2172 37564
rect 2172 37508 2176 37564
rect 2112 37504 2176 37508
rect 2192 37564 2256 37568
rect 2192 37508 2196 37564
rect 2196 37508 2252 37564
rect 2252 37508 2256 37564
rect 2192 37504 2256 37508
rect 6952 37564 7016 37568
rect 6952 37508 6956 37564
rect 6956 37508 7012 37564
rect 7012 37508 7016 37564
rect 6952 37504 7016 37508
rect 7032 37564 7096 37568
rect 7032 37508 7036 37564
rect 7036 37508 7092 37564
rect 7092 37508 7096 37564
rect 7032 37504 7096 37508
rect 7112 37564 7176 37568
rect 7112 37508 7116 37564
rect 7116 37508 7172 37564
rect 7172 37508 7176 37564
rect 7112 37504 7176 37508
rect 7192 37564 7256 37568
rect 7192 37508 7196 37564
rect 7196 37508 7252 37564
rect 7252 37508 7256 37564
rect 7192 37504 7256 37508
rect 11952 37564 12016 37568
rect 11952 37508 11956 37564
rect 11956 37508 12012 37564
rect 12012 37508 12016 37564
rect 11952 37504 12016 37508
rect 12032 37564 12096 37568
rect 12032 37508 12036 37564
rect 12036 37508 12092 37564
rect 12092 37508 12096 37564
rect 12032 37504 12096 37508
rect 12112 37564 12176 37568
rect 12112 37508 12116 37564
rect 12116 37508 12172 37564
rect 12172 37508 12176 37564
rect 12112 37504 12176 37508
rect 12192 37564 12256 37568
rect 12192 37508 12196 37564
rect 12196 37508 12252 37564
rect 12252 37508 12256 37564
rect 12192 37504 12256 37508
rect 16952 37564 17016 37568
rect 16952 37508 16956 37564
rect 16956 37508 17012 37564
rect 17012 37508 17016 37564
rect 16952 37504 17016 37508
rect 17032 37564 17096 37568
rect 17032 37508 17036 37564
rect 17036 37508 17092 37564
rect 17092 37508 17096 37564
rect 17032 37504 17096 37508
rect 17112 37564 17176 37568
rect 17112 37508 17116 37564
rect 17116 37508 17172 37564
rect 17172 37508 17176 37564
rect 17112 37504 17176 37508
rect 17192 37564 17256 37568
rect 17192 37508 17196 37564
rect 17196 37508 17252 37564
rect 17252 37508 17256 37564
rect 17192 37504 17256 37508
rect 21952 37564 22016 37568
rect 21952 37508 21956 37564
rect 21956 37508 22012 37564
rect 22012 37508 22016 37564
rect 21952 37504 22016 37508
rect 22032 37564 22096 37568
rect 22032 37508 22036 37564
rect 22036 37508 22092 37564
rect 22092 37508 22096 37564
rect 22032 37504 22096 37508
rect 22112 37564 22176 37568
rect 22112 37508 22116 37564
rect 22116 37508 22172 37564
rect 22172 37508 22176 37564
rect 22112 37504 22176 37508
rect 22192 37564 22256 37568
rect 22192 37508 22196 37564
rect 22196 37508 22252 37564
rect 22252 37508 22256 37564
rect 22192 37504 22256 37508
rect 26952 37564 27016 37568
rect 26952 37508 26956 37564
rect 26956 37508 27012 37564
rect 27012 37508 27016 37564
rect 26952 37504 27016 37508
rect 27032 37564 27096 37568
rect 27032 37508 27036 37564
rect 27036 37508 27092 37564
rect 27092 37508 27096 37564
rect 27032 37504 27096 37508
rect 27112 37564 27176 37568
rect 27112 37508 27116 37564
rect 27116 37508 27172 37564
rect 27172 37508 27176 37564
rect 27112 37504 27176 37508
rect 27192 37564 27256 37568
rect 27192 37508 27196 37564
rect 27196 37508 27252 37564
rect 27252 37508 27256 37564
rect 27192 37504 27256 37508
rect 31952 37564 32016 37568
rect 31952 37508 31956 37564
rect 31956 37508 32012 37564
rect 32012 37508 32016 37564
rect 31952 37504 32016 37508
rect 32032 37564 32096 37568
rect 32032 37508 32036 37564
rect 32036 37508 32092 37564
rect 32092 37508 32096 37564
rect 32032 37504 32096 37508
rect 32112 37564 32176 37568
rect 32112 37508 32116 37564
rect 32116 37508 32172 37564
rect 32172 37508 32176 37564
rect 32112 37504 32176 37508
rect 32192 37564 32256 37568
rect 32192 37508 32196 37564
rect 32196 37508 32252 37564
rect 32252 37508 32256 37564
rect 32192 37504 32256 37508
rect 36952 37564 37016 37568
rect 36952 37508 36956 37564
rect 36956 37508 37012 37564
rect 37012 37508 37016 37564
rect 36952 37504 37016 37508
rect 37032 37564 37096 37568
rect 37032 37508 37036 37564
rect 37036 37508 37092 37564
rect 37092 37508 37096 37564
rect 37032 37504 37096 37508
rect 37112 37564 37176 37568
rect 37112 37508 37116 37564
rect 37116 37508 37172 37564
rect 37172 37508 37176 37564
rect 37112 37504 37176 37508
rect 37192 37564 37256 37568
rect 37192 37508 37196 37564
rect 37196 37508 37252 37564
rect 37252 37508 37256 37564
rect 37192 37504 37256 37508
rect 2612 37020 2676 37024
rect 2612 36964 2616 37020
rect 2616 36964 2672 37020
rect 2672 36964 2676 37020
rect 2612 36960 2676 36964
rect 2692 37020 2756 37024
rect 2692 36964 2696 37020
rect 2696 36964 2752 37020
rect 2752 36964 2756 37020
rect 2692 36960 2756 36964
rect 2772 37020 2836 37024
rect 2772 36964 2776 37020
rect 2776 36964 2832 37020
rect 2832 36964 2836 37020
rect 2772 36960 2836 36964
rect 2852 37020 2916 37024
rect 2852 36964 2856 37020
rect 2856 36964 2912 37020
rect 2912 36964 2916 37020
rect 2852 36960 2916 36964
rect 7612 37020 7676 37024
rect 7612 36964 7616 37020
rect 7616 36964 7672 37020
rect 7672 36964 7676 37020
rect 7612 36960 7676 36964
rect 7692 37020 7756 37024
rect 7692 36964 7696 37020
rect 7696 36964 7752 37020
rect 7752 36964 7756 37020
rect 7692 36960 7756 36964
rect 7772 37020 7836 37024
rect 7772 36964 7776 37020
rect 7776 36964 7832 37020
rect 7832 36964 7836 37020
rect 7772 36960 7836 36964
rect 7852 37020 7916 37024
rect 7852 36964 7856 37020
rect 7856 36964 7912 37020
rect 7912 36964 7916 37020
rect 7852 36960 7916 36964
rect 12612 37020 12676 37024
rect 12612 36964 12616 37020
rect 12616 36964 12672 37020
rect 12672 36964 12676 37020
rect 12612 36960 12676 36964
rect 12692 37020 12756 37024
rect 12692 36964 12696 37020
rect 12696 36964 12752 37020
rect 12752 36964 12756 37020
rect 12692 36960 12756 36964
rect 12772 37020 12836 37024
rect 12772 36964 12776 37020
rect 12776 36964 12832 37020
rect 12832 36964 12836 37020
rect 12772 36960 12836 36964
rect 12852 37020 12916 37024
rect 12852 36964 12856 37020
rect 12856 36964 12912 37020
rect 12912 36964 12916 37020
rect 12852 36960 12916 36964
rect 17612 37020 17676 37024
rect 17612 36964 17616 37020
rect 17616 36964 17672 37020
rect 17672 36964 17676 37020
rect 17612 36960 17676 36964
rect 17692 37020 17756 37024
rect 17692 36964 17696 37020
rect 17696 36964 17752 37020
rect 17752 36964 17756 37020
rect 17692 36960 17756 36964
rect 17772 37020 17836 37024
rect 17772 36964 17776 37020
rect 17776 36964 17832 37020
rect 17832 36964 17836 37020
rect 17772 36960 17836 36964
rect 17852 37020 17916 37024
rect 17852 36964 17856 37020
rect 17856 36964 17912 37020
rect 17912 36964 17916 37020
rect 17852 36960 17916 36964
rect 22612 37020 22676 37024
rect 22612 36964 22616 37020
rect 22616 36964 22672 37020
rect 22672 36964 22676 37020
rect 22612 36960 22676 36964
rect 22692 37020 22756 37024
rect 22692 36964 22696 37020
rect 22696 36964 22752 37020
rect 22752 36964 22756 37020
rect 22692 36960 22756 36964
rect 22772 37020 22836 37024
rect 22772 36964 22776 37020
rect 22776 36964 22832 37020
rect 22832 36964 22836 37020
rect 22772 36960 22836 36964
rect 22852 37020 22916 37024
rect 22852 36964 22856 37020
rect 22856 36964 22912 37020
rect 22912 36964 22916 37020
rect 22852 36960 22916 36964
rect 27612 37020 27676 37024
rect 27612 36964 27616 37020
rect 27616 36964 27672 37020
rect 27672 36964 27676 37020
rect 27612 36960 27676 36964
rect 27692 37020 27756 37024
rect 27692 36964 27696 37020
rect 27696 36964 27752 37020
rect 27752 36964 27756 37020
rect 27692 36960 27756 36964
rect 27772 37020 27836 37024
rect 27772 36964 27776 37020
rect 27776 36964 27832 37020
rect 27832 36964 27836 37020
rect 27772 36960 27836 36964
rect 27852 37020 27916 37024
rect 27852 36964 27856 37020
rect 27856 36964 27912 37020
rect 27912 36964 27916 37020
rect 27852 36960 27916 36964
rect 32612 37020 32676 37024
rect 32612 36964 32616 37020
rect 32616 36964 32672 37020
rect 32672 36964 32676 37020
rect 32612 36960 32676 36964
rect 32692 37020 32756 37024
rect 32692 36964 32696 37020
rect 32696 36964 32752 37020
rect 32752 36964 32756 37020
rect 32692 36960 32756 36964
rect 32772 37020 32836 37024
rect 32772 36964 32776 37020
rect 32776 36964 32832 37020
rect 32832 36964 32836 37020
rect 32772 36960 32836 36964
rect 32852 37020 32916 37024
rect 32852 36964 32856 37020
rect 32856 36964 32912 37020
rect 32912 36964 32916 37020
rect 32852 36960 32916 36964
rect 37612 37020 37676 37024
rect 37612 36964 37616 37020
rect 37616 36964 37672 37020
rect 37672 36964 37676 37020
rect 37612 36960 37676 36964
rect 37692 37020 37756 37024
rect 37692 36964 37696 37020
rect 37696 36964 37752 37020
rect 37752 36964 37756 37020
rect 37692 36960 37756 36964
rect 37772 37020 37836 37024
rect 37772 36964 37776 37020
rect 37776 36964 37832 37020
rect 37832 36964 37836 37020
rect 37772 36960 37836 36964
rect 37852 37020 37916 37024
rect 37852 36964 37856 37020
rect 37856 36964 37912 37020
rect 37912 36964 37916 37020
rect 37852 36960 37916 36964
rect 1952 36476 2016 36480
rect 1952 36420 1956 36476
rect 1956 36420 2012 36476
rect 2012 36420 2016 36476
rect 1952 36416 2016 36420
rect 2032 36476 2096 36480
rect 2032 36420 2036 36476
rect 2036 36420 2092 36476
rect 2092 36420 2096 36476
rect 2032 36416 2096 36420
rect 2112 36476 2176 36480
rect 2112 36420 2116 36476
rect 2116 36420 2172 36476
rect 2172 36420 2176 36476
rect 2112 36416 2176 36420
rect 2192 36476 2256 36480
rect 2192 36420 2196 36476
rect 2196 36420 2252 36476
rect 2252 36420 2256 36476
rect 2192 36416 2256 36420
rect 6952 36476 7016 36480
rect 6952 36420 6956 36476
rect 6956 36420 7012 36476
rect 7012 36420 7016 36476
rect 6952 36416 7016 36420
rect 7032 36476 7096 36480
rect 7032 36420 7036 36476
rect 7036 36420 7092 36476
rect 7092 36420 7096 36476
rect 7032 36416 7096 36420
rect 7112 36476 7176 36480
rect 7112 36420 7116 36476
rect 7116 36420 7172 36476
rect 7172 36420 7176 36476
rect 7112 36416 7176 36420
rect 7192 36476 7256 36480
rect 7192 36420 7196 36476
rect 7196 36420 7252 36476
rect 7252 36420 7256 36476
rect 7192 36416 7256 36420
rect 11952 36476 12016 36480
rect 11952 36420 11956 36476
rect 11956 36420 12012 36476
rect 12012 36420 12016 36476
rect 11952 36416 12016 36420
rect 12032 36476 12096 36480
rect 12032 36420 12036 36476
rect 12036 36420 12092 36476
rect 12092 36420 12096 36476
rect 12032 36416 12096 36420
rect 12112 36476 12176 36480
rect 12112 36420 12116 36476
rect 12116 36420 12172 36476
rect 12172 36420 12176 36476
rect 12112 36416 12176 36420
rect 12192 36476 12256 36480
rect 12192 36420 12196 36476
rect 12196 36420 12252 36476
rect 12252 36420 12256 36476
rect 12192 36416 12256 36420
rect 16952 36476 17016 36480
rect 16952 36420 16956 36476
rect 16956 36420 17012 36476
rect 17012 36420 17016 36476
rect 16952 36416 17016 36420
rect 17032 36476 17096 36480
rect 17032 36420 17036 36476
rect 17036 36420 17092 36476
rect 17092 36420 17096 36476
rect 17032 36416 17096 36420
rect 17112 36476 17176 36480
rect 17112 36420 17116 36476
rect 17116 36420 17172 36476
rect 17172 36420 17176 36476
rect 17112 36416 17176 36420
rect 17192 36476 17256 36480
rect 17192 36420 17196 36476
rect 17196 36420 17252 36476
rect 17252 36420 17256 36476
rect 17192 36416 17256 36420
rect 21952 36476 22016 36480
rect 21952 36420 21956 36476
rect 21956 36420 22012 36476
rect 22012 36420 22016 36476
rect 21952 36416 22016 36420
rect 22032 36476 22096 36480
rect 22032 36420 22036 36476
rect 22036 36420 22092 36476
rect 22092 36420 22096 36476
rect 22032 36416 22096 36420
rect 22112 36476 22176 36480
rect 22112 36420 22116 36476
rect 22116 36420 22172 36476
rect 22172 36420 22176 36476
rect 22112 36416 22176 36420
rect 22192 36476 22256 36480
rect 22192 36420 22196 36476
rect 22196 36420 22252 36476
rect 22252 36420 22256 36476
rect 22192 36416 22256 36420
rect 26952 36476 27016 36480
rect 26952 36420 26956 36476
rect 26956 36420 27012 36476
rect 27012 36420 27016 36476
rect 26952 36416 27016 36420
rect 27032 36476 27096 36480
rect 27032 36420 27036 36476
rect 27036 36420 27092 36476
rect 27092 36420 27096 36476
rect 27032 36416 27096 36420
rect 27112 36476 27176 36480
rect 27112 36420 27116 36476
rect 27116 36420 27172 36476
rect 27172 36420 27176 36476
rect 27112 36416 27176 36420
rect 27192 36476 27256 36480
rect 27192 36420 27196 36476
rect 27196 36420 27252 36476
rect 27252 36420 27256 36476
rect 27192 36416 27256 36420
rect 31952 36476 32016 36480
rect 31952 36420 31956 36476
rect 31956 36420 32012 36476
rect 32012 36420 32016 36476
rect 31952 36416 32016 36420
rect 32032 36476 32096 36480
rect 32032 36420 32036 36476
rect 32036 36420 32092 36476
rect 32092 36420 32096 36476
rect 32032 36416 32096 36420
rect 32112 36476 32176 36480
rect 32112 36420 32116 36476
rect 32116 36420 32172 36476
rect 32172 36420 32176 36476
rect 32112 36416 32176 36420
rect 32192 36476 32256 36480
rect 32192 36420 32196 36476
rect 32196 36420 32252 36476
rect 32252 36420 32256 36476
rect 32192 36416 32256 36420
rect 36952 36476 37016 36480
rect 36952 36420 36956 36476
rect 36956 36420 37012 36476
rect 37012 36420 37016 36476
rect 36952 36416 37016 36420
rect 37032 36476 37096 36480
rect 37032 36420 37036 36476
rect 37036 36420 37092 36476
rect 37092 36420 37096 36476
rect 37032 36416 37096 36420
rect 37112 36476 37176 36480
rect 37112 36420 37116 36476
rect 37116 36420 37172 36476
rect 37172 36420 37176 36476
rect 37112 36416 37176 36420
rect 37192 36476 37256 36480
rect 37192 36420 37196 36476
rect 37196 36420 37252 36476
rect 37252 36420 37256 36476
rect 37192 36416 37256 36420
rect 18092 36076 18156 36140
rect 2612 35932 2676 35936
rect 2612 35876 2616 35932
rect 2616 35876 2672 35932
rect 2672 35876 2676 35932
rect 2612 35872 2676 35876
rect 2692 35932 2756 35936
rect 2692 35876 2696 35932
rect 2696 35876 2752 35932
rect 2752 35876 2756 35932
rect 2692 35872 2756 35876
rect 2772 35932 2836 35936
rect 2772 35876 2776 35932
rect 2776 35876 2832 35932
rect 2832 35876 2836 35932
rect 2772 35872 2836 35876
rect 2852 35932 2916 35936
rect 2852 35876 2856 35932
rect 2856 35876 2912 35932
rect 2912 35876 2916 35932
rect 2852 35872 2916 35876
rect 7612 35932 7676 35936
rect 7612 35876 7616 35932
rect 7616 35876 7672 35932
rect 7672 35876 7676 35932
rect 7612 35872 7676 35876
rect 7692 35932 7756 35936
rect 7692 35876 7696 35932
rect 7696 35876 7752 35932
rect 7752 35876 7756 35932
rect 7692 35872 7756 35876
rect 7772 35932 7836 35936
rect 7772 35876 7776 35932
rect 7776 35876 7832 35932
rect 7832 35876 7836 35932
rect 7772 35872 7836 35876
rect 7852 35932 7916 35936
rect 7852 35876 7856 35932
rect 7856 35876 7912 35932
rect 7912 35876 7916 35932
rect 7852 35872 7916 35876
rect 12612 35932 12676 35936
rect 12612 35876 12616 35932
rect 12616 35876 12672 35932
rect 12672 35876 12676 35932
rect 12612 35872 12676 35876
rect 12692 35932 12756 35936
rect 12692 35876 12696 35932
rect 12696 35876 12752 35932
rect 12752 35876 12756 35932
rect 12692 35872 12756 35876
rect 12772 35932 12836 35936
rect 12772 35876 12776 35932
rect 12776 35876 12832 35932
rect 12832 35876 12836 35932
rect 12772 35872 12836 35876
rect 12852 35932 12916 35936
rect 12852 35876 12856 35932
rect 12856 35876 12912 35932
rect 12912 35876 12916 35932
rect 12852 35872 12916 35876
rect 17612 35932 17676 35936
rect 17612 35876 17616 35932
rect 17616 35876 17672 35932
rect 17672 35876 17676 35932
rect 17612 35872 17676 35876
rect 17692 35932 17756 35936
rect 17692 35876 17696 35932
rect 17696 35876 17752 35932
rect 17752 35876 17756 35932
rect 17692 35872 17756 35876
rect 17772 35932 17836 35936
rect 17772 35876 17776 35932
rect 17776 35876 17832 35932
rect 17832 35876 17836 35932
rect 17772 35872 17836 35876
rect 17852 35932 17916 35936
rect 17852 35876 17856 35932
rect 17856 35876 17912 35932
rect 17912 35876 17916 35932
rect 17852 35872 17916 35876
rect 22612 35932 22676 35936
rect 22612 35876 22616 35932
rect 22616 35876 22672 35932
rect 22672 35876 22676 35932
rect 22612 35872 22676 35876
rect 22692 35932 22756 35936
rect 22692 35876 22696 35932
rect 22696 35876 22752 35932
rect 22752 35876 22756 35932
rect 22692 35872 22756 35876
rect 22772 35932 22836 35936
rect 22772 35876 22776 35932
rect 22776 35876 22832 35932
rect 22832 35876 22836 35932
rect 22772 35872 22836 35876
rect 22852 35932 22916 35936
rect 22852 35876 22856 35932
rect 22856 35876 22912 35932
rect 22912 35876 22916 35932
rect 22852 35872 22916 35876
rect 27612 35932 27676 35936
rect 27612 35876 27616 35932
rect 27616 35876 27672 35932
rect 27672 35876 27676 35932
rect 27612 35872 27676 35876
rect 27692 35932 27756 35936
rect 27692 35876 27696 35932
rect 27696 35876 27752 35932
rect 27752 35876 27756 35932
rect 27692 35872 27756 35876
rect 27772 35932 27836 35936
rect 27772 35876 27776 35932
rect 27776 35876 27832 35932
rect 27832 35876 27836 35932
rect 27772 35872 27836 35876
rect 27852 35932 27916 35936
rect 27852 35876 27856 35932
rect 27856 35876 27912 35932
rect 27912 35876 27916 35932
rect 27852 35872 27916 35876
rect 32612 35932 32676 35936
rect 32612 35876 32616 35932
rect 32616 35876 32672 35932
rect 32672 35876 32676 35932
rect 32612 35872 32676 35876
rect 32692 35932 32756 35936
rect 32692 35876 32696 35932
rect 32696 35876 32752 35932
rect 32752 35876 32756 35932
rect 32692 35872 32756 35876
rect 32772 35932 32836 35936
rect 32772 35876 32776 35932
rect 32776 35876 32832 35932
rect 32832 35876 32836 35932
rect 32772 35872 32836 35876
rect 32852 35932 32916 35936
rect 32852 35876 32856 35932
rect 32856 35876 32912 35932
rect 32912 35876 32916 35932
rect 32852 35872 32916 35876
rect 37612 35932 37676 35936
rect 37612 35876 37616 35932
rect 37616 35876 37672 35932
rect 37672 35876 37676 35932
rect 37612 35872 37676 35876
rect 37692 35932 37756 35936
rect 37692 35876 37696 35932
rect 37696 35876 37752 35932
rect 37752 35876 37756 35932
rect 37692 35872 37756 35876
rect 37772 35932 37836 35936
rect 37772 35876 37776 35932
rect 37776 35876 37832 35932
rect 37832 35876 37836 35932
rect 37772 35872 37836 35876
rect 37852 35932 37916 35936
rect 37852 35876 37856 35932
rect 37856 35876 37912 35932
rect 37912 35876 37916 35932
rect 37852 35872 37916 35876
rect 1952 35388 2016 35392
rect 1952 35332 1956 35388
rect 1956 35332 2012 35388
rect 2012 35332 2016 35388
rect 1952 35328 2016 35332
rect 2032 35388 2096 35392
rect 2032 35332 2036 35388
rect 2036 35332 2092 35388
rect 2092 35332 2096 35388
rect 2032 35328 2096 35332
rect 2112 35388 2176 35392
rect 2112 35332 2116 35388
rect 2116 35332 2172 35388
rect 2172 35332 2176 35388
rect 2112 35328 2176 35332
rect 2192 35388 2256 35392
rect 2192 35332 2196 35388
rect 2196 35332 2252 35388
rect 2252 35332 2256 35388
rect 2192 35328 2256 35332
rect 6952 35388 7016 35392
rect 6952 35332 6956 35388
rect 6956 35332 7012 35388
rect 7012 35332 7016 35388
rect 6952 35328 7016 35332
rect 7032 35388 7096 35392
rect 7032 35332 7036 35388
rect 7036 35332 7092 35388
rect 7092 35332 7096 35388
rect 7032 35328 7096 35332
rect 7112 35388 7176 35392
rect 7112 35332 7116 35388
rect 7116 35332 7172 35388
rect 7172 35332 7176 35388
rect 7112 35328 7176 35332
rect 7192 35388 7256 35392
rect 7192 35332 7196 35388
rect 7196 35332 7252 35388
rect 7252 35332 7256 35388
rect 7192 35328 7256 35332
rect 11952 35388 12016 35392
rect 11952 35332 11956 35388
rect 11956 35332 12012 35388
rect 12012 35332 12016 35388
rect 11952 35328 12016 35332
rect 12032 35388 12096 35392
rect 12032 35332 12036 35388
rect 12036 35332 12092 35388
rect 12092 35332 12096 35388
rect 12032 35328 12096 35332
rect 12112 35388 12176 35392
rect 12112 35332 12116 35388
rect 12116 35332 12172 35388
rect 12172 35332 12176 35388
rect 12112 35328 12176 35332
rect 12192 35388 12256 35392
rect 12192 35332 12196 35388
rect 12196 35332 12252 35388
rect 12252 35332 12256 35388
rect 12192 35328 12256 35332
rect 16952 35388 17016 35392
rect 16952 35332 16956 35388
rect 16956 35332 17012 35388
rect 17012 35332 17016 35388
rect 16952 35328 17016 35332
rect 17032 35388 17096 35392
rect 17032 35332 17036 35388
rect 17036 35332 17092 35388
rect 17092 35332 17096 35388
rect 17032 35328 17096 35332
rect 17112 35388 17176 35392
rect 17112 35332 17116 35388
rect 17116 35332 17172 35388
rect 17172 35332 17176 35388
rect 17112 35328 17176 35332
rect 17192 35388 17256 35392
rect 17192 35332 17196 35388
rect 17196 35332 17252 35388
rect 17252 35332 17256 35388
rect 17192 35328 17256 35332
rect 21952 35388 22016 35392
rect 21952 35332 21956 35388
rect 21956 35332 22012 35388
rect 22012 35332 22016 35388
rect 21952 35328 22016 35332
rect 22032 35388 22096 35392
rect 22032 35332 22036 35388
rect 22036 35332 22092 35388
rect 22092 35332 22096 35388
rect 22032 35328 22096 35332
rect 22112 35388 22176 35392
rect 22112 35332 22116 35388
rect 22116 35332 22172 35388
rect 22172 35332 22176 35388
rect 22112 35328 22176 35332
rect 22192 35388 22256 35392
rect 22192 35332 22196 35388
rect 22196 35332 22252 35388
rect 22252 35332 22256 35388
rect 22192 35328 22256 35332
rect 26952 35388 27016 35392
rect 26952 35332 26956 35388
rect 26956 35332 27012 35388
rect 27012 35332 27016 35388
rect 26952 35328 27016 35332
rect 27032 35388 27096 35392
rect 27032 35332 27036 35388
rect 27036 35332 27092 35388
rect 27092 35332 27096 35388
rect 27032 35328 27096 35332
rect 27112 35388 27176 35392
rect 27112 35332 27116 35388
rect 27116 35332 27172 35388
rect 27172 35332 27176 35388
rect 27112 35328 27176 35332
rect 27192 35388 27256 35392
rect 27192 35332 27196 35388
rect 27196 35332 27252 35388
rect 27252 35332 27256 35388
rect 27192 35328 27256 35332
rect 31952 35388 32016 35392
rect 31952 35332 31956 35388
rect 31956 35332 32012 35388
rect 32012 35332 32016 35388
rect 31952 35328 32016 35332
rect 32032 35388 32096 35392
rect 32032 35332 32036 35388
rect 32036 35332 32092 35388
rect 32092 35332 32096 35388
rect 32032 35328 32096 35332
rect 32112 35388 32176 35392
rect 32112 35332 32116 35388
rect 32116 35332 32172 35388
rect 32172 35332 32176 35388
rect 32112 35328 32176 35332
rect 32192 35388 32256 35392
rect 32192 35332 32196 35388
rect 32196 35332 32252 35388
rect 32252 35332 32256 35388
rect 32192 35328 32256 35332
rect 36952 35388 37016 35392
rect 36952 35332 36956 35388
rect 36956 35332 37012 35388
rect 37012 35332 37016 35388
rect 36952 35328 37016 35332
rect 37032 35388 37096 35392
rect 37032 35332 37036 35388
rect 37036 35332 37092 35388
rect 37092 35332 37096 35388
rect 37032 35328 37096 35332
rect 37112 35388 37176 35392
rect 37112 35332 37116 35388
rect 37116 35332 37172 35388
rect 37172 35332 37176 35388
rect 37112 35328 37176 35332
rect 37192 35388 37256 35392
rect 37192 35332 37196 35388
rect 37196 35332 37252 35388
rect 37252 35332 37256 35388
rect 37192 35328 37256 35332
rect 2612 34844 2676 34848
rect 2612 34788 2616 34844
rect 2616 34788 2672 34844
rect 2672 34788 2676 34844
rect 2612 34784 2676 34788
rect 2692 34844 2756 34848
rect 2692 34788 2696 34844
rect 2696 34788 2752 34844
rect 2752 34788 2756 34844
rect 2692 34784 2756 34788
rect 2772 34844 2836 34848
rect 2772 34788 2776 34844
rect 2776 34788 2832 34844
rect 2832 34788 2836 34844
rect 2772 34784 2836 34788
rect 2852 34844 2916 34848
rect 2852 34788 2856 34844
rect 2856 34788 2912 34844
rect 2912 34788 2916 34844
rect 2852 34784 2916 34788
rect 7612 34844 7676 34848
rect 7612 34788 7616 34844
rect 7616 34788 7672 34844
rect 7672 34788 7676 34844
rect 7612 34784 7676 34788
rect 7692 34844 7756 34848
rect 7692 34788 7696 34844
rect 7696 34788 7752 34844
rect 7752 34788 7756 34844
rect 7692 34784 7756 34788
rect 7772 34844 7836 34848
rect 7772 34788 7776 34844
rect 7776 34788 7832 34844
rect 7832 34788 7836 34844
rect 7772 34784 7836 34788
rect 7852 34844 7916 34848
rect 7852 34788 7856 34844
rect 7856 34788 7912 34844
rect 7912 34788 7916 34844
rect 7852 34784 7916 34788
rect 12612 34844 12676 34848
rect 12612 34788 12616 34844
rect 12616 34788 12672 34844
rect 12672 34788 12676 34844
rect 12612 34784 12676 34788
rect 12692 34844 12756 34848
rect 12692 34788 12696 34844
rect 12696 34788 12752 34844
rect 12752 34788 12756 34844
rect 12692 34784 12756 34788
rect 12772 34844 12836 34848
rect 12772 34788 12776 34844
rect 12776 34788 12832 34844
rect 12832 34788 12836 34844
rect 12772 34784 12836 34788
rect 12852 34844 12916 34848
rect 12852 34788 12856 34844
rect 12856 34788 12912 34844
rect 12912 34788 12916 34844
rect 12852 34784 12916 34788
rect 17612 34844 17676 34848
rect 17612 34788 17616 34844
rect 17616 34788 17672 34844
rect 17672 34788 17676 34844
rect 17612 34784 17676 34788
rect 17692 34844 17756 34848
rect 17692 34788 17696 34844
rect 17696 34788 17752 34844
rect 17752 34788 17756 34844
rect 17692 34784 17756 34788
rect 17772 34844 17836 34848
rect 17772 34788 17776 34844
rect 17776 34788 17832 34844
rect 17832 34788 17836 34844
rect 17772 34784 17836 34788
rect 17852 34844 17916 34848
rect 17852 34788 17856 34844
rect 17856 34788 17912 34844
rect 17912 34788 17916 34844
rect 17852 34784 17916 34788
rect 22612 34844 22676 34848
rect 22612 34788 22616 34844
rect 22616 34788 22672 34844
rect 22672 34788 22676 34844
rect 22612 34784 22676 34788
rect 22692 34844 22756 34848
rect 22692 34788 22696 34844
rect 22696 34788 22752 34844
rect 22752 34788 22756 34844
rect 22692 34784 22756 34788
rect 22772 34844 22836 34848
rect 22772 34788 22776 34844
rect 22776 34788 22832 34844
rect 22832 34788 22836 34844
rect 22772 34784 22836 34788
rect 22852 34844 22916 34848
rect 22852 34788 22856 34844
rect 22856 34788 22912 34844
rect 22912 34788 22916 34844
rect 22852 34784 22916 34788
rect 27612 34844 27676 34848
rect 27612 34788 27616 34844
rect 27616 34788 27672 34844
rect 27672 34788 27676 34844
rect 27612 34784 27676 34788
rect 27692 34844 27756 34848
rect 27692 34788 27696 34844
rect 27696 34788 27752 34844
rect 27752 34788 27756 34844
rect 27692 34784 27756 34788
rect 27772 34844 27836 34848
rect 27772 34788 27776 34844
rect 27776 34788 27832 34844
rect 27832 34788 27836 34844
rect 27772 34784 27836 34788
rect 27852 34844 27916 34848
rect 27852 34788 27856 34844
rect 27856 34788 27912 34844
rect 27912 34788 27916 34844
rect 27852 34784 27916 34788
rect 32612 34844 32676 34848
rect 32612 34788 32616 34844
rect 32616 34788 32672 34844
rect 32672 34788 32676 34844
rect 32612 34784 32676 34788
rect 32692 34844 32756 34848
rect 32692 34788 32696 34844
rect 32696 34788 32752 34844
rect 32752 34788 32756 34844
rect 32692 34784 32756 34788
rect 32772 34844 32836 34848
rect 32772 34788 32776 34844
rect 32776 34788 32832 34844
rect 32832 34788 32836 34844
rect 32772 34784 32836 34788
rect 32852 34844 32916 34848
rect 32852 34788 32856 34844
rect 32856 34788 32912 34844
rect 32912 34788 32916 34844
rect 32852 34784 32916 34788
rect 37612 34844 37676 34848
rect 37612 34788 37616 34844
rect 37616 34788 37672 34844
rect 37672 34788 37676 34844
rect 37612 34784 37676 34788
rect 37692 34844 37756 34848
rect 37692 34788 37696 34844
rect 37696 34788 37752 34844
rect 37752 34788 37756 34844
rect 37692 34784 37756 34788
rect 37772 34844 37836 34848
rect 37772 34788 37776 34844
rect 37776 34788 37832 34844
rect 37832 34788 37836 34844
rect 37772 34784 37836 34788
rect 37852 34844 37916 34848
rect 37852 34788 37856 34844
rect 37856 34788 37912 34844
rect 37912 34788 37916 34844
rect 37852 34784 37916 34788
rect 18092 34444 18156 34508
rect 1952 34300 2016 34304
rect 1952 34244 1956 34300
rect 1956 34244 2012 34300
rect 2012 34244 2016 34300
rect 1952 34240 2016 34244
rect 2032 34300 2096 34304
rect 2032 34244 2036 34300
rect 2036 34244 2092 34300
rect 2092 34244 2096 34300
rect 2032 34240 2096 34244
rect 2112 34300 2176 34304
rect 2112 34244 2116 34300
rect 2116 34244 2172 34300
rect 2172 34244 2176 34300
rect 2112 34240 2176 34244
rect 2192 34300 2256 34304
rect 2192 34244 2196 34300
rect 2196 34244 2252 34300
rect 2252 34244 2256 34300
rect 2192 34240 2256 34244
rect 6952 34300 7016 34304
rect 6952 34244 6956 34300
rect 6956 34244 7012 34300
rect 7012 34244 7016 34300
rect 6952 34240 7016 34244
rect 7032 34300 7096 34304
rect 7032 34244 7036 34300
rect 7036 34244 7092 34300
rect 7092 34244 7096 34300
rect 7032 34240 7096 34244
rect 7112 34300 7176 34304
rect 7112 34244 7116 34300
rect 7116 34244 7172 34300
rect 7172 34244 7176 34300
rect 7112 34240 7176 34244
rect 7192 34300 7256 34304
rect 7192 34244 7196 34300
rect 7196 34244 7252 34300
rect 7252 34244 7256 34300
rect 7192 34240 7256 34244
rect 11952 34300 12016 34304
rect 11952 34244 11956 34300
rect 11956 34244 12012 34300
rect 12012 34244 12016 34300
rect 11952 34240 12016 34244
rect 12032 34300 12096 34304
rect 12032 34244 12036 34300
rect 12036 34244 12092 34300
rect 12092 34244 12096 34300
rect 12032 34240 12096 34244
rect 12112 34300 12176 34304
rect 12112 34244 12116 34300
rect 12116 34244 12172 34300
rect 12172 34244 12176 34300
rect 12112 34240 12176 34244
rect 12192 34300 12256 34304
rect 12192 34244 12196 34300
rect 12196 34244 12252 34300
rect 12252 34244 12256 34300
rect 12192 34240 12256 34244
rect 16952 34300 17016 34304
rect 16952 34244 16956 34300
rect 16956 34244 17012 34300
rect 17012 34244 17016 34300
rect 16952 34240 17016 34244
rect 17032 34300 17096 34304
rect 17032 34244 17036 34300
rect 17036 34244 17092 34300
rect 17092 34244 17096 34300
rect 17032 34240 17096 34244
rect 17112 34300 17176 34304
rect 17112 34244 17116 34300
rect 17116 34244 17172 34300
rect 17172 34244 17176 34300
rect 17112 34240 17176 34244
rect 17192 34300 17256 34304
rect 17192 34244 17196 34300
rect 17196 34244 17252 34300
rect 17252 34244 17256 34300
rect 17192 34240 17256 34244
rect 21952 34300 22016 34304
rect 21952 34244 21956 34300
rect 21956 34244 22012 34300
rect 22012 34244 22016 34300
rect 21952 34240 22016 34244
rect 22032 34300 22096 34304
rect 22032 34244 22036 34300
rect 22036 34244 22092 34300
rect 22092 34244 22096 34300
rect 22032 34240 22096 34244
rect 22112 34300 22176 34304
rect 22112 34244 22116 34300
rect 22116 34244 22172 34300
rect 22172 34244 22176 34300
rect 22112 34240 22176 34244
rect 22192 34300 22256 34304
rect 22192 34244 22196 34300
rect 22196 34244 22252 34300
rect 22252 34244 22256 34300
rect 22192 34240 22256 34244
rect 26952 34300 27016 34304
rect 26952 34244 26956 34300
rect 26956 34244 27012 34300
rect 27012 34244 27016 34300
rect 26952 34240 27016 34244
rect 27032 34300 27096 34304
rect 27032 34244 27036 34300
rect 27036 34244 27092 34300
rect 27092 34244 27096 34300
rect 27032 34240 27096 34244
rect 27112 34300 27176 34304
rect 27112 34244 27116 34300
rect 27116 34244 27172 34300
rect 27172 34244 27176 34300
rect 27112 34240 27176 34244
rect 27192 34300 27256 34304
rect 27192 34244 27196 34300
rect 27196 34244 27252 34300
rect 27252 34244 27256 34300
rect 27192 34240 27256 34244
rect 31952 34300 32016 34304
rect 31952 34244 31956 34300
rect 31956 34244 32012 34300
rect 32012 34244 32016 34300
rect 31952 34240 32016 34244
rect 32032 34300 32096 34304
rect 32032 34244 32036 34300
rect 32036 34244 32092 34300
rect 32092 34244 32096 34300
rect 32032 34240 32096 34244
rect 32112 34300 32176 34304
rect 32112 34244 32116 34300
rect 32116 34244 32172 34300
rect 32172 34244 32176 34300
rect 32112 34240 32176 34244
rect 32192 34300 32256 34304
rect 32192 34244 32196 34300
rect 32196 34244 32252 34300
rect 32252 34244 32256 34300
rect 32192 34240 32256 34244
rect 36952 34300 37016 34304
rect 36952 34244 36956 34300
rect 36956 34244 37012 34300
rect 37012 34244 37016 34300
rect 36952 34240 37016 34244
rect 37032 34300 37096 34304
rect 37032 34244 37036 34300
rect 37036 34244 37092 34300
rect 37092 34244 37096 34300
rect 37032 34240 37096 34244
rect 37112 34300 37176 34304
rect 37112 34244 37116 34300
rect 37116 34244 37172 34300
rect 37172 34244 37176 34300
rect 37112 34240 37176 34244
rect 37192 34300 37256 34304
rect 37192 34244 37196 34300
rect 37196 34244 37252 34300
rect 37252 34244 37256 34300
rect 37192 34240 37256 34244
rect 21036 33824 21100 33828
rect 21036 33768 21086 33824
rect 21086 33768 21100 33824
rect 21036 33764 21100 33768
rect 2612 33756 2676 33760
rect 2612 33700 2616 33756
rect 2616 33700 2672 33756
rect 2672 33700 2676 33756
rect 2612 33696 2676 33700
rect 2692 33756 2756 33760
rect 2692 33700 2696 33756
rect 2696 33700 2752 33756
rect 2752 33700 2756 33756
rect 2692 33696 2756 33700
rect 2772 33756 2836 33760
rect 2772 33700 2776 33756
rect 2776 33700 2832 33756
rect 2832 33700 2836 33756
rect 2772 33696 2836 33700
rect 2852 33756 2916 33760
rect 2852 33700 2856 33756
rect 2856 33700 2912 33756
rect 2912 33700 2916 33756
rect 2852 33696 2916 33700
rect 7612 33756 7676 33760
rect 7612 33700 7616 33756
rect 7616 33700 7672 33756
rect 7672 33700 7676 33756
rect 7612 33696 7676 33700
rect 7692 33756 7756 33760
rect 7692 33700 7696 33756
rect 7696 33700 7752 33756
rect 7752 33700 7756 33756
rect 7692 33696 7756 33700
rect 7772 33756 7836 33760
rect 7772 33700 7776 33756
rect 7776 33700 7832 33756
rect 7832 33700 7836 33756
rect 7772 33696 7836 33700
rect 7852 33756 7916 33760
rect 7852 33700 7856 33756
rect 7856 33700 7912 33756
rect 7912 33700 7916 33756
rect 7852 33696 7916 33700
rect 12612 33756 12676 33760
rect 12612 33700 12616 33756
rect 12616 33700 12672 33756
rect 12672 33700 12676 33756
rect 12612 33696 12676 33700
rect 12692 33756 12756 33760
rect 12692 33700 12696 33756
rect 12696 33700 12752 33756
rect 12752 33700 12756 33756
rect 12692 33696 12756 33700
rect 12772 33756 12836 33760
rect 12772 33700 12776 33756
rect 12776 33700 12832 33756
rect 12832 33700 12836 33756
rect 12772 33696 12836 33700
rect 12852 33756 12916 33760
rect 12852 33700 12856 33756
rect 12856 33700 12912 33756
rect 12912 33700 12916 33756
rect 12852 33696 12916 33700
rect 17612 33756 17676 33760
rect 17612 33700 17616 33756
rect 17616 33700 17672 33756
rect 17672 33700 17676 33756
rect 17612 33696 17676 33700
rect 17692 33756 17756 33760
rect 17692 33700 17696 33756
rect 17696 33700 17752 33756
rect 17752 33700 17756 33756
rect 17692 33696 17756 33700
rect 17772 33756 17836 33760
rect 17772 33700 17776 33756
rect 17776 33700 17832 33756
rect 17832 33700 17836 33756
rect 17772 33696 17836 33700
rect 17852 33756 17916 33760
rect 17852 33700 17856 33756
rect 17856 33700 17912 33756
rect 17912 33700 17916 33756
rect 17852 33696 17916 33700
rect 22612 33756 22676 33760
rect 22612 33700 22616 33756
rect 22616 33700 22672 33756
rect 22672 33700 22676 33756
rect 22612 33696 22676 33700
rect 22692 33756 22756 33760
rect 22692 33700 22696 33756
rect 22696 33700 22752 33756
rect 22752 33700 22756 33756
rect 22692 33696 22756 33700
rect 22772 33756 22836 33760
rect 22772 33700 22776 33756
rect 22776 33700 22832 33756
rect 22832 33700 22836 33756
rect 22772 33696 22836 33700
rect 22852 33756 22916 33760
rect 22852 33700 22856 33756
rect 22856 33700 22912 33756
rect 22912 33700 22916 33756
rect 22852 33696 22916 33700
rect 27612 33756 27676 33760
rect 27612 33700 27616 33756
rect 27616 33700 27672 33756
rect 27672 33700 27676 33756
rect 27612 33696 27676 33700
rect 27692 33756 27756 33760
rect 27692 33700 27696 33756
rect 27696 33700 27752 33756
rect 27752 33700 27756 33756
rect 27692 33696 27756 33700
rect 27772 33756 27836 33760
rect 27772 33700 27776 33756
rect 27776 33700 27832 33756
rect 27832 33700 27836 33756
rect 27772 33696 27836 33700
rect 27852 33756 27916 33760
rect 27852 33700 27856 33756
rect 27856 33700 27912 33756
rect 27912 33700 27916 33756
rect 27852 33696 27916 33700
rect 32612 33756 32676 33760
rect 32612 33700 32616 33756
rect 32616 33700 32672 33756
rect 32672 33700 32676 33756
rect 32612 33696 32676 33700
rect 32692 33756 32756 33760
rect 32692 33700 32696 33756
rect 32696 33700 32752 33756
rect 32752 33700 32756 33756
rect 32692 33696 32756 33700
rect 32772 33756 32836 33760
rect 32772 33700 32776 33756
rect 32776 33700 32832 33756
rect 32832 33700 32836 33756
rect 32772 33696 32836 33700
rect 32852 33756 32916 33760
rect 32852 33700 32856 33756
rect 32856 33700 32912 33756
rect 32912 33700 32916 33756
rect 32852 33696 32916 33700
rect 37612 33756 37676 33760
rect 37612 33700 37616 33756
rect 37616 33700 37672 33756
rect 37672 33700 37676 33756
rect 37612 33696 37676 33700
rect 37692 33756 37756 33760
rect 37692 33700 37696 33756
rect 37696 33700 37752 33756
rect 37752 33700 37756 33756
rect 37692 33696 37756 33700
rect 37772 33756 37836 33760
rect 37772 33700 37776 33756
rect 37776 33700 37832 33756
rect 37832 33700 37836 33756
rect 37772 33696 37836 33700
rect 37852 33756 37916 33760
rect 37852 33700 37856 33756
rect 37856 33700 37912 33756
rect 37912 33700 37916 33756
rect 37852 33696 37916 33700
rect 1952 33212 2016 33216
rect 1952 33156 1956 33212
rect 1956 33156 2012 33212
rect 2012 33156 2016 33212
rect 1952 33152 2016 33156
rect 2032 33212 2096 33216
rect 2032 33156 2036 33212
rect 2036 33156 2092 33212
rect 2092 33156 2096 33212
rect 2032 33152 2096 33156
rect 2112 33212 2176 33216
rect 2112 33156 2116 33212
rect 2116 33156 2172 33212
rect 2172 33156 2176 33212
rect 2112 33152 2176 33156
rect 2192 33212 2256 33216
rect 2192 33156 2196 33212
rect 2196 33156 2252 33212
rect 2252 33156 2256 33212
rect 2192 33152 2256 33156
rect 6952 33212 7016 33216
rect 6952 33156 6956 33212
rect 6956 33156 7012 33212
rect 7012 33156 7016 33212
rect 6952 33152 7016 33156
rect 7032 33212 7096 33216
rect 7032 33156 7036 33212
rect 7036 33156 7092 33212
rect 7092 33156 7096 33212
rect 7032 33152 7096 33156
rect 7112 33212 7176 33216
rect 7112 33156 7116 33212
rect 7116 33156 7172 33212
rect 7172 33156 7176 33212
rect 7112 33152 7176 33156
rect 7192 33212 7256 33216
rect 7192 33156 7196 33212
rect 7196 33156 7252 33212
rect 7252 33156 7256 33212
rect 7192 33152 7256 33156
rect 11952 33212 12016 33216
rect 11952 33156 11956 33212
rect 11956 33156 12012 33212
rect 12012 33156 12016 33212
rect 11952 33152 12016 33156
rect 12032 33212 12096 33216
rect 12032 33156 12036 33212
rect 12036 33156 12092 33212
rect 12092 33156 12096 33212
rect 12032 33152 12096 33156
rect 12112 33212 12176 33216
rect 12112 33156 12116 33212
rect 12116 33156 12172 33212
rect 12172 33156 12176 33212
rect 12112 33152 12176 33156
rect 12192 33212 12256 33216
rect 12192 33156 12196 33212
rect 12196 33156 12252 33212
rect 12252 33156 12256 33212
rect 12192 33152 12256 33156
rect 16952 33212 17016 33216
rect 16952 33156 16956 33212
rect 16956 33156 17012 33212
rect 17012 33156 17016 33212
rect 16952 33152 17016 33156
rect 17032 33212 17096 33216
rect 17032 33156 17036 33212
rect 17036 33156 17092 33212
rect 17092 33156 17096 33212
rect 17032 33152 17096 33156
rect 17112 33212 17176 33216
rect 17112 33156 17116 33212
rect 17116 33156 17172 33212
rect 17172 33156 17176 33212
rect 17112 33152 17176 33156
rect 17192 33212 17256 33216
rect 17192 33156 17196 33212
rect 17196 33156 17252 33212
rect 17252 33156 17256 33212
rect 17192 33152 17256 33156
rect 21952 33212 22016 33216
rect 21952 33156 21956 33212
rect 21956 33156 22012 33212
rect 22012 33156 22016 33212
rect 21952 33152 22016 33156
rect 22032 33212 22096 33216
rect 22032 33156 22036 33212
rect 22036 33156 22092 33212
rect 22092 33156 22096 33212
rect 22032 33152 22096 33156
rect 22112 33212 22176 33216
rect 22112 33156 22116 33212
rect 22116 33156 22172 33212
rect 22172 33156 22176 33212
rect 22112 33152 22176 33156
rect 22192 33212 22256 33216
rect 22192 33156 22196 33212
rect 22196 33156 22252 33212
rect 22252 33156 22256 33212
rect 22192 33152 22256 33156
rect 26952 33212 27016 33216
rect 26952 33156 26956 33212
rect 26956 33156 27012 33212
rect 27012 33156 27016 33212
rect 26952 33152 27016 33156
rect 27032 33212 27096 33216
rect 27032 33156 27036 33212
rect 27036 33156 27092 33212
rect 27092 33156 27096 33212
rect 27032 33152 27096 33156
rect 27112 33212 27176 33216
rect 27112 33156 27116 33212
rect 27116 33156 27172 33212
rect 27172 33156 27176 33212
rect 27112 33152 27176 33156
rect 27192 33212 27256 33216
rect 27192 33156 27196 33212
rect 27196 33156 27252 33212
rect 27252 33156 27256 33212
rect 27192 33152 27256 33156
rect 31952 33212 32016 33216
rect 31952 33156 31956 33212
rect 31956 33156 32012 33212
rect 32012 33156 32016 33212
rect 31952 33152 32016 33156
rect 32032 33212 32096 33216
rect 32032 33156 32036 33212
rect 32036 33156 32092 33212
rect 32092 33156 32096 33212
rect 32032 33152 32096 33156
rect 32112 33212 32176 33216
rect 32112 33156 32116 33212
rect 32116 33156 32172 33212
rect 32172 33156 32176 33212
rect 32112 33152 32176 33156
rect 32192 33212 32256 33216
rect 32192 33156 32196 33212
rect 32196 33156 32252 33212
rect 32252 33156 32256 33212
rect 32192 33152 32256 33156
rect 36952 33212 37016 33216
rect 36952 33156 36956 33212
rect 36956 33156 37012 33212
rect 37012 33156 37016 33212
rect 36952 33152 37016 33156
rect 37032 33212 37096 33216
rect 37032 33156 37036 33212
rect 37036 33156 37092 33212
rect 37092 33156 37096 33212
rect 37032 33152 37096 33156
rect 37112 33212 37176 33216
rect 37112 33156 37116 33212
rect 37116 33156 37172 33212
rect 37172 33156 37176 33212
rect 37112 33152 37176 33156
rect 37192 33212 37256 33216
rect 37192 33156 37196 33212
rect 37196 33156 37252 33212
rect 37252 33156 37256 33212
rect 37192 33152 37256 33156
rect 2612 32668 2676 32672
rect 2612 32612 2616 32668
rect 2616 32612 2672 32668
rect 2672 32612 2676 32668
rect 2612 32608 2676 32612
rect 2692 32668 2756 32672
rect 2692 32612 2696 32668
rect 2696 32612 2752 32668
rect 2752 32612 2756 32668
rect 2692 32608 2756 32612
rect 2772 32668 2836 32672
rect 2772 32612 2776 32668
rect 2776 32612 2832 32668
rect 2832 32612 2836 32668
rect 2772 32608 2836 32612
rect 2852 32668 2916 32672
rect 2852 32612 2856 32668
rect 2856 32612 2912 32668
rect 2912 32612 2916 32668
rect 2852 32608 2916 32612
rect 7612 32668 7676 32672
rect 7612 32612 7616 32668
rect 7616 32612 7672 32668
rect 7672 32612 7676 32668
rect 7612 32608 7676 32612
rect 7692 32668 7756 32672
rect 7692 32612 7696 32668
rect 7696 32612 7752 32668
rect 7752 32612 7756 32668
rect 7692 32608 7756 32612
rect 7772 32668 7836 32672
rect 7772 32612 7776 32668
rect 7776 32612 7832 32668
rect 7832 32612 7836 32668
rect 7772 32608 7836 32612
rect 7852 32668 7916 32672
rect 7852 32612 7856 32668
rect 7856 32612 7912 32668
rect 7912 32612 7916 32668
rect 7852 32608 7916 32612
rect 12612 32668 12676 32672
rect 12612 32612 12616 32668
rect 12616 32612 12672 32668
rect 12672 32612 12676 32668
rect 12612 32608 12676 32612
rect 12692 32668 12756 32672
rect 12692 32612 12696 32668
rect 12696 32612 12752 32668
rect 12752 32612 12756 32668
rect 12692 32608 12756 32612
rect 12772 32668 12836 32672
rect 12772 32612 12776 32668
rect 12776 32612 12832 32668
rect 12832 32612 12836 32668
rect 12772 32608 12836 32612
rect 12852 32668 12916 32672
rect 12852 32612 12856 32668
rect 12856 32612 12912 32668
rect 12912 32612 12916 32668
rect 12852 32608 12916 32612
rect 17612 32668 17676 32672
rect 17612 32612 17616 32668
rect 17616 32612 17672 32668
rect 17672 32612 17676 32668
rect 17612 32608 17676 32612
rect 17692 32668 17756 32672
rect 17692 32612 17696 32668
rect 17696 32612 17752 32668
rect 17752 32612 17756 32668
rect 17692 32608 17756 32612
rect 17772 32668 17836 32672
rect 17772 32612 17776 32668
rect 17776 32612 17832 32668
rect 17832 32612 17836 32668
rect 17772 32608 17836 32612
rect 17852 32668 17916 32672
rect 17852 32612 17856 32668
rect 17856 32612 17912 32668
rect 17912 32612 17916 32668
rect 17852 32608 17916 32612
rect 22612 32668 22676 32672
rect 22612 32612 22616 32668
rect 22616 32612 22672 32668
rect 22672 32612 22676 32668
rect 22612 32608 22676 32612
rect 22692 32668 22756 32672
rect 22692 32612 22696 32668
rect 22696 32612 22752 32668
rect 22752 32612 22756 32668
rect 22692 32608 22756 32612
rect 22772 32668 22836 32672
rect 22772 32612 22776 32668
rect 22776 32612 22832 32668
rect 22832 32612 22836 32668
rect 22772 32608 22836 32612
rect 22852 32668 22916 32672
rect 22852 32612 22856 32668
rect 22856 32612 22912 32668
rect 22912 32612 22916 32668
rect 22852 32608 22916 32612
rect 27612 32668 27676 32672
rect 27612 32612 27616 32668
rect 27616 32612 27672 32668
rect 27672 32612 27676 32668
rect 27612 32608 27676 32612
rect 27692 32668 27756 32672
rect 27692 32612 27696 32668
rect 27696 32612 27752 32668
rect 27752 32612 27756 32668
rect 27692 32608 27756 32612
rect 27772 32668 27836 32672
rect 27772 32612 27776 32668
rect 27776 32612 27832 32668
rect 27832 32612 27836 32668
rect 27772 32608 27836 32612
rect 27852 32668 27916 32672
rect 27852 32612 27856 32668
rect 27856 32612 27912 32668
rect 27912 32612 27916 32668
rect 27852 32608 27916 32612
rect 32612 32668 32676 32672
rect 32612 32612 32616 32668
rect 32616 32612 32672 32668
rect 32672 32612 32676 32668
rect 32612 32608 32676 32612
rect 32692 32668 32756 32672
rect 32692 32612 32696 32668
rect 32696 32612 32752 32668
rect 32752 32612 32756 32668
rect 32692 32608 32756 32612
rect 32772 32668 32836 32672
rect 32772 32612 32776 32668
rect 32776 32612 32832 32668
rect 32832 32612 32836 32668
rect 32772 32608 32836 32612
rect 32852 32668 32916 32672
rect 32852 32612 32856 32668
rect 32856 32612 32912 32668
rect 32912 32612 32916 32668
rect 32852 32608 32916 32612
rect 37612 32668 37676 32672
rect 37612 32612 37616 32668
rect 37616 32612 37672 32668
rect 37672 32612 37676 32668
rect 37612 32608 37676 32612
rect 37692 32668 37756 32672
rect 37692 32612 37696 32668
rect 37696 32612 37752 32668
rect 37752 32612 37756 32668
rect 37692 32608 37756 32612
rect 37772 32668 37836 32672
rect 37772 32612 37776 32668
rect 37776 32612 37832 32668
rect 37832 32612 37836 32668
rect 37772 32608 37836 32612
rect 37852 32668 37916 32672
rect 37852 32612 37856 32668
rect 37856 32612 37912 32668
rect 37912 32612 37916 32668
rect 37852 32608 37916 32612
rect 1952 32124 2016 32128
rect 1952 32068 1956 32124
rect 1956 32068 2012 32124
rect 2012 32068 2016 32124
rect 1952 32064 2016 32068
rect 2032 32124 2096 32128
rect 2032 32068 2036 32124
rect 2036 32068 2092 32124
rect 2092 32068 2096 32124
rect 2032 32064 2096 32068
rect 2112 32124 2176 32128
rect 2112 32068 2116 32124
rect 2116 32068 2172 32124
rect 2172 32068 2176 32124
rect 2112 32064 2176 32068
rect 2192 32124 2256 32128
rect 2192 32068 2196 32124
rect 2196 32068 2252 32124
rect 2252 32068 2256 32124
rect 2192 32064 2256 32068
rect 6952 32124 7016 32128
rect 6952 32068 6956 32124
rect 6956 32068 7012 32124
rect 7012 32068 7016 32124
rect 6952 32064 7016 32068
rect 7032 32124 7096 32128
rect 7032 32068 7036 32124
rect 7036 32068 7092 32124
rect 7092 32068 7096 32124
rect 7032 32064 7096 32068
rect 7112 32124 7176 32128
rect 7112 32068 7116 32124
rect 7116 32068 7172 32124
rect 7172 32068 7176 32124
rect 7112 32064 7176 32068
rect 7192 32124 7256 32128
rect 7192 32068 7196 32124
rect 7196 32068 7252 32124
rect 7252 32068 7256 32124
rect 7192 32064 7256 32068
rect 11952 32124 12016 32128
rect 11952 32068 11956 32124
rect 11956 32068 12012 32124
rect 12012 32068 12016 32124
rect 11952 32064 12016 32068
rect 12032 32124 12096 32128
rect 12032 32068 12036 32124
rect 12036 32068 12092 32124
rect 12092 32068 12096 32124
rect 12032 32064 12096 32068
rect 12112 32124 12176 32128
rect 12112 32068 12116 32124
rect 12116 32068 12172 32124
rect 12172 32068 12176 32124
rect 12112 32064 12176 32068
rect 12192 32124 12256 32128
rect 12192 32068 12196 32124
rect 12196 32068 12252 32124
rect 12252 32068 12256 32124
rect 12192 32064 12256 32068
rect 16952 32124 17016 32128
rect 16952 32068 16956 32124
rect 16956 32068 17012 32124
rect 17012 32068 17016 32124
rect 16952 32064 17016 32068
rect 17032 32124 17096 32128
rect 17032 32068 17036 32124
rect 17036 32068 17092 32124
rect 17092 32068 17096 32124
rect 17032 32064 17096 32068
rect 17112 32124 17176 32128
rect 17112 32068 17116 32124
rect 17116 32068 17172 32124
rect 17172 32068 17176 32124
rect 17112 32064 17176 32068
rect 17192 32124 17256 32128
rect 17192 32068 17196 32124
rect 17196 32068 17252 32124
rect 17252 32068 17256 32124
rect 17192 32064 17256 32068
rect 21952 32124 22016 32128
rect 21952 32068 21956 32124
rect 21956 32068 22012 32124
rect 22012 32068 22016 32124
rect 21952 32064 22016 32068
rect 22032 32124 22096 32128
rect 22032 32068 22036 32124
rect 22036 32068 22092 32124
rect 22092 32068 22096 32124
rect 22032 32064 22096 32068
rect 22112 32124 22176 32128
rect 22112 32068 22116 32124
rect 22116 32068 22172 32124
rect 22172 32068 22176 32124
rect 22112 32064 22176 32068
rect 22192 32124 22256 32128
rect 22192 32068 22196 32124
rect 22196 32068 22252 32124
rect 22252 32068 22256 32124
rect 22192 32064 22256 32068
rect 26952 32124 27016 32128
rect 26952 32068 26956 32124
rect 26956 32068 27012 32124
rect 27012 32068 27016 32124
rect 26952 32064 27016 32068
rect 27032 32124 27096 32128
rect 27032 32068 27036 32124
rect 27036 32068 27092 32124
rect 27092 32068 27096 32124
rect 27032 32064 27096 32068
rect 27112 32124 27176 32128
rect 27112 32068 27116 32124
rect 27116 32068 27172 32124
rect 27172 32068 27176 32124
rect 27112 32064 27176 32068
rect 27192 32124 27256 32128
rect 27192 32068 27196 32124
rect 27196 32068 27252 32124
rect 27252 32068 27256 32124
rect 27192 32064 27256 32068
rect 31952 32124 32016 32128
rect 31952 32068 31956 32124
rect 31956 32068 32012 32124
rect 32012 32068 32016 32124
rect 31952 32064 32016 32068
rect 32032 32124 32096 32128
rect 32032 32068 32036 32124
rect 32036 32068 32092 32124
rect 32092 32068 32096 32124
rect 32032 32064 32096 32068
rect 32112 32124 32176 32128
rect 32112 32068 32116 32124
rect 32116 32068 32172 32124
rect 32172 32068 32176 32124
rect 32112 32064 32176 32068
rect 32192 32124 32256 32128
rect 32192 32068 32196 32124
rect 32196 32068 32252 32124
rect 32252 32068 32256 32124
rect 32192 32064 32256 32068
rect 36952 32124 37016 32128
rect 36952 32068 36956 32124
rect 36956 32068 37012 32124
rect 37012 32068 37016 32124
rect 36952 32064 37016 32068
rect 37032 32124 37096 32128
rect 37032 32068 37036 32124
rect 37036 32068 37092 32124
rect 37092 32068 37096 32124
rect 37032 32064 37096 32068
rect 37112 32124 37176 32128
rect 37112 32068 37116 32124
rect 37116 32068 37172 32124
rect 37172 32068 37176 32124
rect 37112 32064 37176 32068
rect 37192 32124 37256 32128
rect 37192 32068 37196 32124
rect 37196 32068 37252 32124
rect 37252 32068 37256 32124
rect 37192 32064 37256 32068
rect 2612 31580 2676 31584
rect 2612 31524 2616 31580
rect 2616 31524 2672 31580
rect 2672 31524 2676 31580
rect 2612 31520 2676 31524
rect 2692 31580 2756 31584
rect 2692 31524 2696 31580
rect 2696 31524 2752 31580
rect 2752 31524 2756 31580
rect 2692 31520 2756 31524
rect 2772 31580 2836 31584
rect 2772 31524 2776 31580
rect 2776 31524 2832 31580
rect 2832 31524 2836 31580
rect 2772 31520 2836 31524
rect 2852 31580 2916 31584
rect 2852 31524 2856 31580
rect 2856 31524 2912 31580
rect 2912 31524 2916 31580
rect 2852 31520 2916 31524
rect 7612 31580 7676 31584
rect 7612 31524 7616 31580
rect 7616 31524 7672 31580
rect 7672 31524 7676 31580
rect 7612 31520 7676 31524
rect 7692 31580 7756 31584
rect 7692 31524 7696 31580
rect 7696 31524 7752 31580
rect 7752 31524 7756 31580
rect 7692 31520 7756 31524
rect 7772 31580 7836 31584
rect 7772 31524 7776 31580
rect 7776 31524 7832 31580
rect 7832 31524 7836 31580
rect 7772 31520 7836 31524
rect 7852 31580 7916 31584
rect 7852 31524 7856 31580
rect 7856 31524 7912 31580
rect 7912 31524 7916 31580
rect 7852 31520 7916 31524
rect 12612 31580 12676 31584
rect 12612 31524 12616 31580
rect 12616 31524 12672 31580
rect 12672 31524 12676 31580
rect 12612 31520 12676 31524
rect 12692 31580 12756 31584
rect 12692 31524 12696 31580
rect 12696 31524 12752 31580
rect 12752 31524 12756 31580
rect 12692 31520 12756 31524
rect 12772 31580 12836 31584
rect 12772 31524 12776 31580
rect 12776 31524 12832 31580
rect 12832 31524 12836 31580
rect 12772 31520 12836 31524
rect 12852 31580 12916 31584
rect 12852 31524 12856 31580
rect 12856 31524 12912 31580
rect 12912 31524 12916 31580
rect 12852 31520 12916 31524
rect 17612 31580 17676 31584
rect 17612 31524 17616 31580
rect 17616 31524 17672 31580
rect 17672 31524 17676 31580
rect 17612 31520 17676 31524
rect 17692 31580 17756 31584
rect 17692 31524 17696 31580
rect 17696 31524 17752 31580
rect 17752 31524 17756 31580
rect 17692 31520 17756 31524
rect 17772 31580 17836 31584
rect 17772 31524 17776 31580
rect 17776 31524 17832 31580
rect 17832 31524 17836 31580
rect 17772 31520 17836 31524
rect 17852 31580 17916 31584
rect 17852 31524 17856 31580
rect 17856 31524 17912 31580
rect 17912 31524 17916 31580
rect 17852 31520 17916 31524
rect 22612 31580 22676 31584
rect 22612 31524 22616 31580
rect 22616 31524 22672 31580
rect 22672 31524 22676 31580
rect 22612 31520 22676 31524
rect 22692 31580 22756 31584
rect 22692 31524 22696 31580
rect 22696 31524 22752 31580
rect 22752 31524 22756 31580
rect 22692 31520 22756 31524
rect 22772 31580 22836 31584
rect 22772 31524 22776 31580
rect 22776 31524 22832 31580
rect 22832 31524 22836 31580
rect 22772 31520 22836 31524
rect 22852 31580 22916 31584
rect 22852 31524 22856 31580
rect 22856 31524 22912 31580
rect 22912 31524 22916 31580
rect 22852 31520 22916 31524
rect 27612 31580 27676 31584
rect 27612 31524 27616 31580
rect 27616 31524 27672 31580
rect 27672 31524 27676 31580
rect 27612 31520 27676 31524
rect 27692 31580 27756 31584
rect 27692 31524 27696 31580
rect 27696 31524 27752 31580
rect 27752 31524 27756 31580
rect 27692 31520 27756 31524
rect 27772 31580 27836 31584
rect 27772 31524 27776 31580
rect 27776 31524 27832 31580
rect 27832 31524 27836 31580
rect 27772 31520 27836 31524
rect 27852 31580 27916 31584
rect 27852 31524 27856 31580
rect 27856 31524 27912 31580
rect 27912 31524 27916 31580
rect 27852 31520 27916 31524
rect 32612 31580 32676 31584
rect 32612 31524 32616 31580
rect 32616 31524 32672 31580
rect 32672 31524 32676 31580
rect 32612 31520 32676 31524
rect 32692 31580 32756 31584
rect 32692 31524 32696 31580
rect 32696 31524 32752 31580
rect 32752 31524 32756 31580
rect 32692 31520 32756 31524
rect 32772 31580 32836 31584
rect 32772 31524 32776 31580
rect 32776 31524 32832 31580
rect 32832 31524 32836 31580
rect 32772 31520 32836 31524
rect 32852 31580 32916 31584
rect 32852 31524 32856 31580
rect 32856 31524 32912 31580
rect 32912 31524 32916 31580
rect 32852 31520 32916 31524
rect 37612 31580 37676 31584
rect 37612 31524 37616 31580
rect 37616 31524 37672 31580
rect 37672 31524 37676 31580
rect 37612 31520 37676 31524
rect 37692 31580 37756 31584
rect 37692 31524 37696 31580
rect 37696 31524 37752 31580
rect 37752 31524 37756 31580
rect 37692 31520 37756 31524
rect 37772 31580 37836 31584
rect 37772 31524 37776 31580
rect 37776 31524 37832 31580
rect 37832 31524 37836 31580
rect 37772 31520 37836 31524
rect 37852 31580 37916 31584
rect 37852 31524 37856 31580
rect 37856 31524 37912 31580
rect 37912 31524 37916 31580
rect 37852 31520 37916 31524
rect 1952 31036 2016 31040
rect 1952 30980 1956 31036
rect 1956 30980 2012 31036
rect 2012 30980 2016 31036
rect 1952 30976 2016 30980
rect 2032 31036 2096 31040
rect 2032 30980 2036 31036
rect 2036 30980 2092 31036
rect 2092 30980 2096 31036
rect 2032 30976 2096 30980
rect 2112 31036 2176 31040
rect 2112 30980 2116 31036
rect 2116 30980 2172 31036
rect 2172 30980 2176 31036
rect 2112 30976 2176 30980
rect 2192 31036 2256 31040
rect 2192 30980 2196 31036
rect 2196 30980 2252 31036
rect 2252 30980 2256 31036
rect 2192 30976 2256 30980
rect 6952 31036 7016 31040
rect 6952 30980 6956 31036
rect 6956 30980 7012 31036
rect 7012 30980 7016 31036
rect 6952 30976 7016 30980
rect 7032 31036 7096 31040
rect 7032 30980 7036 31036
rect 7036 30980 7092 31036
rect 7092 30980 7096 31036
rect 7032 30976 7096 30980
rect 7112 31036 7176 31040
rect 7112 30980 7116 31036
rect 7116 30980 7172 31036
rect 7172 30980 7176 31036
rect 7112 30976 7176 30980
rect 7192 31036 7256 31040
rect 7192 30980 7196 31036
rect 7196 30980 7252 31036
rect 7252 30980 7256 31036
rect 7192 30976 7256 30980
rect 11952 31036 12016 31040
rect 11952 30980 11956 31036
rect 11956 30980 12012 31036
rect 12012 30980 12016 31036
rect 11952 30976 12016 30980
rect 12032 31036 12096 31040
rect 12032 30980 12036 31036
rect 12036 30980 12092 31036
rect 12092 30980 12096 31036
rect 12032 30976 12096 30980
rect 12112 31036 12176 31040
rect 12112 30980 12116 31036
rect 12116 30980 12172 31036
rect 12172 30980 12176 31036
rect 12112 30976 12176 30980
rect 12192 31036 12256 31040
rect 12192 30980 12196 31036
rect 12196 30980 12252 31036
rect 12252 30980 12256 31036
rect 12192 30976 12256 30980
rect 16952 31036 17016 31040
rect 16952 30980 16956 31036
rect 16956 30980 17012 31036
rect 17012 30980 17016 31036
rect 16952 30976 17016 30980
rect 17032 31036 17096 31040
rect 17032 30980 17036 31036
rect 17036 30980 17092 31036
rect 17092 30980 17096 31036
rect 17032 30976 17096 30980
rect 17112 31036 17176 31040
rect 17112 30980 17116 31036
rect 17116 30980 17172 31036
rect 17172 30980 17176 31036
rect 17112 30976 17176 30980
rect 17192 31036 17256 31040
rect 17192 30980 17196 31036
rect 17196 30980 17252 31036
rect 17252 30980 17256 31036
rect 17192 30976 17256 30980
rect 21952 31036 22016 31040
rect 21952 30980 21956 31036
rect 21956 30980 22012 31036
rect 22012 30980 22016 31036
rect 21952 30976 22016 30980
rect 22032 31036 22096 31040
rect 22032 30980 22036 31036
rect 22036 30980 22092 31036
rect 22092 30980 22096 31036
rect 22032 30976 22096 30980
rect 22112 31036 22176 31040
rect 22112 30980 22116 31036
rect 22116 30980 22172 31036
rect 22172 30980 22176 31036
rect 22112 30976 22176 30980
rect 22192 31036 22256 31040
rect 22192 30980 22196 31036
rect 22196 30980 22252 31036
rect 22252 30980 22256 31036
rect 22192 30976 22256 30980
rect 26952 31036 27016 31040
rect 26952 30980 26956 31036
rect 26956 30980 27012 31036
rect 27012 30980 27016 31036
rect 26952 30976 27016 30980
rect 27032 31036 27096 31040
rect 27032 30980 27036 31036
rect 27036 30980 27092 31036
rect 27092 30980 27096 31036
rect 27032 30976 27096 30980
rect 27112 31036 27176 31040
rect 27112 30980 27116 31036
rect 27116 30980 27172 31036
rect 27172 30980 27176 31036
rect 27112 30976 27176 30980
rect 27192 31036 27256 31040
rect 27192 30980 27196 31036
rect 27196 30980 27252 31036
rect 27252 30980 27256 31036
rect 27192 30976 27256 30980
rect 31952 31036 32016 31040
rect 31952 30980 31956 31036
rect 31956 30980 32012 31036
rect 32012 30980 32016 31036
rect 31952 30976 32016 30980
rect 32032 31036 32096 31040
rect 32032 30980 32036 31036
rect 32036 30980 32092 31036
rect 32092 30980 32096 31036
rect 32032 30976 32096 30980
rect 32112 31036 32176 31040
rect 32112 30980 32116 31036
rect 32116 30980 32172 31036
rect 32172 30980 32176 31036
rect 32112 30976 32176 30980
rect 32192 31036 32256 31040
rect 32192 30980 32196 31036
rect 32196 30980 32252 31036
rect 32252 30980 32256 31036
rect 32192 30976 32256 30980
rect 36952 31036 37016 31040
rect 36952 30980 36956 31036
rect 36956 30980 37012 31036
rect 37012 30980 37016 31036
rect 36952 30976 37016 30980
rect 37032 31036 37096 31040
rect 37032 30980 37036 31036
rect 37036 30980 37092 31036
rect 37092 30980 37096 31036
rect 37032 30976 37096 30980
rect 37112 31036 37176 31040
rect 37112 30980 37116 31036
rect 37116 30980 37172 31036
rect 37172 30980 37176 31036
rect 37112 30976 37176 30980
rect 37192 31036 37256 31040
rect 37192 30980 37196 31036
rect 37196 30980 37252 31036
rect 37252 30980 37256 31036
rect 37192 30976 37256 30980
rect 2612 30492 2676 30496
rect 2612 30436 2616 30492
rect 2616 30436 2672 30492
rect 2672 30436 2676 30492
rect 2612 30432 2676 30436
rect 2692 30492 2756 30496
rect 2692 30436 2696 30492
rect 2696 30436 2752 30492
rect 2752 30436 2756 30492
rect 2692 30432 2756 30436
rect 2772 30492 2836 30496
rect 2772 30436 2776 30492
rect 2776 30436 2832 30492
rect 2832 30436 2836 30492
rect 2772 30432 2836 30436
rect 2852 30492 2916 30496
rect 2852 30436 2856 30492
rect 2856 30436 2912 30492
rect 2912 30436 2916 30492
rect 2852 30432 2916 30436
rect 7612 30492 7676 30496
rect 7612 30436 7616 30492
rect 7616 30436 7672 30492
rect 7672 30436 7676 30492
rect 7612 30432 7676 30436
rect 7692 30492 7756 30496
rect 7692 30436 7696 30492
rect 7696 30436 7752 30492
rect 7752 30436 7756 30492
rect 7692 30432 7756 30436
rect 7772 30492 7836 30496
rect 7772 30436 7776 30492
rect 7776 30436 7832 30492
rect 7832 30436 7836 30492
rect 7772 30432 7836 30436
rect 7852 30492 7916 30496
rect 7852 30436 7856 30492
rect 7856 30436 7912 30492
rect 7912 30436 7916 30492
rect 7852 30432 7916 30436
rect 12612 30492 12676 30496
rect 12612 30436 12616 30492
rect 12616 30436 12672 30492
rect 12672 30436 12676 30492
rect 12612 30432 12676 30436
rect 12692 30492 12756 30496
rect 12692 30436 12696 30492
rect 12696 30436 12752 30492
rect 12752 30436 12756 30492
rect 12692 30432 12756 30436
rect 12772 30492 12836 30496
rect 12772 30436 12776 30492
rect 12776 30436 12832 30492
rect 12832 30436 12836 30492
rect 12772 30432 12836 30436
rect 12852 30492 12916 30496
rect 12852 30436 12856 30492
rect 12856 30436 12912 30492
rect 12912 30436 12916 30492
rect 12852 30432 12916 30436
rect 17612 30492 17676 30496
rect 17612 30436 17616 30492
rect 17616 30436 17672 30492
rect 17672 30436 17676 30492
rect 17612 30432 17676 30436
rect 17692 30492 17756 30496
rect 17692 30436 17696 30492
rect 17696 30436 17752 30492
rect 17752 30436 17756 30492
rect 17692 30432 17756 30436
rect 17772 30492 17836 30496
rect 17772 30436 17776 30492
rect 17776 30436 17832 30492
rect 17832 30436 17836 30492
rect 17772 30432 17836 30436
rect 17852 30492 17916 30496
rect 17852 30436 17856 30492
rect 17856 30436 17912 30492
rect 17912 30436 17916 30492
rect 17852 30432 17916 30436
rect 22612 30492 22676 30496
rect 22612 30436 22616 30492
rect 22616 30436 22672 30492
rect 22672 30436 22676 30492
rect 22612 30432 22676 30436
rect 22692 30492 22756 30496
rect 22692 30436 22696 30492
rect 22696 30436 22752 30492
rect 22752 30436 22756 30492
rect 22692 30432 22756 30436
rect 22772 30492 22836 30496
rect 22772 30436 22776 30492
rect 22776 30436 22832 30492
rect 22832 30436 22836 30492
rect 22772 30432 22836 30436
rect 22852 30492 22916 30496
rect 22852 30436 22856 30492
rect 22856 30436 22912 30492
rect 22912 30436 22916 30492
rect 22852 30432 22916 30436
rect 27612 30492 27676 30496
rect 27612 30436 27616 30492
rect 27616 30436 27672 30492
rect 27672 30436 27676 30492
rect 27612 30432 27676 30436
rect 27692 30492 27756 30496
rect 27692 30436 27696 30492
rect 27696 30436 27752 30492
rect 27752 30436 27756 30492
rect 27692 30432 27756 30436
rect 27772 30492 27836 30496
rect 27772 30436 27776 30492
rect 27776 30436 27832 30492
rect 27832 30436 27836 30492
rect 27772 30432 27836 30436
rect 27852 30492 27916 30496
rect 27852 30436 27856 30492
rect 27856 30436 27912 30492
rect 27912 30436 27916 30492
rect 27852 30432 27916 30436
rect 32612 30492 32676 30496
rect 32612 30436 32616 30492
rect 32616 30436 32672 30492
rect 32672 30436 32676 30492
rect 32612 30432 32676 30436
rect 32692 30492 32756 30496
rect 32692 30436 32696 30492
rect 32696 30436 32752 30492
rect 32752 30436 32756 30492
rect 32692 30432 32756 30436
rect 32772 30492 32836 30496
rect 32772 30436 32776 30492
rect 32776 30436 32832 30492
rect 32832 30436 32836 30492
rect 32772 30432 32836 30436
rect 32852 30492 32916 30496
rect 32852 30436 32856 30492
rect 32856 30436 32912 30492
rect 32912 30436 32916 30492
rect 32852 30432 32916 30436
rect 37612 30492 37676 30496
rect 37612 30436 37616 30492
rect 37616 30436 37672 30492
rect 37672 30436 37676 30492
rect 37612 30432 37676 30436
rect 37692 30492 37756 30496
rect 37692 30436 37696 30492
rect 37696 30436 37752 30492
rect 37752 30436 37756 30492
rect 37692 30432 37756 30436
rect 37772 30492 37836 30496
rect 37772 30436 37776 30492
rect 37776 30436 37832 30492
rect 37832 30436 37836 30492
rect 37772 30432 37836 30436
rect 37852 30492 37916 30496
rect 37852 30436 37856 30492
rect 37856 30436 37912 30492
rect 37912 30436 37916 30492
rect 37852 30432 37916 30436
rect 1952 29948 2016 29952
rect 1952 29892 1956 29948
rect 1956 29892 2012 29948
rect 2012 29892 2016 29948
rect 1952 29888 2016 29892
rect 2032 29948 2096 29952
rect 2032 29892 2036 29948
rect 2036 29892 2092 29948
rect 2092 29892 2096 29948
rect 2032 29888 2096 29892
rect 2112 29948 2176 29952
rect 2112 29892 2116 29948
rect 2116 29892 2172 29948
rect 2172 29892 2176 29948
rect 2112 29888 2176 29892
rect 2192 29948 2256 29952
rect 2192 29892 2196 29948
rect 2196 29892 2252 29948
rect 2252 29892 2256 29948
rect 2192 29888 2256 29892
rect 6952 29948 7016 29952
rect 6952 29892 6956 29948
rect 6956 29892 7012 29948
rect 7012 29892 7016 29948
rect 6952 29888 7016 29892
rect 7032 29948 7096 29952
rect 7032 29892 7036 29948
rect 7036 29892 7092 29948
rect 7092 29892 7096 29948
rect 7032 29888 7096 29892
rect 7112 29948 7176 29952
rect 7112 29892 7116 29948
rect 7116 29892 7172 29948
rect 7172 29892 7176 29948
rect 7112 29888 7176 29892
rect 7192 29948 7256 29952
rect 7192 29892 7196 29948
rect 7196 29892 7252 29948
rect 7252 29892 7256 29948
rect 7192 29888 7256 29892
rect 11952 29948 12016 29952
rect 11952 29892 11956 29948
rect 11956 29892 12012 29948
rect 12012 29892 12016 29948
rect 11952 29888 12016 29892
rect 12032 29948 12096 29952
rect 12032 29892 12036 29948
rect 12036 29892 12092 29948
rect 12092 29892 12096 29948
rect 12032 29888 12096 29892
rect 12112 29948 12176 29952
rect 12112 29892 12116 29948
rect 12116 29892 12172 29948
rect 12172 29892 12176 29948
rect 12112 29888 12176 29892
rect 12192 29948 12256 29952
rect 12192 29892 12196 29948
rect 12196 29892 12252 29948
rect 12252 29892 12256 29948
rect 12192 29888 12256 29892
rect 16952 29948 17016 29952
rect 16952 29892 16956 29948
rect 16956 29892 17012 29948
rect 17012 29892 17016 29948
rect 16952 29888 17016 29892
rect 17032 29948 17096 29952
rect 17032 29892 17036 29948
rect 17036 29892 17092 29948
rect 17092 29892 17096 29948
rect 17032 29888 17096 29892
rect 17112 29948 17176 29952
rect 17112 29892 17116 29948
rect 17116 29892 17172 29948
rect 17172 29892 17176 29948
rect 17112 29888 17176 29892
rect 17192 29948 17256 29952
rect 17192 29892 17196 29948
rect 17196 29892 17252 29948
rect 17252 29892 17256 29948
rect 17192 29888 17256 29892
rect 21952 29948 22016 29952
rect 21952 29892 21956 29948
rect 21956 29892 22012 29948
rect 22012 29892 22016 29948
rect 21952 29888 22016 29892
rect 22032 29948 22096 29952
rect 22032 29892 22036 29948
rect 22036 29892 22092 29948
rect 22092 29892 22096 29948
rect 22032 29888 22096 29892
rect 22112 29948 22176 29952
rect 22112 29892 22116 29948
rect 22116 29892 22172 29948
rect 22172 29892 22176 29948
rect 22112 29888 22176 29892
rect 22192 29948 22256 29952
rect 22192 29892 22196 29948
rect 22196 29892 22252 29948
rect 22252 29892 22256 29948
rect 22192 29888 22256 29892
rect 26952 29948 27016 29952
rect 26952 29892 26956 29948
rect 26956 29892 27012 29948
rect 27012 29892 27016 29948
rect 26952 29888 27016 29892
rect 27032 29948 27096 29952
rect 27032 29892 27036 29948
rect 27036 29892 27092 29948
rect 27092 29892 27096 29948
rect 27032 29888 27096 29892
rect 27112 29948 27176 29952
rect 27112 29892 27116 29948
rect 27116 29892 27172 29948
rect 27172 29892 27176 29948
rect 27112 29888 27176 29892
rect 27192 29948 27256 29952
rect 27192 29892 27196 29948
rect 27196 29892 27252 29948
rect 27252 29892 27256 29948
rect 27192 29888 27256 29892
rect 31952 29948 32016 29952
rect 31952 29892 31956 29948
rect 31956 29892 32012 29948
rect 32012 29892 32016 29948
rect 31952 29888 32016 29892
rect 32032 29948 32096 29952
rect 32032 29892 32036 29948
rect 32036 29892 32092 29948
rect 32092 29892 32096 29948
rect 32032 29888 32096 29892
rect 32112 29948 32176 29952
rect 32112 29892 32116 29948
rect 32116 29892 32172 29948
rect 32172 29892 32176 29948
rect 32112 29888 32176 29892
rect 32192 29948 32256 29952
rect 32192 29892 32196 29948
rect 32196 29892 32252 29948
rect 32252 29892 32256 29948
rect 32192 29888 32256 29892
rect 36952 29948 37016 29952
rect 36952 29892 36956 29948
rect 36956 29892 37012 29948
rect 37012 29892 37016 29948
rect 36952 29888 37016 29892
rect 37032 29948 37096 29952
rect 37032 29892 37036 29948
rect 37036 29892 37092 29948
rect 37092 29892 37096 29948
rect 37032 29888 37096 29892
rect 37112 29948 37176 29952
rect 37112 29892 37116 29948
rect 37116 29892 37172 29948
rect 37172 29892 37176 29948
rect 37112 29888 37176 29892
rect 37192 29948 37256 29952
rect 37192 29892 37196 29948
rect 37196 29892 37252 29948
rect 37252 29892 37256 29948
rect 37192 29888 37256 29892
rect 2612 29404 2676 29408
rect 2612 29348 2616 29404
rect 2616 29348 2672 29404
rect 2672 29348 2676 29404
rect 2612 29344 2676 29348
rect 2692 29404 2756 29408
rect 2692 29348 2696 29404
rect 2696 29348 2752 29404
rect 2752 29348 2756 29404
rect 2692 29344 2756 29348
rect 2772 29404 2836 29408
rect 2772 29348 2776 29404
rect 2776 29348 2832 29404
rect 2832 29348 2836 29404
rect 2772 29344 2836 29348
rect 2852 29404 2916 29408
rect 2852 29348 2856 29404
rect 2856 29348 2912 29404
rect 2912 29348 2916 29404
rect 2852 29344 2916 29348
rect 7612 29404 7676 29408
rect 7612 29348 7616 29404
rect 7616 29348 7672 29404
rect 7672 29348 7676 29404
rect 7612 29344 7676 29348
rect 7692 29404 7756 29408
rect 7692 29348 7696 29404
rect 7696 29348 7752 29404
rect 7752 29348 7756 29404
rect 7692 29344 7756 29348
rect 7772 29404 7836 29408
rect 7772 29348 7776 29404
rect 7776 29348 7832 29404
rect 7832 29348 7836 29404
rect 7772 29344 7836 29348
rect 7852 29404 7916 29408
rect 7852 29348 7856 29404
rect 7856 29348 7912 29404
rect 7912 29348 7916 29404
rect 7852 29344 7916 29348
rect 12612 29404 12676 29408
rect 12612 29348 12616 29404
rect 12616 29348 12672 29404
rect 12672 29348 12676 29404
rect 12612 29344 12676 29348
rect 12692 29404 12756 29408
rect 12692 29348 12696 29404
rect 12696 29348 12752 29404
rect 12752 29348 12756 29404
rect 12692 29344 12756 29348
rect 12772 29404 12836 29408
rect 12772 29348 12776 29404
rect 12776 29348 12832 29404
rect 12832 29348 12836 29404
rect 12772 29344 12836 29348
rect 12852 29404 12916 29408
rect 12852 29348 12856 29404
rect 12856 29348 12912 29404
rect 12912 29348 12916 29404
rect 12852 29344 12916 29348
rect 17612 29404 17676 29408
rect 17612 29348 17616 29404
rect 17616 29348 17672 29404
rect 17672 29348 17676 29404
rect 17612 29344 17676 29348
rect 17692 29404 17756 29408
rect 17692 29348 17696 29404
rect 17696 29348 17752 29404
rect 17752 29348 17756 29404
rect 17692 29344 17756 29348
rect 17772 29404 17836 29408
rect 17772 29348 17776 29404
rect 17776 29348 17832 29404
rect 17832 29348 17836 29404
rect 17772 29344 17836 29348
rect 17852 29404 17916 29408
rect 17852 29348 17856 29404
rect 17856 29348 17912 29404
rect 17912 29348 17916 29404
rect 17852 29344 17916 29348
rect 22612 29404 22676 29408
rect 22612 29348 22616 29404
rect 22616 29348 22672 29404
rect 22672 29348 22676 29404
rect 22612 29344 22676 29348
rect 22692 29404 22756 29408
rect 22692 29348 22696 29404
rect 22696 29348 22752 29404
rect 22752 29348 22756 29404
rect 22692 29344 22756 29348
rect 22772 29404 22836 29408
rect 22772 29348 22776 29404
rect 22776 29348 22832 29404
rect 22832 29348 22836 29404
rect 22772 29344 22836 29348
rect 22852 29404 22916 29408
rect 22852 29348 22856 29404
rect 22856 29348 22912 29404
rect 22912 29348 22916 29404
rect 22852 29344 22916 29348
rect 27612 29404 27676 29408
rect 27612 29348 27616 29404
rect 27616 29348 27672 29404
rect 27672 29348 27676 29404
rect 27612 29344 27676 29348
rect 27692 29404 27756 29408
rect 27692 29348 27696 29404
rect 27696 29348 27752 29404
rect 27752 29348 27756 29404
rect 27692 29344 27756 29348
rect 27772 29404 27836 29408
rect 27772 29348 27776 29404
rect 27776 29348 27832 29404
rect 27832 29348 27836 29404
rect 27772 29344 27836 29348
rect 27852 29404 27916 29408
rect 27852 29348 27856 29404
rect 27856 29348 27912 29404
rect 27912 29348 27916 29404
rect 27852 29344 27916 29348
rect 32612 29404 32676 29408
rect 32612 29348 32616 29404
rect 32616 29348 32672 29404
rect 32672 29348 32676 29404
rect 32612 29344 32676 29348
rect 32692 29404 32756 29408
rect 32692 29348 32696 29404
rect 32696 29348 32752 29404
rect 32752 29348 32756 29404
rect 32692 29344 32756 29348
rect 32772 29404 32836 29408
rect 32772 29348 32776 29404
rect 32776 29348 32832 29404
rect 32832 29348 32836 29404
rect 32772 29344 32836 29348
rect 32852 29404 32916 29408
rect 32852 29348 32856 29404
rect 32856 29348 32912 29404
rect 32912 29348 32916 29404
rect 32852 29344 32916 29348
rect 37612 29404 37676 29408
rect 37612 29348 37616 29404
rect 37616 29348 37672 29404
rect 37672 29348 37676 29404
rect 37612 29344 37676 29348
rect 37692 29404 37756 29408
rect 37692 29348 37696 29404
rect 37696 29348 37752 29404
rect 37752 29348 37756 29404
rect 37692 29344 37756 29348
rect 37772 29404 37836 29408
rect 37772 29348 37776 29404
rect 37776 29348 37832 29404
rect 37832 29348 37836 29404
rect 37772 29344 37836 29348
rect 37852 29404 37916 29408
rect 37852 29348 37856 29404
rect 37856 29348 37912 29404
rect 37912 29348 37916 29404
rect 37852 29344 37916 29348
rect 1952 28860 2016 28864
rect 1952 28804 1956 28860
rect 1956 28804 2012 28860
rect 2012 28804 2016 28860
rect 1952 28800 2016 28804
rect 2032 28860 2096 28864
rect 2032 28804 2036 28860
rect 2036 28804 2092 28860
rect 2092 28804 2096 28860
rect 2032 28800 2096 28804
rect 2112 28860 2176 28864
rect 2112 28804 2116 28860
rect 2116 28804 2172 28860
rect 2172 28804 2176 28860
rect 2112 28800 2176 28804
rect 2192 28860 2256 28864
rect 2192 28804 2196 28860
rect 2196 28804 2252 28860
rect 2252 28804 2256 28860
rect 2192 28800 2256 28804
rect 6952 28860 7016 28864
rect 6952 28804 6956 28860
rect 6956 28804 7012 28860
rect 7012 28804 7016 28860
rect 6952 28800 7016 28804
rect 7032 28860 7096 28864
rect 7032 28804 7036 28860
rect 7036 28804 7092 28860
rect 7092 28804 7096 28860
rect 7032 28800 7096 28804
rect 7112 28860 7176 28864
rect 7112 28804 7116 28860
rect 7116 28804 7172 28860
rect 7172 28804 7176 28860
rect 7112 28800 7176 28804
rect 7192 28860 7256 28864
rect 7192 28804 7196 28860
rect 7196 28804 7252 28860
rect 7252 28804 7256 28860
rect 7192 28800 7256 28804
rect 11952 28860 12016 28864
rect 11952 28804 11956 28860
rect 11956 28804 12012 28860
rect 12012 28804 12016 28860
rect 11952 28800 12016 28804
rect 12032 28860 12096 28864
rect 12032 28804 12036 28860
rect 12036 28804 12092 28860
rect 12092 28804 12096 28860
rect 12032 28800 12096 28804
rect 12112 28860 12176 28864
rect 12112 28804 12116 28860
rect 12116 28804 12172 28860
rect 12172 28804 12176 28860
rect 12112 28800 12176 28804
rect 12192 28860 12256 28864
rect 12192 28804 12196 28860
rect 12196 28804 12252 28860
rect 12252 28804 12256 28860
rect 12192 28800 12256 28804
rect 16952 28860 17016 28864
rect 16952 28804 16956 28860
rect 16956 28804 17012 28860
rect 17012 28804 17016 28860
rect 16952 28800 17016 28804
rect 17032 28860 17096 28864
rect 17032 28804 17036 28860
rect 17036 28804 17092 28860
rect 17092 28804 17096 28860
rect 17032 28800 17096 28804
rect 17112 28860 17176 28864
rect 17112 28804 17116 28860
rect 17116 28804 17172 28860
rect 17172 28804 17176 28860
rect 17112 28800 17176 28804
rect 17192 28860 17256 28864
rect 17192 28804 17196 28860
rect 17196 28804 17252 28860
rect 17252 28804 17256 28860
rect 17192 28800 17256 28804
rect 21952 28860 22016 28864
rect 21952 28804 21956 28860
rect 21956 28804 22012 28860
rect 22012 28804 22016 28860
rect 21952 28800 22016 28804
rect 22032 28860 22096 28864
rect 22032 28804 22036 28860
rect 22036 28804 22092 28860
rect 22092 28804 22096 28860
rect 22032 28800 22096 28804
rect 22112 28860 22176 28864
rect 22112 28804 22116 28860
rect 22116 28804 22172 28860
rect 22172 28804 22176 28860
rect 22112 28800 22176 28804
rect 22192 28860 22256 28864
rect 22192 28804 22196 28860
rect 22196 28804 22252 28860
rect 22252 28804 22256 28860
rect 22192 28800 22256 28804
rect 26952 28860 27016 28864
rect 26952 28804 26956 28860
rect 26956 28804 27012 28860
rect 27012 28804 27016 28860
rect 26952 28800 27016 28804
rect 27032 28860 27096 28864
rect 27032 28804 27036 28860
rect 27036 28804 27092 28860
rect 27092 28804 27096 28860
rect 27032 28800 27096 28804
rect 27112 28860 27176 28864
rect 27112 28804 27116 28860
rect 27116 28804 27172 28860
rect 27172 28804 27176 28860
rect 27112 28800 27176 28804
rect 27192 28860 27256 28864
rect 27192 28804 27196 28860
rect 27196 28804 27252 28860
rect 27252 28804 27256 28860
rect 27192 28800 27256 28804
rect 31952 28860 32016 28864
rect 31952 28804 31956 28860
rect 31956 28804 32012 28860
rect 32012 28804 32016 28860
rect 31952 28800 32016 28804
rect 32032 28860 32096 28864
rect 32032 28804 32036 28860
rect 32036 28804 32092 28860
rect 32092 28804 32096 28860
rect 32032 28800 32096 28804
rect 32112 28860 32176 28864
rect 32112 28804 32116 28860
rect 32116 28804 32172 28860
rect 32172 28804 32176 28860
rect 32112 28800 32176 28804
rect 32192 28860 32256 28864
rect 32192 28804 32196 28860
rect 32196 28804 32252 28860
rect 32252 28804 32256 28860
rect 32192 28800 32256 28804
rect 36952 28860 37016 28864
rect 36952 28804 36956 28860
rect 36956 28804 37012 28860
rect 37012 28804 37016 28860
rect 36952 28800 37016 28804
rect 37032 28860 37096 28864
rect 37032 28804 37036 28860
rect 37036 28804 37092 28860
rect 37092 28804 37096 28860
rect 37032 28800 37096 28804
rect 37112 28860 37176 28864
rect 37112 28804 37116 28860
rect 37116 28804 37172 28860
rect 37172 28804 37176 28860
rect 37112 28800 37176 28804
rect 37192 28860 37256 28864
rect 37192 28804 37196 28860
rect 37196 28804 37252 28860
rect 37252 28804 37256 28860
rect 37192 28800 37256 28804
rect 31708 28732 31772 28796
rect 2612 28316 2676 28320
rect 2612 28260 2616 28316
rect 2616 28260 2672 28316
rect 2672 28260 2676 28316
rect 2612 28256 2676 28260
rect 2692 28316 2756 28320
rect 2692 28260 2696 28316
rect 2696 28260 2752 28316
rect 2752 28260 2756 28316
rect 2692 28256 2756 28260
rect 2772 28316 2836 28320
rect 2772 28260 2776 28316
rect 2776 28260 2832 28316
rect 2832 28260 2836 28316
rect 2772 28256 2836 28260
rect 2852 28316 2916 28320
rect 2852 28260 2856 28316
rect 2856 28260 2912 28316
rect 2912 28260 2916 28316
rect 2852 28256 2916 28260
rect 7612 28316 7676 28320
rect 7612 28260 7616 28316
rect 7616 28260 7672 28316
rect 7672 28260 7676 28316
rect 7612 28256 7676 28260
rect 7692 28316 7756 28320
rect 7692 28260 7696 28316
rect 7696 28260 7752 28316
rect 7752 28260 7756 28316
rect 7692 28256 7756 28260
rect 7772 28316 7836 28320
rect 7772 28260 7776 28316
rect 7776 28260 7832 28316
rect 7832 28260 7836 28316
rect 7772 28256 7836 28260
rect 7852 28316 7916 28320
rect 7852 28260 7856 28316
rect 7856 28260 7912 28316
rect 7912 28260 7916 28316
rect 7852 28256 7916 28260
rect 12612 28316 12676 28320
rect 12612 28260 12616 28316
rect 12616 28260 12672 28316
rect 12672 28260 12676 28316
rect 12612 28256 12676 28260
rect 12692 28316 12756 28320
rect 12692 28260 12696 28316
rect 12696 28260 12752 28316
rect 12752 28260 12756 28316
rect 12692 28256 12756 28260
rect 12772 28316 12836 28320
rect 12772 28260 12776 28316
rect 12776 28260 12832 28316
rect 12832 28260 12836 28316
rect 12772 28256 12836 28260
rect 12852 28316 12916 28320
rect 12852 28260 12856 28316
rect 12856 28260 12912 28316
rect 12912 28260 12916 28316
rect 12852 28256 12916 28260
rect 17612 28316 17676 28320
rect 17612 28260 17616 28316
rect 17616 28260 17672 28316
rect 17672 28260 17676 28316
rect 17612 28256 17676 28260
rect 17692 28316 17756 28320
rect 17692 28260 17696 28316
rect 17696 28260 17752 28316
rect 17752 28260 17756 28316
rect 17692 28256 17756 28260
rect 17772 28316 17836 28320
rect 17772 28260 17776 28316
rect 17776 28260 17832 28316
rect 17832 28260 17836 28316
rect 17772 28256 17836 28260
rect 17852 28316 17916 28320
rect 17852 28260 17856 28316
rect 17856 28260 17912 28316
rect 17912 28260 17916 28316
rect 17852 28256 17916 28260
rect 22612 28316 22676 28320
rect 22612 28260 22616 28316
rect 22616 28260 22672 28316
rect 22672 28260 22676 28316
rect 22612 28256 22676 28260
rect 22692 28316 22756 28320
rect 22692 28260 22696 28316
rect 22696 28260 22752 28316
rect 22752 28260 22756 28316
rect 22692 28256 22756 28260
rect 22772 28316 22836 28320
rect 22772 28260 22776 28316
rect 22776 28260 22832 28316
rect 22832 28260 22836 28316
rect 22772 28256 22836 28260
rect 22852 28316 22916 28320
rect 22852 28260 22856 28316
rect 22856 28260 22912 28316
rect 22912 28260 22916 28316
rect 22852 28256 22916 28260
rect 27612 28316 27676 28320
rect 27612 28260 27616 28316
rect 27616 28260 27672 28316
rect 27672 28260 27676 28316
rect 27612 28256 27676 28260
rect 27692 28316 27756 28320
rect 27692 28260 27696 28316
rect 27696 28260 27752 28316
rect 27752 28260 27756 28316
rect 27692 28256 27756 28260
rect 27772 28316 27836 28320
rect 27772 28260 27776 28316
rect 27776 28260 27832 28316
rect 27832 28260 27836 28316
rect 27772 28256 27836 28260
rect 27852 28316 27916 28320
rect 27852 28260 27856 28316
rect 27856 28260 27912 28316
rect 27912 28260 27916 28316
rect 27852 28256 27916 28260
rect 32612 28316 32676 28320
rect 32612 28260 32616 28316
rect 32616 28260 32672 28316
rect 32672 28260 32676 28316
rect 32612 28256 32676 28260
rect 32692 28316 32756 28320
rect 32692 28260 32696 28316
rect 32696 28260 32752 28316
rect 32752 28260 32756 28316
rect 32692 28256 32756 28260
rect 32772 28316 32836 28320
rect 32772 28260 32776 28316
rect 32776 28260 32832 28316
rect 32832 28260 32836 28316
rect 32772 28256 32836 28260
rect 32852 28316 32916 28320
rect 32852 28260 32856 28316
rect 32856 28260 32912 28316
rect 32912 28260 32916 28316
rect 32852 28256 32916 28260
rect 37612 28316 37676 28320
rect 37612 28260 37616 28316
rect 37616 28260 37672 28316
rect 37672 28260 37676 28316
rect 37612 28256 37676 28260
rect 37692 28316 37756 28320
rect 37692 28260 37696 28316
rect 37696 28260 37752 28316
rect 37752 28260 37756 28316
rect 37692 28256 37756 28260
rect 37772 28316 37836 28320
rect 37772 28260 37776 28316
rect 37776 28260 37832 28316
rect 37832 28260 37836 28316
rect 37772 28256 37836 28260
rect 37852 28316 37916 28320
rect 37852 28260 37856 28316
rect 37856 28260 37912 28316
rect 37912 28260 37916 28316
rect 37852 28256 37916 28260
rect 1952 27772 2016 27776
rect 1952 27716 1956 27772
rect 1956 27716 2012 27772
rect 2012 27716 2016 27772
rect 1952 27712 2016 27716
rect 2032 27772 2096 27776
rect 2032 27716 2036 27772
rect 2036 27716 2092 27772
rect 2092 27716 2096 27772
rect 2032 27712 2096 27716
rect 2112 27772 2176 27776
rect 2112 27716 2116 27772
rect 2116 27716 2172 27772
rect 2172 27716 2176 27772
rect 2112 27712 2176 27716
rect 2192 27772 2256 27776
rect 2192 27716 2196 27772
rect 2196 27716 2252 27772
rect 2252 27716 2256 27772
rect 2192 27712 2256 27716
rect 6952 27772 7016 27776
rect 6952 27716 6956 27772
rect 6956 27716 7012 27772
rect 7012 27716 7016 27772
rect 6952 27712 7016 27716
rect 7032 27772 7096 27776
rect 7032 27716 7036 27772
rect 7036 27716 7092 27772
rect 7092 27716 7096 27772
rect 7032 27712 7096 27716
rect 7112 27772 7176 27776
rect 7112 27716 7116 27772
rect 7116 27716 7172 27772
rect 7172 27716 7176 27772
rect 7112 27712 7176 27716
rect 7192 27772 7256 27776
rect 7192 27716 7196 27772
rect 7196 27716 7252 27772
rect 7252 27716 7256 27772
rect 7192 27712 7256 27716
rect 11952 27772 12016 27776
rect 11952 27716 11956 27772
rect 11956 27716 12012 27772
rect 12012 27716 12016 27772
rect 11952 27712 12016 27716
rect 12032 27772 12096 27776
rect 12032 27716 12036 27772
rect 12036 27716 12092 27772
rect 12092 27716 12096 27772
rect 12032 27712 12096 27716
rect 12112 27772 12176 27776
rect 12112 27716 12116 27772
rect 12116 27716 12172 27772
rect 12172 27716 12176 27772
rect 12112 27712 12176 27716
rect 12192 27772 12256 27776
rect 12192 27716 12196 27772
rect 12196 27716 12252 27772
rect 12252 27716 12256 27772
rect 12192 27712 12256 27716
rect 16952 27772 17016 27776
rect 16952 27716 16956 27772
rect 16956 27716 17012 27772
rect 17012 27716 17016 27772
rect 16952 27712 17016 27716
rect 17032 27772 17096 27776
rect 17032 27716 17036 27772
rect 17036 27716 17092 27772
rect 17092 27716 17096 27772
rect 17032 27712 17096 27716
rect 17112 27772 17176 27776
rect 17112 27716 17116 27772
rect 17116 27716 17172 27772
rect 17172 27716 17176 27772
rect 17112 27712 17176 27716
rect 17192 27772 17256 27776
rect 17192 27716 17196 27772
rect 17196 27716 17252 27772
rect 17252 27716 17256 27772
rect 17192 27712 17256 27716
rect 21952 27772 22016 27776
rect 21952 27716 21956 27772
rect 21956 27716 22012 27772
rect 22012 27716 22016 27772
rect 21952 27712 22016 27716
rect 22032 27772 22096 27776
rect 22032 27716 22036 27772
rect 22036 27716 22092 27772
rect 22092 27716 22096 27772
rect 22032 27712 22096 27716
rect 22112 27772 22176 27776
rect 22112 27716 22116 27772
rect 22116 27716 22172 27772
rect 22172 27716 22176 27772
rect 22112 27712 22176 27716
rect 22192 27772 22256 27776
rect 22192 27716 22196 27772
rect 22196 27716 22252 27772
rect 22252 27716 22256 27772
rect 22192 27712 22256 27716
rect 26952 27772 27016 27776
rect 26952 27716 26956 27772
rect 26956 27716 27012 27772
rect 27012 27716 27016 27772
rect 26952 27712 27016 27716
rect 27032 27772 27096 27776
rect 27032 27716 27036 27772
rect 27036 27716 27092 27772
rect 27092 27716 27096 27772
rect 27032 27712 27096 27716
rect 27112 27772 27176 27776
rect 27112 27716 27116 27772
rect 27116 27716 27172 27772
rect 27172 27716 27176 27772
rect 27112 27712 27176 27716
rect 27192 27772 27256 27776
rect 27192 27716 27196 27772
rect 27196 27716 27252 27772
rect 27252 27716 27256 27772
rect 27192 27712 27256 27716
rect 31952 27772 32016 27776
rect 31952 27716 31956 27772
rect 31956 27716 32012 27772
rect 32012 27716 32016 27772
rect 31952 27712 32016 27716
rect 32032 27772 32096 27776
rect 32032 27716 32036 27772
rect 32036 27716 32092 27772
rect 32092 27716 32096 27772
rect 32032 27712 32096 27716
rect 32112 27772 32176 27776
rect 32112 27716 32116 27772
rect 32116 27716 32172 27772
rect 32172 27716 32176 27772
rect 32112 27712 32176 27716
rect 32192 27772 32256 27776
rect 32192 27716 32196 27772
rect 32196 27716 32252 27772
rect 32252 27716 32256 27772
rect 32192 27712 32256 27716
rect 36952 27772 37016 27776
rect 36952 27716 36956 27772
rect 36956 27716 37012 27772
rect 37012 27716 37016 27772
rect 36952 27712 37016 27716
rect 37032 27772 37096 27776
rect 37032 27716 37036 27772
rect 37036 27716 37092 27772
rect 37092 27716 37096 27772
rect 37032 27712 37096 27716
rect 37112 27772 37176 27776
rect 37112 27716 37116 27772
rect 37116 27716 37172 27772
rect 37172 27716 37176 27772
rect 37112 27712 37176 27716
rect 37192 27772 37256 27776
rect 37192 27716 37196 27772
rect 37196 27716 37252 27772
rect 37252 27716 37256 27772
rect 37192 27712 37256 27716
rect 2612 27228 2676 27232
rect 2612 27172 2616 27228
rect 2616 27172 2672 27228
rect 2672 27172 2676 27228
rect 2612 27168 2676 27172
rect 2692 27228 2756 27232
rect 2692 27172 2696 27228
rect 2696 27172 2752 27228
rect 2752 27172 2756 27228
rect 2692 27168 2756 27172
rect 2772 27228 2836 27232
rect 2772 27172 2776 27228
rect 2776 27172 2832 27228
rect 2832 27172 2836 27228
rect 2772 27168 2836 27172
rect 2852 27228 2916 27232
rect 2852 27172 2856 27228
rect 2856 27172 2912 27228
rect 2912 27172 2916 27228
rect 2852 27168 2916 27172
rect 7612 27228 7676 27232
rect 7612 27172 7616 27228
rect 7616 27172 7672 27228
rect 7672 27172 7676 27228
rect 7612 27168 7676 27172
rect 7692 27228 7756 27232
rect 7692 27172 7696 27228
rect 7696 27172 7752 27228
rect 7752 27172 7756 27228
rect 7692 27168 7756 27172
rect 7772 27228 7836 27232
rect 7772 27172 7776 27228
rect 7776 27172 7832 27228
rect 7832 27172 7836 27228
rect 7772 27168 7836 27172
rect 7852 27228 7916 27232
rect 7852 27172 7856 27228
rect 7856 27172 7912 27228
rect 7912 27172 7916 27228
rect 7852 27168 7916 27172
rect 12612 27228 12676 27232
rect 12612 27172 12616 27228
rect 12616 27172 12672 27228
rect 12672 27172 12676 27228
rect 12612 27168 12676 27172
rect 12692 27228 12756 27232
rect 12692 27172 12696 27228
rect 12696 27172 12752 27228
rect 12752 27172 12756 27228
rect 12692 27168 12756 27172
rect 12772 27228 12836 27232
rect 12772 27172 12776 27228
rect 12776 27172 12832 27228
rect 12832 27172 12836 27228
rect 12772 27168 12836 27172
rect 12852 27228 12916 27232
rect 12852 27172 12856 27228
rect 12856 27172 12912 27228
rect 12912 27172 12916 27228
rect 12852 27168 12916 27172
rect 17612 27228 17676 27232
rect 17612 27172 17616 27228
rect 17616 27172 17672 27228
rect 17672 27172 17676 27228
rect 17612 27168 17676 27172
rect 17692 27228 17756 27232
rect 17692 27172 17696 27228
rect 17696 27172 17752 27228
rect 17752 27172 17756 27228
rect 17692 27168 17756 27172
rect 17772 27228 17836 27232
rect 17772 27172 17776 27228
rect 17776 27172 17832 27228
rect 17832 27172 17836 27228
rect 17772 27168 17836 27172
rect 17852 27228 17916 27232
rect 17852 27172 17856 27228
rect 17856 27172 17912 27228
rect 17912 27172 17916 27228
rect 17852 27168 17916 27172
rect 22612 27228 22676 27232
rect 22612 27172 22616 27228
rect 22616 27172 22672 27228
rect 22672 27172 22676 27228
rect 22612 27168 22676 27172
rect 22692 27228 22756 27232
rect 22692 27172 22696 27228
rect 22696 27172 22752 27228
rect 22752 27172 22756 27228
rect 22692 27168 22756 27172
rect 22772 27228 22836 27232
rect 22772 27172 22776 27228
rect 22776 27172 22832 27228
rect 22832 27172 22836 27228
rect 22772 27168 22836 27172
rect 22852 27228 22916 27232
rect 22852 27172 22856 27228
rect 22856 27172 22912 27228
rect 22912 27172 22916 27228
rect 22852 27168 22916 27172
rect 27612 27228 27676 27232
rect 27612 27172 27616 27228
rect 27616 27172 27672 27228
rect 27672 27172 27676 27228
rect 27612 27168 27676 27172
rect 27692 27228 27756 27232
rect 27692 27172 27696 27228
rect 27696 27172 27752 27228
rect 27752 27172 27756 27228
rect 27692 27168 27756 27172
rect 27772 27228 27836 27232
rect 27772 27172 27776 27228
rect 27776 27172 27832 27228
rect 27832 27172 27836 27228
rect 27772 27168 27836 27172
rect 27852 27228 27916 27232
rect 27852 27172 27856 27228
rect 27856 27172 27912 27228
rect 27912 27172 27916 27228
rect 27852 27168 27916 27172
rect 32612 27228 32676 27232
rect 32612 27172 32616 27228
rect 32616 27172 32672 27228
rect 32672 27172 32676 27228
rect 32612 27168 32676 27172
rect 32692 27228 32756 27232
rect 32692 27172 32696 27228
rect 32696 27172 32752 27228
rect 32752 27172 32756 27228
rect 32692 27168 32756 27172
rect 32772 27228 32836 27232
rect 32772 27172 32776 27228
rect 32776 27172 32832 27228
rect 32832 27172 32836 27228
rect 32772 27168 32836 27172
rect 32852 27228 32916 27232
rect 32852 27172 32856 27228
rect 32856 27172 32912 27228
rect 32912 27172 32916 27228
rect 32852 27168 32916 27172
rect 37612 27228 37676 27232
rect 37612 27172 37616 27228
rect 37616 27172 37672 27228
rect 37672 27172 37676 27228
rect 37612 27168 37676 27172
rect 37692 27228 37756 27232
rect 37692 27172 37696 27228
rect 37696 27172 37752 27228
rect 37752 27172 37756 27228
rect 37692 27168 37756 27172
rect 37772 27228 37836 27232
rect 37772 27172 37776 27228
rect 37776 27172 37832 27228
rect 37832 27172 37836 27228
rect 37772 27168 37836 27172
rect 37852 27228 37916 27232
rect 37852 27172 37856 27228
rect 37856 27172 37912 27228
rect 37912 27172 37916 27228
rect 37852 27168 37916 27172
rect 1952 26684 2016 26688
rect 1952 26628 1956 26684
rect 1956 26628 2012 26684
rect 2012 26628 2016 26684
rect 1952 26624 2016 26628
rect 2032 26684 2096 26688
rect 2032 26628 2036 26684
rect 2036 26628 2092 26684
rect 2092 26628 2096 26684
rect 2032 26624 2096 26628
rect 2112 26684 2176 26688
rect 2112 26628 2116 26684
rect 2116 26628 2172 26684
rect 2172 26628 2176 26684
rect 2112 26624 2176 26628
rect 2192 26684 2256 26688
rect 2192 26628 2196 26684
rect 2196 26628 2252 26684
rect 2252 26628 2256 26684
rect 2192 26624 2256 26628
rect 6952 26684 7016 26688
rect 6952 26628 6956 26684
rect 6956 26628 7012 26684
rect 7012 26628 7016 26684
rect 6952 26624 7016 26628
rect 7032 26684 7096 26688
rect 7032 26628 7036 26684
rect 7036 26628 7092 26684
rect 7092 26628 7096 26684
rect 7032 26624 7096 26628
rect 7112 26684 7176 26688
rect 7112 26628 7116 26684
rect 7116 26628 7172 26684
rect 7172 26628 7176 26684
rect 7112 26624 7176 26628
rect 7192 26684 7256 26688
rect 7192 26628 7196 26684
rect 7196 26628 7252 26684
rect 7252 26628 7256 26684
rect 7192 26624 7256 26628
rect 11952 26684 12016 26688
rect 11952 26628 11956 26684
rect 11956 26628 12012 26684
rect 12012 26628 12016 26684
rect 11952 26624 12016 26628
rect 12032 26684 12096 26688
rect 12032 26628 12036 26684
rect 12036 26628 12092 26684
rect 12092 26628 12096 26684
rect 12032 26624 12096 26628
rect 12112 26684 12176 26688
rect 12112 26628 12116 26684
rect 12116 26628 12172 26684
rect 12172 26628 12176 26684
rect 12112 26624 12176 26628
rect 12192 26684 12256 26688
rect 12192 26628 12196 26684
rect 12196 26628 12252 26684
rect 12252 26628 12256 26684
rect 12192 26624 12256 26628
rect 16952 26684 17016 26688
rect 16952 26628 16956 26684
rect 16956 26628 17012 26684
rect 17012 26628 17016 26684
rect 16952 26624 17016 26628
rect 17032 26684 17096 26688
rect 17032 26628 17036 26684
rect 17036 26628 17092 26684
rect 17092 26628 17096 26684
rect 17032 26624 17096 26628
rect 17112 26684 17176 26688
rect 17112 26628 17116 26684
rect 17116 26628 17172 26684
rect 17172 26628 17176 26684
rect 17112 26624 17176 26628
rect 17192 26684 17256 26688
rect 17192 26628 17196 26684
rect 17196 26628 17252 26684
rect 17252 26628 17256 26684
rect 17192 26624 17256 26628
rect 21952 26684 22016 26688
rect 21952 26628 21956 26684
rect 21956 26628 22012 26684
rect 22012 26628 22016 26684
rect 21952 26624 22016 26628
rect 22032 26684 22096 26688
rect 22032 26628 22036 26684
rect 22036 26628 22092 26684
rect 22092 26628 22096 26684
rect 22032 26624 22096 26628
rect 22112 26684 22176 26688
rect 22112 26628 22116 26684
rect 22116 26628 22172 26684
rect 22172 26628 22176 26684
rect 22112 26624 22176 26628
rect 22192 26684 22256 26688
rect 22192 26628 22196 26684
rect 22196 26628 22252 26684
rect 22252 26628 22256 26684
rect 22192 26624 22256 26628
rect 26952 26684 27016 26688
rect 26952 26628 26956 26684
rect 26956 26628 27012 26684
rect 27012 26628 27016 26684
rect 26952 26624 27016 26628
rect 27032 26684 27096 26688
rect 27032 26628 27036 26684
rect 27036 26628 27092 26684
rect 27092 26628 27096 26684
rect 27032 26624 27096 26628
rect 27112 26684 27176 26688
rect 27112 26628 27116 26684
rect 27116 26628 27172 26684
rect 27172 26628 27176 26684
rect 27112 26624 27176 26628
rect 27192 26684 27256 26688
rect 27192 26628 27196 26684
rect 27196 26628 27252 26684
rect 27252 26628 27256 26684
rect 27192 26624 27256 26628
rect 31952 26684 32016 26688
rect 31952 26628 31956 26684
rect 31956 26628 32012 26684
rect 32012 26628 32016 26684
rect 31952 26624 32016 26628
rect 32032 26684 32096 26688
rect 32032 26628 32036 26684
rect 32036 26628 32092 26684
rect 32092 26628 32096 26684
rect 32032 26624 32096 26628
rect 32112 26684 32176 26688
rect 32112 26628 32116 26684
rect 32116 26628 32172 26684
rect 32172 26628 32176 26684
rect 32112 26624 32176 26628
rect 32192 26684 32256 26688
rect 32192 26628 32196 26684
rect 32196 26628 32252 26684
rect 32252 26628 32256 26684
rect 32192 26624 32256 26628
rect 36952 26684 37016 26688
rect 36952 26628 36956 26684
rect 36956 26628 37012 26684
rect 37012 26628 37016 26684
rect 36952 26624 37016 26628
rect 37032 26684 37096 26688
rect 37032 26628 37036 26684
rect 37036 26628 37092 26684
rect 37092 26628 37096 26684
rect 37032 26624 37096 26628
rect 37112 26684 37176 26688
rect 37112 26628 37116 26684
rect 37116 26628 37172 26684
rect 37172 26628 37176 26684
rect 37112 26624 37176 26628
rect 37192 26684 37256 26688
rect 37192 26628 37196 26684
rect 37196 26628 37252 26684
rect 37252 26628 37256 26684
rect 37192 26624 37256 26628
rect 2612 26140 2676 26144
rect 2612 26084 2616 26140
rect 2616 26084 2672 26140
rect 2672 26084 2676 26140
rect 2612 26080 2676 26084
rect 2692 26140 2756 26144
rect 2692 26084 2696 26140
rect 2696 26084 2752 26140
rect 2752 26084 2756 26140
rect 2692 26080 2756 26084
rect 2772 26140 2836 26144
rect 2772 26084 2776 26140
rect 2776 26084 2832 26140
rect 2832 26084 2836 26140
rect 2772 26080 2836 26084
rect 2852 26140 2916 26144
rect 2852 26084 2856 26140
rect 2856 26084 2912 26140
rect 2912 26084 2916 26140
rect 2852 26080 2916 26084
rect 7612 26140 7676 26144
rect 7612 26084 7616 26140
rect 7616 26084 7672 26140
rect 7672 26084 7676 26140
rect 7612 26080 7676 26084
rect 7692 26140 7756 26144
rect 7692 26084 7696 26140
rect 7696 26084 7752 26140
rect 7752 26084 7756 26140
rect 7692 26080 7756 26084
rect 7772 26140 7836 26144
rect 7772 26084 7776 26140
rect 7776 26084 7832 26140
rect 7832 26084 7836 26140
rect 7772 26080 7836 26084
rect 7852 26140 7916 26144
rect 7852 26084 7856 26140
rect 7856 26084 7912 26140
rect 7912 26084 7916 26140
rect 7852 26080 7916 26084
rect 12612 26140 12676 26144
rect 12612 26084 12616 26140
rect 12616 26084 12672 26140
rect 12672 26084 12676 26140
rect 12612 26080 12676 26084
rect 12692 26140 12756 26144
rect 12692 26084 12696 26140
rect 12696 26084 12752 26140
rect 12752 26084 12756 26140
rect 12692 26080 12756 26084
rect 12772 26140 12836 26144
rect 12772 26084 12776 26140
rect 12776 26084 12832 26140
rect 12832 26084 12836 26140
rect 12772 26080 12836 26084
rect 12852 26140 12916 26144
rect 12852 26084 12856 26140
rect 12856 26084 12912 26140
rect 12912 26084 12916 26140
rect 12852 26080 12916 26084
rect 17612 26140 17676 26144
rect 17612 26084 17616 26140
rect 17616 26084 17672 26140
rect 17672 26084 17676 26140
rect 17612 26080 17676 26084
rect 17692 26140 17756 26144
rect 17692 26084 17696 26140
rect 17696 26084 17752 26140
rect 17752 26084 17756 26140
rect 17692 26080 17756 26084
rect 17772 26140 17836 26144
rect 17772 26084 17776 26140
rect 17776 26084 17832 26140
rect 17832 26084 17836 26140
rect 17772 26080 17836 26084
rect 17852 26140 17916 26144
rect 17852 26084 17856 26140
rect 17856 26084 17912 26140
rect 17912 26084 17916 26140
rect 17852 26080 17916 26084
rect 22612 26140 22676 26144
rect 22612 26084 22616 26140
rect 22616 26084 22672 26140
rect 22672 26084 22676 26140
rect 22612 26080 22676 26084
rect 22692 26140 22756 26144
rect 22692 26084 22696 26140
rect 22696 26084 22752 26140
rect 22752 26084 22756 26140
rect 22692 26080 22756 26084
rect 22772 26140 22836 26144
rect 22772 26084 22776 26140
rect 22776 26084 22832 26140
rect 22832 26084 22836 26140
rect 22772 26080 22836 26084
rect 22852 26140 22916 26144
rect 22852 26084 22856 26140
rect 22856 26084 22912 26140
rect 22912 26084 22916 26140
rect 22852 26080 22916 26084
rect 27612 26140 27676 26144
rect 27612 26084 27616 26140
rect 27616 26084 27672 26140
rect 27672 26084 27676 26140
rect 27612 26080 27676 26084
rect 27692 26140 27756 26144
rect 27692 26084 27696 26140
rect 27696 26084 27752 26140
rect 27752 26084 27756 26140
rect 27692 26080 27756 26084
rect 27772 26140 27836 26144
rect 27772 26084 27776 26140
rect 27776 26084 27832 26140
rect 27832 26084 27836 26140
rect 27772 26080 27836 26084
rect 27852 26140 27916 26144
rect 27852 26084 27856 26140
rect 27856 26084 27912 26140
rect 27912 26084 27916 26140
rect 27852 26080 27916 26084
rect 32612 26140 32676 26144
rect 32612 26084 32616 26140
rect 32616 26084 32672 26140
rect 32672 26084 32676 26140
rect 32612 26080 32676 26084
rect 32692 26140 32756 26144
rect 32692 26084 32696 26140
rect 32696 26084 32752 26140
rect 32752 26084 32756 26140
rect 32692 26080 32756 26084
rect 32772 26140 32836 26144
rect 32772 26084 32776 26140
rect 32776 26084 32832 26140
rect 32832 26084 32836 26140
rect 32772 26080 32836 26084
rect 32852 26140 32916 26144
rect 32852 26084 32856 26140
rect 32856 26084 32912 26140
rect 32912 26084 32916 26140
rect 32852 26080 32916 26084
rect 37612 26140 37676 26144
rect 37612 26084 37616 26140
rect 37616 26084 37672 26140
rect 37672 26084 37676 26140
rect 37612 26080 37676 26084
rect 37692 26140 37756 26144
rect 37692 26084 37696 26140
rect 37696 26084 37752 26140
rect 37752 26084 37756 26140
rect 37692 26080 37756 26084
rect 37772 26140 37836 26144
rect 37772 26084 37776 26140
rect 37776 26084 37832 26140
rect 37832 26084 37836 26140
rect 37772 26080 37836 26084
rect 37852 26140 37916 26144
rect 37852 26084 37856 26140
rect 37856 26084 37912 26140
rect 37912 26084 37916 26140
rect 37852 26080 37916 26084
rect 1952 25596 2016 25600
rect 1952 25540 1956 25596
rect 1956 25540 2012 25596
rect 2012 25540 2016 25596
rect 1952 25536 2016 25540
rect 2032 25596 2096 25600
rect 2032 25540 2036 25596
rect 2036 25540 2092 25596
rect 2092 25540 2096 25596
rect 2032 25536 2096 25540
rect 2112 25596 2176 25600
rect 2112 25540 2116 25596
rect 2116 25540 2172 25596
rect 2172 25540 2176 25596
rect 2112 25536 2176 25540
rect 2192 25596 2256 25600
rect 2192 25540 2196 25596
rect 2196 25540 2252 25596
rect 2252 25540 2256 25596
rect 2192 25536 2256 25540
rect 6952 25596 7016 25600
rect 6952 25540 6956 25596
rect 6956 25540 7012 25596
rect 7012 25540 7016 25596
rect 6952 25536 7016 25540
rect 7032 25596 7096 25600
rect 7032 25540 7036 25596
rect 7036 25540 7092 25596
rect 7092 25540 7096 25596
rect 7032 25536 7096 25540
rect 7112 25596 7176 25600
rect 7112 25540 7116 25596
rect 7116 25540 7172 25596
rect 7172 25540 7176 25596
rect 7112 25536 7176 25540
rect 7192 25596 7256 25600
rect 7192 25540 7196 25596
rect 7196 25540 7252 25596
rect 7252 25540 7256 25596
rect 7192 25536 7256 25540
rect 11952 25596 12016 25600
rect 11952 25540 11956 25596
rect 11956 25540 12012 25596
rect 12012 25540 12016 25596
rect 11952 25536 12016 25540
rect 12032 25596 12096 25600
rect 12032 25540 12036 25596
rect 12036 25540 12092 25596
rect 12092 25540 12096 25596
rect 12032 25536 12096 25540
rect 12112 25596 12176 25600
rect 12112 25540 12116 25596
rect 12116 25540 12172 25596
rect 12172 25540 12176 25596
rect 12112 25536 12176 25540
rect 12192 25596 12256 25600
rect 12192 25540 12196 25596
rect 12196 25540 12252 25596
rect 12252 25540 12256 25596
rect 12192 25536 12256 25540
rect 16952 25596 17016 25600
rect 16952 25540 16956 25596
rect 16956 25540 17012 25596
rect 17012 25540 17016 25596
rect 16952 25536 17016 25540
rect 17032 25596 17096 25600
rect 17032 25540 17036 25596
rect 17036 25540 17092 25596
rect 17092 25540 17096 25596
rect 17032 25536 17096 25540
rect 17112 25596 17176 25600
rect 17112 25540 17116 25596
rect 17116 25540 17172 25596
rect 17172 25540 17176 25596
rect 17112 25536 17176 25540
rect 17192 25596 17256 25600
rect 17192 25540 17196 25596
rect 17196 25540 17252 25596
rect 17252 25540 17256 25596
rect 17192 25536 17256 25540
rect 21952 25596 22016 25600
rect 21952 25540 21956 25596
rect 21956 25540 22012 25596
rect 22012 25540 22016 25596
rect 21952 25536 22016 25540
rect 22032 25596 22096 25600
rect 22032 25540 22036 25596
rect 22036 25540 22092 25596
rect 22092 25540 22096 25596
rect 22032 25536 22096 25540
rect 22112 25596 22176 25600
rect 22112 25540 22116 25596
rect 22116 25540 22172 25596
rect 22172 25540 22176 25596
rect 22112 25536 22176 25540
rect 22192 25596 22256 25600
rect 22192 25540 22196 25596
rect 22196 25540 22252 25596
rect 22252 25540 22256 25596
rect 22192 25536 22256 25540
rect 26952 25596 27016 25600
rect 26952 25540 26956 25596
rect 26956 25540 27012 25596
rect 27012 25540 27016 25596
rect 26952 25536 27016 25540
rect 27032 25596 27096 25600
rect 27032 25540 27036 25596
rect 27036 25540 27092 25596
rect 27092 25540 27096 25596
rect 27032 25536 27096 25540
rect 27112 25596 27176 25600
rect 27112 25540 27116 25596
rect 27116 25540 27172 25596
rect 27172 25540 27176 25596
rect 27112 25536 27176 25540
rect 27192 25596 27256 25600
rect 27192 25540 27196 25596
rect 27196 25540 27252 25596
rect 27252 25540 27256 25596
rect 27192 25536 27256 25540
rect 31952 25596 32016 25600
rect 31952 25540 31956 25596
rect 31956 25540 32012 25596
rect 32012 25540 32016 25596
rect 31952 25536 32016 25540
rect 32032 25596 32096 25600
rect 32032 25540 32036 25596
rect 32036 25540 32092 25596
rect 32092 25540 32096 25596
rect 32032 25536 32096 25540
rect 32112 25596 32176 25600
rect 32112 25540 32116 25596
rect 32116 25540 32172 25596
rect 32172 25540 32176 25596
rect 32112 25536 32176 25540
rect 32192 25596 32256 25600
rect 32192 25540 32196 25596
rect 32196 25540 32252 25596
rect 32252 25540 32256 25596
rect 32192 25536 32256 25540
rect 36952 25596 37016 25600
rect 36952 25540 36956 25596
rect 36956 25540 37012 25596
rect 37012 25540 37016 25596
rect 36952 25536 37016 25540
rect 37032 25596 37096 25600
rect 37032 25540 37036 25596
rect 37036 25540 37092 25596
rect 37092 25540 37096 25596
rect 37032 25536 37096 25540
rect 37112 25596 37176 25600
rect 37112 25540 37116 25596
rect 37116 25540 37172 25596
rect 37172 25540 37176 25596
rect 37112 25536 37176 25540
rect 37192 25596 37256 25600
rect 37192 25540 37196 25596
rect 37196 25540 37252 25596
rect 37252 25540 37256 25596
rect 37192 25536 37256 25540
rect 2612 25052 2676 25056
rect 2612 24996 2616 25052
rect 2616 24996 2672 25052
rect 2672 24996 2676 25052
rect 2612 24992 2676 24996
rect 2692 25052 2756 25056
rect 2692 24996 2696 25052
rect 2696 24996 2752 25052
rect 2752 24996 2756 25052
rect 2692 24992 2756 24996
rect 2772 25052 2836 25056
rect 2772 24996 2776 25052
rect 2776 24996 2832 25052
rect 2832 24996 2836 25052
rect 2772 24992 2836 24996
rect 2852 25052 2916 25056
rect 2852 24996 2856 25052
rect 2856 24996 2912 25052
rect 2912 24996 2916 25052
rect 2852 24992 2916 24996
rect 7612 25052 7676 25056
rect 7612 24996 7616 25052
rect 7616 24996 7672 25052
rect 7672 24996 7676 25052
rect 7612 24992 7676 24996
rect 7692 25052 7756 25056
rect 7692 24996 7696 25052
rect 7696 24996 7752 25052
rect 7752 24996 7756 25052
rect 7692 24992 7756 24996
rect 7772 25052 7836 25056
rect 7772 24996 7776 25052
rect 7776 24996 7832 25052
rect 7832 24996 7836 25052
rect 7772 24992 7836 24996
rect 7852 25052 7916 25056
rect 7852 24996 7856 25052
rect 7856 24996 7912 25052
rect 7912 24996 7916 25052
rect 7852 24992 7916 24996
rect 12612 25052 12676 25056
rect 12612 24996 12616 25052
rect 12616 24996 12672 25052
rect 12672 24996 12676 25052
rect 12612 24992 12676 24996
rect 12692 25052 12756 25056
rect 12692 24996 12696 25052
rect 12696 24996 12752 25052
rect 12752 24996 12756 25052
rect 12692 24992 12756 24996
rect 12772 25052 12836 25056
rect 12772 24996 12776 25052
rect 12776 24996 12832 25052
rect 12832 24996 12836 25052
rect 12772 24992 12836 24996
rect 12852 25052 12916 25056
rect 12852 24996 12856 25052
rect 12856 24996 12912 25052
rect 12912 24996 12916 25052
rect 12852 24992 12916 24996
rect 17612 25052 17676 25056
rect 17612 24996 17616 25052
rect 17616 24996 17672 25052
rect 17672 24996 17676 25052
rect 17612 24992 17676 24996
rect 17692 25052 17756 25056
rect 17692 24996 17696 25052
rect 17696 24996 17752 25052
rect 17752 24996 17756 25052
rect 17692 24992 17756 24996
rect 17772 25052 17836 25056
rect 17772 24996 17776 25052
rect 17776 24996 17832 25052
rect 17832 24996 17836 25052
rect 17772 24992 17836 24996
rect 17852 25052 17916 25056
rect 17852 24996 17856 25052
rect 17856 24996 17912 25052
rect 17912 24996 17916 25052
rect 17852 24992 17916 24996
rect 22612 25052 22676 25056
rect 22612 24996 22616 25052
rect 22616 24996 22672 25052
rect 22672 24996 22676 25052
rect 22612 24992 22676 24996
rect 22692 25052 22756 25056
rect 22692 24996 22696 25052
rect 22696 24996 22752 25052
rect 22752 24996 22756 25052
rect 22692 24992 22756 24996
rect 22772 25052 22836 25056
rect 22772 24996 22776 25052
rect 22776 24996 22832 25052
rect 22832 24996 22836 25052
rect 22772 24992 22836 24996
rect 22852 25052 22916 25056
rect 22852 24996 22856 25052
rect 22856 24996 22912 25052
rect 22912 24996 22916 25052
rect 22852 24992 22916 24996
rect 27612 25052 27676 25056
rect 27612 24996 27616 25052
rect 27616 24996 27672 25052
rect 27672 24996 27676 25052
rect 27612 24992 27676 24996
rect 27692 25052 27756 25056
rect 27692 24996 27696 25052
rect 27696 24996 27752 25052
rect 27752 24996 27756 25052
rect 27692 24992 27756 24996
rect 27772 25052 27836 25056
rect 27772 24996 27776 25052
rect 27776 24996 27832 25052
rect 27832 24996 27836 25052
rect 27772 24992 27836 24996
rect 27852 25052 27916 25056
rect 27852 24996 27856 25052
rect 27856 24996 27912 25052
rect 27912 24996 27916 25052
rect 27852 24992 27916 24996
rect 32612 25052 32676 25056
rect 32612 24996 32616 25052
rect 32616 24996 32672 25052
rect 32672 24996 32676 25052
rect 32612 24992 32676 24996
rect 32692 25052 32756 25056
rect 32692 24996 32696 25052
rect 32696 24996 32752 25052
rect 32752 24996 32756 25052
rect 32692 24992 32756 24996
rect 32772 25052 32836 25056
rect 32772 24996 32776 25052
rect 32776 24996 32832 25052
rect 32832 24996 32836 25052
rect 32772 24992 32836 24996
rect 32852 25052 32916 25056
rect 32852 24996 32856 25052
rect 32856 24996 32912 25052
rect 32912 24996 32916 25052
rect 32852 24992 32916 24996
rect 37612 25052 37676 25056
rect 37612 24996 37616 25052
rect 37616 24996 37672 25052
rect 37672 24996 37676 25052
rect 37612 24992 37676 24996
rect 37692 25052 37756 25056
rect 37692 24996 37696 25052
rect 37696 24996 37752 25052
rect 37752 24996 37756 25052
rect 37692 24992 37756 24996
rect 37772 25052 37836 25056
rect 37772 24996 37776 25052
rect 37776 24996 37832 25052
rect 37832 24996 37836 25052
rect 37772 24992 37836 24996
rect 37852 25052 37916 25056
rect 37852 24996 37856 25052
rect 37856 24996 37912 25052
rect 37912 24996 37916 25052
rect 37852 24992 37916 24996
rect 1952 24508 2016 24512
rect 1952 24452 1956 24508
rect 1956 24452 2012 24508
rect 2012 24452 2016 24508
rect 1952 24448 2016 24452
rect 2032 24508 2096 24512
rect 2032 24452 2036 24508
rect 2036 24452 2092 24508
rect 2092 24452 2096 24508
rect 2032 24448 2096 24452
rect 2112 24508 2176 24512
rect 2112 24452 2116 24508
rect 2116 24452 2172 24508
rect 2172 24452 2176 24508
rect 2112 24448 2176 24452
rect 2192 24508 2256 24512
rect 2192 24452 2196 24508
rect 2196 24452 2252 24508
rect 2252 24452 2256 24508
rect 2192 24448 2256 24452
rect 6952 24508 7016 24512
rect 6952 24452 6956 24508
rect 6956 24452 7012 24508
rect 7012 24452 7016 24508
rect 6952 24448 7016 24452
rect 7032 24508 7096 24512
rect 7032 24452 7036 24508
rect 7036 24452 7092 24508
rect 7092 24452 7096 24508
rect 7032 24448 7096 24452
rect 7112 24508 7176 24512
rect 7112 24452 7116 24508
rect 7116 24452 7172 24508
rect 7172 24452 7176 24508
rect 7112 24448 7176 24452
rect 7192 24508 7256 24512
rect 7192 24452 7196 24508
rect 7196 24452 7252 24508
rect 7252 24452 7256 24508
rect 7192 24448 7256 24452
rect 11952 24508 12016 24512
rect 11952 24452 11956 24508
rect 11956 24452 12012 24508
rect 12012 24452 12016 24508
rect 11952 24448 12016 24452
rect 12032 24508 12096 24512
rect 12032 24452 12036 24508
rect 12036 24452 12092 24508
rect 12092 24452 12096 24508
rect 12032 24448 12096 24452
rect 12112 24508 12176 24512
rect 12112 24452 12116 24508
rect 12116 24452 12172 24508
rect 12172 24452 12176 24508
rect 12112 24448 12176 24452
rect 12192 24508 12256 24512
rect 12192 24452 12196 24508
rect 12196 24452 12252 24508
rect 12252 24452 12256 24508
rect 12192 24448 12256 24452
rect 16952 24508 17016 24512
rect 16952 24452 16956 24508
rect 16956 24452 17012 24508
rect 17012 24452 17016 24508
rect 16952 24448 17016 24452
rect 17032 24508 17096 24512
rect 17032 24452 17036 24508
rect 17036 24452 17092 24508
rect 17092 24452 17096 24508
rect 17032 24448 17096 24452
rect 17112 24508 17176 24512
rect 17112 24452 17116 24508
rect 17116 24452 17172 24508
rect 17172 24452 17176 24508
rect 17112 24448 17176 24452
rect 17192 24508 17256 24512
rect 17192 24452 17196 24508
rect 17196 24452 17252 24508
rect 17252 24452 17256 24508
rect 17192 24448 17256 24452
rect 21952 24508 22016 24512
rect 21952 24452 21956 24508
rect 21956 24452 22012 24508
rect 22012 24452 22016 24508
rect 21952 24448 22016 24452
rect 22032 24508 22096 24512
rect 22032 24452 22036 24508
rect 22036 24452 22092 24508
rect 22092 24452 22096 24508
rect 22032 24448 22096 24452
rect 22112 24508 22176 24512
rect 22112 24452 22116 24508
rect 22116 24452 22172 24508
rect 22172 24452 22176 24508
rect 22112 24448 22176 24452
rect 22192 24508 22256 24512
rect 22192 24452 22196 24508
rect 22196 24452 22252 24508
rect 22252 24452 22256 24508
rect 22192 24448 22256 24452
rect 26952 24508 27016 24512
rect 26952 24452 26956 24508
rect 26956 24452 27012 24508
rect 27012 24452 27016 24508
rect 26952 24448 27016 24452
rect 27032 24508 27096 24512
rect 27032 24452 27036 24508
rect 27036 24452 27092 24508
rect 27092 24452 27096 24508
rect 27032 24448 27096 24452
rect 27112 24508 27176 24512
rect 27112 24452 27116 24508
rect 27116 24452 27172 24508
rect 27172 24452 27176 24508
rect 27112 24448 27176 24452
rect 27192 24508 27256 24512
rect 27192 24452 27196 24508
rect 27196 24452 27252 24508
rect 27252 24452 27256 24508
rect 27192 24448 27256 24452
rect 31952 24508 32016 24512
rect 31952 24452 31956 24508
rect 31956 24452 32012 24508
rect 32012 24452 32016 24508
rect 31952 24448 32016 24452
rect 32032 24508 32096 24512
rect 32032 24452 32036 24508
rect 32036 24452 32092 24508
rect 32092 24452 32096 24508
rect 32032 24448 32096 24452
rect 32112 24508 32176 24512
rect 32112 24452 32116 24508
rect 32116 24452 32172 24508
rect 32172 24452 32176 24508
rect 32112 24448 32176 24452
rect 32192 24508 32256 24512
rect 32192 24452 32196 24508
rect 32196 24452 32252 24508
rect 32252 24452 32256 24508
rect 32192 24448 32256 24452
rect 36952 24508 37016 24512
rect 36952 24452 36956 24508
rect 36956 24452 37012 24508
rect 37012 24452 37016 24508
rect 36952 24448 37016 24452
rect 37032 24508 37096 24512
rect 37032 24452 37036 24508
rect 37036 24452 37092 24508
rect 37092 24452 37096 24508
rect 37032 24448 37096 24452
rect 37112 24508 37176 24512
rect 37112 24452 37116 24508
rect 37116 24452 37172 24508
rect 37172 24452 37176 24508
rect 37112 24448 37176 24452
rect 37192 24508 37256 24512
rect 37192 24452 37196 24508
rect 37196 24452 37252 24508
rect 37252 24452 37256 24508
rect 37192 24448 37256 24452
rect 2612 23964 2676 23968
rect 2612 23908 2616 23964
rect 2616 23908 2672 23964
rect 2672 23908 2676 23964
rect 2612 23904 2676 23908
rect 2692 23964 2756 23968
rect 2692 23908 2696 23964
rect 2696 23908 2752 23964
rect 2752 23908 2756 23964
rect 2692 23904 2756 23908
rect 2772 23964 2836 23968
rect 2772 23908 2776 23964
rect 2776 23908 2832 23964
rect 2832 23908 2836 23964
rect 2772 23904 2836 23908
rect 2852 23964 2916 23968
rect 2852 23908 2856 23964
rect 2856 23908 2912 23964
rect 2912 23908 2916 23964
rect 2852 23904 2916 23908
rect 7612 23964 7676 23968
rect 7612 23908 7616 23964
rect 7616 23908 7672 23964
rect 7672 23908 7676 23964
rect 7612 23904 7676 23908
rect 7692 23964 7756 23968
rect 7692 23908 7696 23964
rect 7696 23908 7752 23964
rect 7752 23908 7756 23964
rect 7692 23904 7756 23908
rect 7772 23964 7836 23968
rect 7772 23908 7776 23964
rect 7776 23908 7832 23964
rect 7832 23908 7836 23964
rect 7772 23904 7836 23908
rect 7852 23964 7916 23968
rect 7852 23908 7856 23964
rect 7856 23908 7912 23964
rect 7912 23908 7916 23964
rect 7852 23904 7916 23908
rect 12612 23964 12676 23968
rect 12612 23908 12616 23964
rect 12616 23908 12672 23964
rect 12672 23908 12676 23964
rect 12612 23904 12676 23908
rect 12692 23964 12756 23968
rect 12692 23908 12696 23964
rect 12696 23908 12752 23964
rect 12752 23908 12756 23964
rect 12692 23904 12756 23908
rect 12772 23964 12836 23968
rect 12772 23908 12776 23964
rect 12776 23908 12832 23964
rect 12832 23908 12836 23964
rect 12772 23904 12836 23908
rect 12852 23964 12916 23968
rect 12852 23908 12856 23964
rect 12856 23908 12912 23964
rect 12912 23908 12916 23964
rect 12852 23904 12916 23908
rect 17612 23964 17676 23968
rect 17612 23908 17616 23964
rect 17616 23908 17672 23964
rect 17672 23908 17676 23964
rect 17612 23904 17676 23908
rect 17692 23964 17756 23968
rect 17692 23908 17696 23964
rect 17696 23908 17752 23964
rect 17752 23908 17756 23964
rect 17692 23904 17756 23908
rect 17772 23964 17836 23968
rect 17772 23908 17776 23964
rect 17776 23908 17832 23964
rect 17832 23908 17836 23964
rect 17772 23904 17836 23908
rect 17852 23964 17916 23968
rect 17852 23908 17856 23964
rect 17856 23908 17912 23964
rect 17912 23908 17916 23964
rect 17852 23904 17916 23908
rect 22612 23964 22676 23968
rect 22612 23908 22616 23964
rect 22616 23908 22672 23964
rect 22672 23908 22676 23964
rect 22612 23904 22676 23908
rect 22692 23964 22756 23968
rect 22692 23908 22696 23964
rect 22696 23908 22752 23964
rect 22752 23908 22756 23964
rect 22692 23904 22756 23908
rect 22772 23964 22836 23968
rect 22772 23908 22776 23964
rect 22776 23908 22832 23964
rect 22832 23908 22836 23964
rect 22772 23904 22836 23908
rect 22852 23964 22916 23968
rect 22852 23908 22856 23964
rect 22856 23908 22912 23964
rect 22912 23908 22916 23964
rect 22852 23904 22916 23908
rect 27612 23964 27676 23968
rect 27612 23908 27616 23964
rect 27616 23908 27672 23964
rect 27672 23908 27676 23964
rect 27612 23904 27676 23908
rect 27692 23964 27756 23968
rect 27692 23908 27696 23964
rect 27696 23908 27752 23964
rect 27752 23908 27756 23964
rect 27692 23904 27756 23908
rect 27772 23964 27836 23968
rect 27772 23908 27776 23964
rect 27776 23908 27832 23964
rect 27832 23908 27836 23964
rect 27772 23904 27836 23908
rect 27852 23964 27916 23968
rect 27852 23908 27856 23964
rect 27856 23908 27912 23964
rect 27912 23908 27916 23964
rect 27852 23904 27916 23908
rect 32612 23964 32676 23968
rect 32612 23908 32616 23964
rect 32616 23908 32672 23964
rect 32672 23908 32676 23964
rect 32612 23904 32676 23908
rect 32692 23964 32756 23968
rect 32692 23908 32696 23964
rect 32696 23908 32752 23964
rect 32752 23908 32756 23964
rect 32692 23904 32756 23908
rect 32772 23964 32836 23968
rect 32772 23908 32776 23964
rect 32776 23908 32832 23964
rect 32832 23908 32836 23964
rect 32772 23904 32836 23908
rect 32852 23964 32916 23968
rect 32852 23908 32856 23964
rect 32856 23908 32912 23964
rect 32912 23908 32916 23964
rect 32852 23904 32916 23908
rect 37612 23964 37676 23968
rect 37612 23908 37616 23964
rect 37616 23908 37672 23964
rect 37672 23908 37676 23964
rect 37612 23904 37676 23908
rect 37692 23964 37756 23968
rect 37692 23908 37696 23964
rect 37696 23908 37752 23964
rect 37752 23908 37756 23964
rect 37692 23904 37756 23908
rect 37772 23964 37836 23968
rect 37772 23908 37776 23964
rect 37776 23908 37832 23964
rect 37832 23908 37836 23964
rect 37772 23904 37836 23908
rect 37852 23964 37916 23968
rect 37852 23908 37856 23964
rect 37856 23908 37912 23964
rect 37912 23908 37916 23964
rect 37852 23904 37916 23908
rect 1952 23420 2016 23424
rect 1952 23364 1956 23420
rect 1956 23364 2012 23420
rect 2012 23364 2016 23420
rect 1952 23360 2016 23364
rect 2032 23420 2096 23424
rect 2032 23364 2036 23420
rect 2036 23364 2092 23420
rect 2092 23364 2096 23420
rect 2032 23360 2096 23364
rect 2112 23420 2176 23424
rect 2112 23364 2116 23420
rect 2116 23364 2172 23420
rect 2172 23364 2176 23420
rect 2112 23360 2176 23364
rect 2192 23420 2256 23424
rect 2192 23364 2196 23420
rect 2196 23364 2252 23420
rect 2252 23364 2256 23420
rect 2192 23360 2256 23364
rect 6952 23420 7016 23424
rect 6952 23364 6956 23420
rect 6956 23364 7012 23420
rect 7012 23364 7016 23420
rect 6952 23360 7016 23364
rect 7032 23420 7096 23424
rect 7032 23364 7036 23420
rect 7036 23364 7092 23420
rect 7092 23364 7096 23420
rect 7032 23360 7096 23364
rect 7112 23420 7176 23424
rect 7112 23364 7116 23420
rect 7116 23364 7172 23420
rect 7172 23364 7176 23420
rect 7112 23360 7176 23364
rect 7192 23420 7256 23424
rect 7192 23364 7196 23420
rect 7196 23364 7252 23420
rect 7252 23364 7256 23420
rect 7192 23360 7256 23364
rect 11952 23420 12016 23424
rect 11952 23364 11956 23420
rect 11956 23364 12012 23420
rect 12012 23364 12016 23420
rect 11952 23360 12016 23364
rect 12032 23420 12096 23424
rect 12032 23364 12036 23420
rect 12036 23364 12092 23420
rect 12092 23364 12096 23420
rect 12032 23360 12096 23364
rect 12112 23420 12176 23424
rect 12112 23364 12116 23420
rect 12116 23364 12172 23420
rect 12172 23364 12176 23420
rect 12112 23360 12176 23364
rect 12192 23420 12256 23424
rect 12192 23364 12196 23420
rect 12196 23364 12252 23420
rect 12252 23364 12256 23420
rect 12192 23360 12256 23364
rect 16952 23420 17016 23424
rect 16952 23364 16956 23420
rect 16956 23364 17012 23420
rect 17012 23364 17016 23420
rect 16952 23360 17016 23364
rect 17032 23420 17096 23424
rect 17032 23364 17036 23420
rect 17036 23364 17092 23420
rect 17092 23364 17096 23420
rect 17032 23360 17096 23364
rect 17112 23420 17176 23424
rect 17112 23364 17116 23420
rect 17116 23364 17172 23420
rect 17172 23364 17176 23420
rect 17112 23360 17176 23364
rect 17192 23420 17256 23424
rect 17192 23364 17196 23420
rect 17196 23364 17252 23420
rect 17252 23364 17256 23420
rect 17192 23360 17256 23364
rect 21952 23420 22016 23424
rect 21952 23364 21956 23420
rect 21956 23364 22012 23420
rect 22012 23364 22016 23420
rect 21952 23360 22016 23364
rect 22032 23420 22096 23424
rect 22032 23364 22036 23420
rect 22036 23364 22092 23420
rect 22092 23364 22096 23420
rect 22032 23360 22096 23364
rect 22112 23420 22176 23424
rect 22112 23364 22116 23420
rect 22116 23364 22172 23420
rect 22172 23364 22176 23420
rect 22112 23360 22176 23364
rect 22192 23420 22256 23424
rect 22192 23364 22196 23420
rect 22196 23364 22252 23420
rect 22252 23364 22256 23420
rect 22192 23360 22256 23364
rect 26952 23420 27016 23424
rect 26952 23364 26956 23420
rect 26956 23364 27012 23420
rect 27012 23364 27016 23420
rect 26952 23360 27016 23364
rect 27032 23420 27096 23424
rect 27032 23364 27036 23420
rect 27036 23364 27092 23420
rect 27092 23364 27096 23420
rect 27032 23360 27096 23364
rect 27112 23420 27176 23424
rect 27112 23364 27116 23420
rect 27116 23364 27172 23420
rect 27172 23364 27176 23420
rect 27112 23360 27176 23364
rect 27192 23420 27256 23424
rect 27192 23364 27196 23420
rect 27196 23364 27252 23420
rect 27252 23364 27256 23420
rect 27192 23360 27256 23364
rect 31952 23420 32016 23424
rect 31952 23364 31956 23420
rect 31956 23364 32012 23420
rect 32012 23364 32016 23420
rect 31952 23360 32016 23364
rect 32032 23420 32096 23424
rect 32032 23364 32036 23420
rect 32036 23364 32092 23420
rect 32092 23364 32096 23420
rect 32032 23360 32096 23364
rect 32112 23420 32176 23424
rect 32112 23364 32116 23420
rect 32116 23364 32172 23420
rect 32172 23364 32176 23420
rect 32112 23360 32176 23364
rect 32192 23420 32256 23424
rect 32192 23364 32196 23420
rect 32196 23364 32252 23420
rect 32252 23364 32256 23420
rect 32192 23360 32256 23364
rect 36952 23420 37016 23424
rect 36952 23364 36956 23420
rect 36956 23364 37012 23420
rect 37012 23364 37016 23420
rect 36952 23360 37016 23364
rect 37032 23420 37096 23424
rect 37032 23364 37036 23420
rect 37036 23364 37092 23420
rect 37092 23364 37096 23420
rect 37032 23360 37096 23364
rect 37112 23420 37176 23424
rect 37112 23364 37116 23420
rect 37116 23364 37172 23420
rect 37172 23364 37176 23420
rect 37112 23360 37176 23364
rect 37192 23420 37256 23424
rect 37192 23364 37196 23420
rect 37196 23364 37252 23420
rect 37252 23364 37256 23420
rect 37192 23360 37256 23364
rect 2612 22876 2676 22880
rect 2612 22820 2616 22876
rect 2616 22820 2672 22876
rect 2672 22820 2676 22876
rect 2612 22816 2676 22820
rect 2692 22876 2756 22880
rect 2692 22820 2696 22876
rect 2696 22820 2752 22876
rect 2752 22820 2756 22876
rect 2692 22816 2756 22820
rect 2772 22876 2836 22880
rect 2772 22820 2776 22876
rect 2776 22820 2832 22876
rect 2832 22820 2836 22876
rect 2772 22816 2836 22820
rect 2852 22876 2916 22880
rect 2852 22820 2856 22876
rect 2856 22820 2912 22876
rect 2912 22820 2916 22876
rect 2852 22816 2916 22820
rect 7612 22876 7676 22880
rect 7612 22820 7616 22876
rect 7616 22820 7672 22876
rect 7672 22820 7676 22876
rect 7612 22816 7676 22820
rect 7692 22876 7756 22880
rect 7692 22820 7696 22876
rect 7696 22820 7752 22876
rect 7752 22820 7756 22876
rect 7692 22816 7756 22820
rect 7772 22876 7836 22880
rect 7772 22820 7776 22876
rect 7776 22820 7832 22876
rect 7832 22820 7836 22876
rect 7772 22816 7836 22820
rect 7852 22876 7916 22880
rect 7852 22820 7856 22876
rect 7856 22820 7912 22876
rect 7912 22820 7916 22876
rect 7852 22816 7916 22820
rect 12612 22876 12676 22880
rect 12612 22820 12616 22876
rect 12616 22820 12672 22876
rect 12672 22820 12676 22876
rect 12612 22816 12676 22820
rect 12692 22876 12756 22880
rect 12692 22820 12696 22876
rect 12696 22820 12752 22876
rect 12752 22820 12756 22876
rect 12692 22816 12756 22820
rect 12772 22876 12836 22880
rect 12772 22820 12776 22876
rect 12776 22820 12832 22876
rect 12832 22820 12836 22876
rect 12772 22816 12836 22820
rect 12852 22876 12916 22880
rect 12852 22820 12856 22876
rect 12856 22820 12912 22876
rect 12912 22820 12916 22876
rect 12852 22816 12916 22820
rect 17612 22876 17676 22880
rect 17612 22820 17616 22876
rect 17616 22820 17672 22876
rect 17672 22820 17676 22876
rect 17612 22816 17676 22820
rect 17692 22876 17756 22880
rect 17692 22820 17696 22876
rect 17696 22820 17752 22876
rect 17752 22820 17756 22876
rect 17692 22816 17756 22820
rect 17772 22876 17836 22880
rect 17772 22820 17776 22876
rect 17776 22820 17832 22876
rect 17832 22820 17836 22876
rect 17772 22816 17836 22820
rect 17852 22876 17916 22880
rect 17852 22820 17856 22876
rect 17856 22820 17912 22876
rect 17912 22820 17916 22876
rect 17852 22816 17916 22820
rect 22612 22876 22676 22880
rect 22612 22820 22616 22876
rect 22616 22820 22672 22876
rect 22672 22820 22676 22876
rect 22612 22816 22676 22820
rect 22692 22876 22756 22880
rect 22692 22820 22696 22876
rect 22696 22820 22752 22876
rect 22752 22820 22756 22876
rect 22692 22816 22756 22820
rect 22772 22876 22836 22880
rect 22772 22820 22776 22876
rect 22776 22820 22832 22876
rect 22832 22820 22836 22876
rect 22772 22816 22836 22820
rect 22852 22876 22916 22880
rect 22852 22820 22856 22876
rect 22856 22820 22912 22876
rect 22912 22820 22916 22876
rect 22852 22816 22916 22820
rect 27612 22876 27676 22880
rect 27612 22820 27616 22876
rect 27616 22820 27672 22876
rect 27672 22820 27676 22876
rect 27612 22816 27676 22820
rect 27692 22876 27756 22880
rect 27692 22820 27696 22876
rect 27696 22820 27752 22876
rect 27752 22820 27756 22876
rect 27692 22816 27756 22820
rect 27772 22876 27836 22880
rect 27772 22820 27776 22876
rect 27776 22820 27832 22876
rect 27832 22820 27836 22876
rect 27772 22816 27836 22820
rect 27852 22876 27916 22880
rect 27852 22820 27856 22876
rect 27856 22820 27912 22876
rect 27912 22820 27916 22876
rect 27852 22816 27916 22820
rect 32612 22876 32676 22880
rect 32612 22820 32616 22876
rect 32616 22820 32672 22876
rect 32672 22820 32676 22876
rect 32612 22816 32676 22820
rect 32692 22876 32756 22880
rect 32692 22820 32696 22876
rect 32696 22820 32752 22876
rect 32752 22820 32756 22876
rect 32692 22816 32756 22820
rect 32772 22876 32836 22880
rect 32772 22820 32776 22876
rect 32776 22820 32832 22876
rect 32832 22820 32836 22876
rect 32772 22816 32836 22820
rect 32852 22876 32916 22880
rect 32852 22820 32856 22876
rect 32856 22820 32912 22876
rect 32912 22820 32916 22876
rect 32852 22816 32916 22820
rect 37612 22876 37676 22880
rect 37612 22820 37616 22876
rect 37616 22820 37672 22876
rect 37672 22820 37676 22876
rect 37612 22816 37676 22820
rect 37692 22876 37756 22880
rect 37692 22820 37696 22876
rect 37696 22820 37752 22876
rect 37752 22820 37756 22876
rect 37692 22816 37756 22820
rect 37772 22876 37836 22880
rect 37772 22820 37776 22876
rect 37776 22820 37832 22876
rect 37832 22820 37836 22876
rect 37772 22816 37836 22820
rect 37852 22876 37916 22880
rect 37852 22820 37856 22876
rect 37856 22820 37912 22876
rect 37912 22820 37916 22876
rect 37852 22816 37916 22820
rect 21036 22612 21100 22676
rect 1952 22332 2016 22336
rect 1952 22276 1956 22332
rect 1956 22276 2012 22332
rect 2012 22276 2016 22332
rect 1952 22272 2016 22276
rect 2032 22332 2096 22336
rect 2032 22276 2036 22332
rect 2036 22276 2092 22332
rect 2092 22276 2096 22332
rect 2032 22272 2096 22276
rect 2112 22332 2176 22336
rect 2112 22276 2116 22332
rect 2116 22276 2172 22332
rect 2172 22276 2176 22332
rect 2112 22272 2176 22276
rect 2192 22332 2256 22336
rect 2192 22276 2196 22332
rect 2196 22276 2252 22332
rect 2252 22276 2256 22332
rect 2192 22272 2256 22276
rect 6952 22332 7016 22336
rect 6952 22276 6956 22332
rect 6956 22276 7012 22332
rect 7012 22276 7016 22332
rect 6952 22272 7016 22276
rect 7032 22332 7096 22336
rect 7032 22276 7036 22332
rect 7036 22276 7092 22332
rect 7092 22276 7096 22332
rect 7032 22272 7096 22276
rect 7112 22332 7176 22336
rect 7112 22276 7116 22332
rect 7116 22276 7172 22332
rect 7172 22276 7176 22332
rect 7112 22272 7176 22276
rect 7192 22332 7256 22336
rect 7192 22276 7196 22332
rect 7196 22276 7252 22332
rect 7252 22276 7256 22332
rect 7192 22272 7256 22276
rect 11952 22332 12016 22336
rect 11952 22276 11956 22332
rect 11956 22276 12012 22332
rect 12012 22276 12016 22332
rect 11952 22272 12016 22276
rect 12032 22332 12096 22336
rect 12032 22276 12036 22332
rect 12036 22276 12092 22332
rect 12092 22276 12096 22332
rect 12032 22272 12096 22276
rect 12112 22332 12176 22336
rect 12112 22276 12116 22332
rect 12116 22276 12172 22332
rect 12172 22276 12176 22332
rect 12112 22272 12176 22276
rect 12192 22332 12256 22336
rect 12192 22276 12196 22332
rect 12196 22276 12252 22332
rect 12252 22276 12256 22332
rect 12192 22272 12256 22276
rect 16952 22332 17016 22336
rect 16952 22276 16956 22332
rect 16956 22276 17012 22332
rect 17012 22276 17016 22332
rect 16952 22272 17016 22276
rect 17032 22332 17096 22336
rect 17032 22276 17036 22332
rect 17036 22276 17092 22332
rect 17092 22276 17096 22332
rect 17032 22272 17096 22276
rect 17112 22332 17176 22336
rect 17112 22276 17116 22332
rect 17116 22276 17172 22332
rect 17172 22276 17176 22332
rect 17112 22272 17176 22276
rect 17192 22332 17256 22336
rect 17192 22276 17196 22332
rect 17196 22276 17252 22332
rect 17252 22276 17256 22332
rect 17192 22272 17256 22276
rect 21952 22332 22016 22336
rect 21952 22276 21956 22332
rect 21956 22276 22012 22332
rect 22012 22276 22016 22332
rect 21952 22272 22016 22276
rect 22032 22332 22096 22336
rect 22032 22276 22036 22332
rect 22036 22276 22092 22332
rect 22092 22276 22096 22332
rect 22032 22272 22096 22276
rect 22112 22332 22176 22336
rect 22112 22276 22116 22332
rect 22116 22276 22172 22332
rect 22172 22276 22176 22332
rect 22112 22272 22176 22276
rect 22192 22332 22256 22336
rect 22192 22276 22196 22332
rect 22196 22276 22252 22332
rect 22252 22276 22256 22332
rect 22192 22272 22256 22276
rect 26952 22332 27016 22336
rect 26952 22276 26956 22332
rect 26956 22276 27012 22332
rect 27012 22276 27016 22332
rect 26952 22272 27016 22276
rect 27032 22332 27096 22336
rect 27032 22276 27036 22332
rect 27036 22276 27092 22332
rect 27092 22276 27096 22332
rect 27032 22272 27096 22276
rect 27112 22332 27176 22336
rect 27112 22276 27116 22332
rect 27116 22276 27172 22332
rect 27172 22276 27176 22332
rect 27112 22272 27176 22276
rect 27192 22332 27256 22336
rect 27192 22276 27196 22332
rect 27196 22276 27252 22332
rect 27252 22276 27256 22332
rect 27192 22272 27256 22276
rect 31952 22332 32016 22336
rect 31952 22276 31956 22332
rect 31956 22276 32012 22332
rect 32012 22276 32016 22332
rect 31952 22272 32016 22276
rect 32032 22332 32096 22336
rect 32032 22276 32036 22332
rect 32036 22276 32092 22332
rect 32092 22276 32096 22332
rect 32032 22272 32096 22276
rect 32112 22332 32176 22336
rect 32112 22276 32116 22332
rect 32116 22276 32172 22332
rect 32172 22276 32176 22332
rect 32112 22272 32176 22276
rect 32192 22332 32256 22336
rect 32192 22276 32196 22332
rect 32196 22276 32252 22332
rect 32252 22276 32256 22332
rect 32192 22272 32256 22276
rect 36952 22332 37016 22336
rect 36952 22276 36956 22332
rect 36956 22276 37012 22332
rect 37012 22276 37016 22332
rect 36952 22272 37016 22276
rect 37032 22332 37096 22336
rect 37032 22276 37036 22332
rect 37036 22276 37092 22332
rect 37092 22276 37096 22332
rect 37032 22272 37096 22276
rect 37112 22332 37176 22336
rect 37112 22276 37116 22332
rect 37116 22276 37172 22332
rect 37172 22276 37176 22332
rect 37112 22272 37176 22276
rect 37192 22332 37256 22336
rect 37192 22276 37196 22332
rect 37196 22276 37252 22332
rect 37252 22276 37256 22332
rect 37192 22272 37256 22276
rect 21036 21932 21100 21996
rect 2612 21788 2676 21792
rect 2612 21732 2616 21788
rect 2616 21732 2672 21788
rect 2672 21732 2676 21788
rect 2612 21728 2676 21732
rect 2692 21788 2756 21792
rect 2692 21732 2696 21788
rect 2696 21732 2752 21788
rect 2752 21732 2756 21788
rect 2692 21728 2756 21732
rect 2772 21788 2836 21792
rect 2772 21732 2776 21788
rect 2776 21732 2832 21788
rect 2832 21732 2836 21788
rect 2772 21728 2836 21732
rect 2852 21788 2916 21792
rect 2852 21732 2856 21788
rect 2856 21732 2912 21788
rect 2912 21732 2916 21788
rect 2852 21728 2916 21732
rect 7612 21788 7676 21792
rect 7612 21732 7616 21788
rect 7616 21732 7672 21788
rect 7672 21732 7676 21788
rect 7612 21728 7676 21732
rect 7692 21788 7756 21792
rect 7692 21732 7696 21788
rect 7696 21732 7752 21788
rect 7752 21732 7756 21788
rect 7692 21728 7756 21732
rect 7772 21788 7836 21792
rect 7772 21732 7776 21788
rect 7776 21732 7832 21788
rect 7832 21732 7836 21788
rect 7772 21728 7836 21732
rect 7852 21788 7916 21792
rect 7852 21732 7856 21788
rect 7856 21732 7912 21788
rect 7912 21732 7916 21788
rect 7852 21728 7916 21732
rect 12612 21788 12676 21792
rect 12612 21732 12616 21788
rect 12616 21732 12672 21788
rect 12672 21732 12676 21788
rect 12612 21728 12676 21732
rect 12692 21788 12756 21792
rect 12692 21732 12696 21788
rect 12696 21732 12752 21788
rect 12752 21732 12756 21788
rect 12692 21728 12756 21732
rect 12772 21788 12836 21792
rect 12772 21732 12776 21788
rect 12776 21732 12832 21788
rect 12832 21732 12836 21788
rect 12772 21728 12836 21732
rect 12852 21788 12916 21792
rect 12852 21732 12856 21788
rect 12856 21732 12912 21788
rect 12912 21732 12916 21788
rect 12852 21728 12916 21732
rect 17612 21788 17676 21792
rect 17612 21732 17616 21788
rect 17616 21732 17672 21788
rect 17672 21732 17676 21788
rect 17612 21728 17676 21732
rect 17692 21788 17756 21792
rect 17692 21732 17696 21788
rect 17696 21732 17752 21788
rect 17752 21732 17756 21788
rect 17692 21728 17756 21732
rect 17772 21788 17836 21792
rect 17772 21732 17776 21788
rect 17776 21732 17832 21788
rect 17832 21732 17836 21788
rect 17772 21728 17836 21732
rect 17852 21788 17916 21792
rect 17852 21732 17856 21788
rect 17856 21732 17912 21788
rect 17912 21732 17916 21788
rect 17852 21728 17916 21732
rect 22612 21788 22676 21792
rect 22612 21732 22616 21788
rect 22616 21732 22672 21788
rect 22672 21732 22676 21788
rect 22612 21728 22676 21732
rect 22692 21788 22756 21792
rect 22692 21732 22696 21788
rect 22696 21732 22752 21788
rect 22752 21732 22756 21788
rect 22692 21728 22756 21732
rect 22772 21788 22836 21792
rect 22772 21732 22776 21788
rect 22776 21732 22832 21788
rect 22832 21732 22836 21788
rect 22772 21728 22836 21732
rect 22852 21788 22916 21792
rect 22852 21732 22856 21788
rect 22856 21732 22912 21788
rect 22912 21732 22916 21788
rect 22852 21728 22916 21732
rect 27612 21788 27676 21792
rect 27612 21732 27616 21788
rect 27616 21732 27672 21788
rect 27672 21732 27676 21788
rect 27612 21728 27676 21732
rect 27692 21788 27756 21792
rect 27692 21732 27696 21788
rect 27696 21732 27752 21788
rect 27752 21732 27756 21788
rect 27692 21728 27756 21732
rect 27772 21788 27836 21792
rect 27772 21732 27776 21788
rect 27776 21732 27832 21788
rect 27832 21732 27836 21788
rect 27772 21728 27836 21732
rect 27852 21788 27916 21792
rect 27852 21732 27856 21788
rect 27856 21732 27912 21788
rect 27912 21732 27916 21788
rect 27852 21728 27916 21732
rect 32612 21788 32676 21792
rect 32612 21732 32616 21788
rect 32616 21732 32672 21788
rect 32672 21732 32676 21788
rect 32612 21728 32676 21732
rect 32692 21788 32756 21792
rect 32692 21732 32696 21788
rect 32696 21732 32752 21788
rect 32752 21732 32756 21788
rect 32692 21728 32756 21732
rect 32772 21788 32836 21792
rect 32772 21732 32776 21788
rect 32776 21732 32832 21788
rect 32832 21732 32836 21788
rect 32772 21728 32836 21732
rect 32852 21788 32916 21792
rect 32852 21732 32856 21788
rect 32856 21732 32912 21788
rect 32912 21732 32916 21788
rect 32852 21728 32916 21732
rect 37612 21788 37676 21792
rect 37612 21732 37616 21788
rect 37616 21732 37672 21788
rect 37672 21732 37676 21788
rect 37612 21728 37676 21732
rect 37692 21788 37756 21792
rect 37692 21732 37696 21788
rect 37696 21732 37752 21788
rect 37752 21732 37756 21788
rect 37692 21728 37756 21732
rect 37772 21788 37836 21792
rect 37772 21732 37776 21788
rect 37776 21732 37832 21788
rect 37832 21732 37836 21788
rect 37772 21728 37836 21732
rect 37852 21788 37916 21792
rect 37852 21732 37856 21788
rect 37856 21732 37912 21788
rect 37912 21732 37916 21788
rect 37852 21728 37916 21732
rect 1952 21244 2016 21248
rect 1952 21188 1956 21244
rect 1956 21188 2012 21244
rect 2012 21188 2016 21244
rect 1952 21184 2016 21188
rect 2032 21244 2096 21248
rect 2032 21188 2036 21244
rect 2036 21188 2092 21244
rect 2092 21188 2096 21244
rect 2032 21184 2096 21188
rect 2112 21244 2176 21248
rect 2112 21188 2116 21244
rect 2116 21188 2172 21244
rect 2172 21188 2176 21244
rect 2112 21184 2176 21188
rect 2192 21244 2256 21248
rect 2192 21188 2196 21244
rect 2196 21188 2252 21244
rect 2252 21188 2256 21244
rect 2192 21184 2256 21188
rect 6952 21244 7016 21248
rect 6952 21188 6956 21244
rect 6956 21188 7012 21244
rect 7012 21188 7016 21244
rect 6952 21184 7016 21188
rect 7032 21244 7096 21248
rect 7032 21188 7036 21244
rect 7036 21188 7092 21244
rect 7092 21188 7096 21244
rect 7032 21184 7096 21188
rect 7112 21244 7176 21248
rect 7112 21188 7116 21244
rect 7116 21188 7172 21244
rect 7172 21188 7176 21244
rect 7112 21184 7176 21188
rect 7192 21244 7256 21248
rect 7192 21188 7196 21244
rect 7196 21188 7252 21244
rect 7252 21188 7256 21244
rect 7192 21184 7256 21188
rect 11952 21244 12016 21248
rect 11952 21188 11956 21244
rect 11956 21188 12012 21244
rect 12012 21188 12016 21244
rect 11952 21184 12016 21188
rect 12032 21244 12096 21248
rect 12032 21188 12036 21244
rect 12036 21188 12092 21244
rect 12092 21188 12096 21244
rect 12032 21184 12096 21188
rect 12112 21244 12176 21248
rect 12112 21188 12116 21244
rect 12116 21188 12172 21244
rect 12172 21188 12176 21244
rect 12112 21184 12176 21188
rect 12192 21244 12256 21248
rect 12192 21188 12196 21244
rect 12196 21188 12252 21244
rect 12252 21188 12256 21244
rect 12192 21184 12256 21188
rect 16952 21244 17016 21248
rect 16952 21188 16956 21244
rect 16956 21188 17012 21244
rect 17012 21188 17016 21244
rect 16952 21184 17016 21188
rect 17032 21244 17096 21248
rect 17032 21188 17036 21244
rect 17036 21188 17092 21244
rect 17092 21188 17096 21244
rect 17032 21184 17096 21188
rect 17112 21244 17176 21248
rect 17112 21188 17116 21244
rect 17116 21188 17172 21244
rect 17172 21188 17176 21244
rect 17112 21184 17176 21188
rect 17192 21244 17256 21248
rect 17192 21188 17196 21244
rect 17196 21188 17252 21244
rect 17252 21188 17256 21244
rect 17192 21184 17256 21188
rect 21952 21244 22016 21248
rect 21952 21188 21956 21244
rect 21956 21188 22012 21244
rect 22012 21188 22016 21244
rect 21952 21184 22016 21188
rect 22032 21244 22096 21248
rect 22032 21188 22036 21244
rect 22036 21188 22092 21244
rect 22092 21188 22096 21244
rect 22032 21184 22096 21188
rect 22112 21244 22176 21248
rect 22112 21188 22116 21244
rect 22116 21188 22172 21244
rect 22172 21188 22176 21244
rect 22112 21184 22176 21188
rect 22192 21244 22256 21248
rect 22192 21188 22196 21244
rect 22196 21188 22252 21244
rect 22252 21188 22256 21244
rect 22192 21184 22256 21188
rect 26952 21244 27016 21248
rect 26952 21188 26956 21244
rect 26956 21188 27012 21244
rect 27012 21188 27016 21244
rect 26952 21184 27016 21188
rect 27032 21244 27096 21248
rect 27032 21188 27036 21244
rect 27036 21188 27092 21244
rect 27092 21188 27096 21244
rect 27032 21184 27096 21188
rect 27112 21244 27176 21248
rect 27112 21188 27116 21244
rect 27116 21188 27172 21244
rect 27172 21188 27176 21244
rect 27112 21184 27176 21188
rect 27192 21244 27256 21248
rect 27192 21188 27196 21244
rect 27196 21188 27252 21244
rect 27252 21188 27256 21244
rect 27192 21184 27256 21188
rect 31952 21244 32016 21248
rect 31952 21188 31956 21244
rect 31956 21188 32012 21244
rect 32012 21188 32016 21244
rect 31952 21184 32016 21188
rect 32032 21244 32096 21248
rect 32032 21188 32036 21244
rect 32036 21188 32092 21244
rect 32092 21188 32096 21244
rect 32032 21184 32096 21188
rect 32112 21244 32176 21248
rect 32112 21188 32116 21244
rect 32116 21188 32172 21244
rect 32172 21188 32176 21244
rect 32112 21184 32176 21188
rect 32192 21244 32256 21248
rect 32192 21188 32196 21244
rect 32196 21188 32252 21244
rect 32252 21188 32256 21244
rect 32192 21184 32256 21188
rect 36952 21244 37016 21248
rect 36952 21188 36956 21244
rect 36956 21188 37012 21244
rect 37012 21188 37016 21244
rect 36952 21184 37016 21188
rect 37032 21244 37096 21248
rect 37032 21188 37036 21244
rect 37036 21188 37092 21244
rect 37092 21188 37096 21244
rect 37032 21184 37096 21188
rect 37112 21244 37176 21248
rect 37112 21188 37116 21244
rect 37116 21188 37172 21244
rect 37172 21188 37176 21244
rect 37112 21184 37176 21188
rect 37192 21244 37256 21248
rect 37192 21188 37196 21244
rect 37196 21188 37252 21244
rect 37252 21188 37256 21244
rect 37192 21184 37256 21188
rect 2612 20700 2676 20704
rect 2612 20644 2616 20700
rect 2616 20644 2672 20700
rect 2672 20644 2676 20700
rect 2612 20640 2676 20644
rect 2692 20700 2756 20704
rect 2692 20644 2696 20700
rect 2696 20644 2752 20700
rect 2752 20644 2756 20700
rect 2692 20640 2756 20644
rect 2772 20700 2836 20704
rect 2772 20644 2776 20700
rect 2776 20644 2832 20700
rect 2832 20644 2836 20700
rect 2772 20640 2836 20644
rect 2852 20700 2916 20704
rect 2852 20644 2856 20700
rect 2856 20644 2912 20700
rect 2912 20644 2916 20700
rect 2852 20640 2916 20644
rect 7612 20700 7676 20704
rect 7612 20644 7616 20700
rect 7616 20644 7672 20700
rect 7672 20644 7676 20700
rect 7612 20640 7676 20644
rect 7692 20700 7756 20704
rect 7692 20644 7696 20700
rect 7696 20644 7752 20700
rect 7752 20644 7756 20700
rect 7692 20640 7756 20644
rect 7772 20700 7836 20704
rect 7772 20644 7776 20700
rect 7776 20644 7832 20700
rect 7832 20644 7836 20700
rect 7772 20640 7836 20644
rect 7852 20700 7916 20704
rect 7852 20644 7856 20700
rect 7856 20644 7912 20700
rect 7912 20644 7916 20700
rect 7852 20640 7916 20644
rect 12612 20700 12676 20704
rect 12612 20644 12616 20700
rect 12616 20644 12672 20700
rect 12672 20644 12676 20700
rect 12612 20640 12676 20644
rect 12692 20700 12756 20704
rect 12692 20644 12696 20700
rect 12696 20644 12752 20700
rect 12752 20644 12756 20700
rect 12692 20640 12756 20644
rect 12772 20700 12836 20704
rect 12772 20644 12776 20700
rect 12776 20644 12832 20700
rect 12832 20644 12836 20700
rect 12772 20640 12836 20644
rect 12852 20700 12916 20704
rect 12852 20644 12856 20700
rect 12856 20644 12912 20700
rect 12912 20644 12916 20700
rect 12852 20640 12916 20644
rect 17612 20700 17676 20704
rect 17612 20644 17616 20700
rect 17616 20644 17672 20700
rect 17672 20644 17676 20700
rect 17612 20640 17676 20644
rect 17692 20700 17756 20704
rect 17692 20644 17696 20700
rect 17696 20644 17752 20700
rect 17752 20644 17756 20700
rect 17692 20640 17756 20644
rect 17772 20700 17836 20704
rect 17772 20644 17776 20700
rect 17776 20644 17832 20700
rect 17832 20644 17836 20700
rect 17772 20640 17836 20644
rect 17852 20700 17916 20704
rect 17852 20644 17856 20700
rect 17856 20644 17912 20700
rect 17912 20644 17916 20700
rect 17852 20640 17916 20644
rect 22612 20700 22676 20704
rect 22612 20644 22616 20700
rect 22616 20644 22672 20700
rect 22672 20644 22676 20700
rect 22612 20640 22676 20644
rect 22692 20700 22756 20704
rect 22692 20644 22696 20700
rect 22696 20644 22752 20700
rect 22752 20644 22756 20700
rect 22692 20640 22756 20644
rect 22772 20700 22836 20704
rect 22772 20644 22776 20700
rect 22776 20644 22832 20700
rect 22832 20644 22836 20700
rect 22772 20640 22836 20644
rect 22852 20700 22916 20704
rect 22852 20644 22856 20700
rect 22856 20644 22912 20700
rect 22912 20644 22916 20700
rect 22852 20640 22916 20644
rect 27612 20700 27676 20704
rect 27612 20644 27616 20700
rect 27616 20644 27672 20700
rect 27672 20644 27676 20700
rect 27612 20640 27676 20644
rect 27692 20700 27756 20704
rect 27692 20644 27696 20700
rect 27696 20644 27752 20700
rect 27752 20644 27756 20700
rect 27692 20640 27756 20644
rect 27772 20700 27836 20704
rect 27772 20644 27776 20700
rect 27776 20644 27832 20700
rect 27832 20644 27836 20700
rect 27772 20640 27836 20644
rect 27852 20700 27916 20704
rect 27852 20644 27856 20700
rect 27856 20644 27912 20700
rect 27912 20644 27916 20700
rect 27852 20640 27916 20644
rect 32612 20700 32676 20704
rect 32612 20644 32616 20700
rect 32616 20644 32672 20700
rect 32672 20644 32676 20700
rect 32612 20640 32676 20644
rect 32692 20700 32756 20704
rect 32692 20644 32696 20700
rect 32696 20644 32752 20700
rect 32752 20644 32756 20700
rect 32692 20640 32756 20644
rect 32772 20700 32836 20704
rect 32772 20644 32776 20700
rect 32776 20644 32832 20700
rect 32832 20644 32836 20700
rect 32772 20640 32836 20644
rect 32852 20700 32916 20704
rect 32852 20644 32856 20700
rect 32856 20644 32912 20700
rect 32912 20644 32916 20700
rect 32852 20640 32916 20644
rect 37612 20700 37676 20704
rect 37612 20644 37616 20700
rect 37616 20644 37672 20700
rect 37672 20644 37676 20700
rect 37612 20640 37676 20644
rect 37692 20700 37756 20704
rect 37692 20644 37696 20700
rect 37696 20644 37752 20700
rect 37752 20644 37756 20700
rect 37692 20640 37756 20644
rect 37772 20700 37836 20704
rect 37772 20644 37776 20700
rect 37776 20644 37832 20700
rect 37832 20644 37836 20700
rect 37772 20640 37836 20644
rect 37852 20700 37916 20704
rect 37852 20644 37856 20700
rect 37856 20644 37912 20700
rect 37912 20644 37916 20700
rect 37852 20640 37916 20644
rect 1952 20156 2016 20160
rect 1952 20100 1956 20156
rect 1956 20100 2012 20156
rect 2012 20100 2016 20156
rect 1952 20096 2016 20100
rect 2032 20156 2096 20160
rect 2032 20100 2036 20156
rect 2036 20100 2092 20156
rect 2092 20100 2096 20156
rect 2032 20096 2096 20100
rect 2112 20156 2176 20160
rect 2112 20100 2116 20156
rect 2116 20100 2172 20156
rect 2172 20100 2176 20156
rect 2112 20096 2176 20100
rect 2192 20156 2256 20160
rect 2192 20100 2196 20156
rect 2196 20100 2252 20156
rect 2252 20100 2256 20156
rect 2192 20096 2256 20100
rect 6952 20156 7016 20160
rect 6952 20100 6956 20156
rect 6956 20100 7012 20156
rect 7012 20100 7016 20156
rect 6952 20096 7016 20100
rect 7032 20156 7096 20160
rect 7032 20100 7036 20156
rect 7036 20100 7092 20156
rect 7092 20100 7096 20156
rect 7032 20096 7096 20100
rect 7112 20156 7176 20160
rect 7112 20100 7116 20156
rect 7116 20100 7172 20156
rect 7172 20100 7176 20156
rect 7112 20096 7176 20100
rect 7192 20156 7256 20160
rect 7192 20100 7196 20156
rect 7196 20100 7252 20156
rect 7252 20100 7256 20156
rect 7192 20096 7256 20100
rect 11952 20156 12016 20160
rect 11952 20100 11956 20156
rect 11956 20100 12012 20156
rect 12012 20100 12016 20156
rect 11952 20096 12016 20100
rect 12032 20156 12096 20160
rect 12032 20100 12036 20156
rect 12036 20100 12092 20156
rect 12092 20100 12096 20156
rect 12032 20096 12096 20100
rect 12112 20156 12176 20160
rect 12112 20100 12116 20156
rect 12116 20100 12172 20156
rect 12172 20100 12176 20156
rect 12112 20096 12176 20100
rect 12192 20156 12256 20160
rect 12192 20100 12196 20156
rect 12196 20100 12252 20156
rect 12252 20100 12256 20156
rect 12192 20096 12256 20100
rect 16952 20156 17016 20160
rect 16952 20100 16956 20156
rect 16956 20100 17012 20156
rect 17012 20100 17016 20156
rect 16952 20096 17016 20100
rect 17032 20156 17096 20160
rect 17032 20100 17036 20156
rect 17036 20100 17092 20156
rect 17092 20100 17096 20156
rect 17032 20096 17096 20100
rect 17112 20156 17176 20160
rect 17112 20100 17116 20156
rect 17116 20100 17172 20156
rect 17172 20100 17176 20156
rect 17112 20096 17176 20100
rect 17192 20156 17256 20160
rect 17192 20100 17196 20156
rect 17196 20100 17252 20156
rect 17252 20100 17256 20156
rect 17192 20096 17256 20100
rect 21952 20156 22016 20160
rect 21952 20100 21956 20156
rect 21956 20100 22012 20156
rect 22012 20100 22016 20156
rect 21952 20096 22016 20100
rect 22032 20156 22096 20160
rect 22032 20100 22036 20156
rect 22036 20100 22092 20156
rect 22092 20100 22096 20156
rect 22032 20096 22096 20100
rect 22112 20156 22176 20160
rect 22112 20100 22116 20156
rect 22116 20100 22172 20156
rect 22172 20100 22176 20156
rect 22112 20096 22176 20100
rect 22192 20156 22256 20160
rect 22192 20100 22196 20156
rect 22196 20100 22252 20156
rect 22252 20100 22256 20156
rect 22192 20096 22256 20100
rect 26952 20156 27016 20160
rect 26952 20100 26956 20156
rect 26956 20100 27012 20156
rect 27012 20100 27016 20156
rect 26952 20096 27016 20100
rect 27032 20156 27096 20160
rect 27032 20100 27036 20156
rect 27036 20100 27092 20156
rect 27092 20100 27096 20156
rect 27032 20096 27096 20100
rect 27112 20156 27176 20160
rect 27112 20100 27116 20156
rect 27116 20100 27172 20156
rect 27172 20100 27176 20156
rect 27112 20096 27176 20100
rect 27192 20156 27256 20160
rect 27192 20100 27196 20156
rect 27196 20100 27252 20156
rect 27252 20100 27256 20156
rect 27192 20096 27256 20100
rect 31952 20156 32016 20160
rect 31952 20100 31956 20156
rect 31956 20100 32012 20156
rect 32012 20100 32016 20156
rect 31952 20096 32016 20100
rect 32032 20156 32096 20160
rect 32032 20100 32036 20156
rect 32036 20100 32092 20156
rect 32092 20100 32096 20156
rect 32032 20096 32096 20100
rect 32112 20156 32176 20160
rect 32112 20100 32116 20156
rect 32116 20100 32172 20156
rect 32172 20100 32176 20156
rect 32112 20096 32176 20100
rect 32192 20156 32256 20160
rect 32192 20100 32196 20156
rect 32196 20100 32252 20156
rect 32252 20100 32256 20156
rect 32192 20096 32256 20100
rect 36952 20156 37016 20160
rect 36952 20100 36956 20156
rect 36956 20100 37012 20156
rect 37012 20100 37016 20156
rect 36952 20096 37016 20100
rect 37032 20156 37096 20160
rect 37032 20100 37036 20156
rect 37036 20100 37092 20156
rect 37092 20100 37096 20156
rect 37032 20096 37096 20100
rect 37112 20156 37176 20160
rect 37112 20100 37116 20156
rect 37116 20100 37172 20156
rect 37172 20100 37176 20156
rect 37112 20096 37176 20100
rect 37192 20156 37256 20160
rect 37192 20100 37196 20156
rect 37196 20100 37252 20156
rect 37252 20100 37256 20156
rect 37192 20096 37256 20100
rect 2612 19612 2676 19616
rect 2612 19556 2616 19612
rect 2616 19556 2672 19612
rect 2672 19556 2676 19612
rect 2612 19552 2676 19556
rect 2692 19612 2756 19616
rect 2692 19556 2696 19612
rect 2696 19556 2752 19612
rect 2752 19556 2756 19612
rect 2692 19552 2756 19556
rect 2772 19612 2836 19616
rect 2772 19556 2776 19612
rect 2776 19556 2832 19612
rect 2832 19556 2836 19612
rect 2772 19552 2836 19556
rect 2852 19612 2916 19616
rect 2852 19556 2856 19612
rect 2856 19556 2912 19612
rect 2912 19556 2916 19612
rect 2852 19552 2916 19556
rect 7612 19612 7676 19616
rect 7612 19556 7616 19612
rect 7616 19556 7672 19612
rect 7672 19556 7676 19612
rect 7612 19552 7676 19556
rect 7692 19612 7756 19616
rect 7692 19556 7696 19612
rect 7696 19556 7752 19612
rect 7752 19556 7756 19612
rect 7692 19552 7756 19556
rect 7772 19612 7836 19616
rect 7772 19556 7776 19612
rect 7776 19556 7832 19612
rect 7832 19556 7836 19612
rect 7772 19552 7836 19556
rect 7852 19612 7916 19616
rect 7852 19556 7856 19612
rect 7856 19556 7912 19612
rect 7912 19556 7916 19612
rect 7852 19552 7916 19556
rect 12612 19612 12676 19616
rect 12612 19556 12616 19612
rect 12616 19556 12672 19612
rect 12672 19556 12676 19612
rect 12612 19552 12676 19556
rect 12692 19612 12756 19616
rect 12692 19556 12696 19612
rect 12696 19556 12752 19612
rect 12752 19556 12756 19612
rect 12692 19552 12756 19556
rect 12772 19612 12836 19616
rect 12772 19556 12776 19612
rect 12776 19556 12832 19612
rect 12832 19556 12836 19612
rect 12772 19552 12836 19556
rect 12852 19612 12916 19616
rect 12852 19556 12856 19612
rect 12856 19556 12912 19612
rect 12912 19556 12916 19612
rect 12852 19552 12916 19556
rect 17612 19612 17676 19616
rect 17612 19556 17616 19612
rect 17616 19556 17672 19612
rect 17672 19556 17676 19612
rect 17612 19552 17676 19556
rect 17692 19612 17756 19616
rect 17692 19556 17696 19612
rect 17696 19556 17752 19612
rect 17752 19556 17756 19612
rect 17692 19552 17756 19556
rect 17772 19612 17836 19616
rect 17772 19556 17776 19612
rect 17776 19556 17832 19612
rect 17832 19556 17836 19612
rect 17772 19552 17836 19556
rect 17852 19612 17916 19616
rect 17852 19556 17856 19612
rect 17856 19556 17912 19612
rect 17912 19556 17916 19612
rect 17852 19552 17916 19556
rect 22612 19612 22676 19616
rect 22612 19556 22616 19612
rect 22616 19556 22672 19612
rect 22672 19556 22676 19612
rect 22612 19552 22676 19556
rect 22692 19612 22756 19616
rect 22692 19556 22696 19612
rect 22696 19556 22752 19612
rect 22752 19556 22756 19612
rect 22692 19552 22756 19556
rect 22772 19612 22836 19616
rect 22772 19556 22776 19612
rect 22776 19556 22832 19612
rect 22832 19556 22836 19612
rect 22772 19552 22836 19556
rect 22852 19612 22916 19616
rect 22852 19556 22856 19612
rect 22856 19556 22912 19612
rect 22912 19556 22916 19612
rect 22852 19552 22916 19556
rect 27612 19612 27676 19616
rect 27612 19556 27616 19612
rect 27616 19556 27672 19612
rect 27672 19556 27676 19612
rect 27612 19552 27676 19556
rect 27692 19612 27756 19616
rect 27692 19556 27696 19612
rect 27696 19556 27752 19612
rect 27752 19556 27756 19612
rect 27692 19552 27756 19556
rect 27772 19612 27836 19616
rect 27772 19556 27776 19612
rect 27776 19556 27832 19612
rect 27832 19556 27836 19612
rect 27772 19552 27836 19556
rect 27852 19612 27916 19616
rect 27852 19556 27856 19612
rect 27856 19556 27912 19612
rect 27912 19556 27916 19612
rect 27852 19552 27916 19556
rect 32612 19612 32676 19616
rect 32612 19556 32616 19612
rect 32616 19556 32672 19612
rect 32672 19556 32676 19612
rect 32612 19552 32676 19556
rect 32692 19612 32756 19616
rect 32692 19556 32696 19612
rect 32696 19556 32752 19612
rect 32752 19556 32756 19612
rect 32692 19552 32756 19556
rect 32772 19612 32836 19616
rect 32772 19556 32776 19612
rect 32776 19556 32832 19612
rect 32832 19556 32836 19612
rect 32772 19552 32836 19556
rect 32852 19612 32916 19616
rect 32852 19556 32856 19612
rect 32856 19556 32912 19612
rect 32912 19556 32916 19612
rect 32852 19552 32916 19556
rect 37612 19612 37676 19616
rect 37612 19556 37616 19612
rect 37616 19556 37672 19612
rect 37672 19556 37676 19612
rect 37612 19552 37676 19556
rect 37692 19612 37756 19616
rect 37692 19556 37696 19612
rect 37696 19556 37752 19612
rect 37752 19556 37756 19612
rect 37692 19552 37756 19556
rect 37772 19612 37836 19616
rect 37772 19556 37776 19612
rect 37776 19556 37832 19612
rect 37832 19556 37836 19612
rect 37772 19552 37836 19556
rect 37852 19612 37916 19616
rect 37852 19556 37856 19612
rect 37856 19556 37912 19612
rect 37912 19556 37916 19612
rect 37852 19552 37916 19556
rect 1952 19068 2016 19072
rect 1952 19012 1956 19068
rect 1956 19012 2012 19068
rect 2012 19012 2016 19068
rect 1952 19008 2016 19012
rect 2032 19068 2096 19072
rect 2032 19012 2036 19068
rect 2036 19012 2092 19068
rect 2092 19012 2096 19068
rect 2032 19008 2096 19012
rect 2112 19068 2176 19072
rect 2112 19012 2116 19068
rect 2116 19012 2172 19068
rect 2172 19012 2176 19068
rect 2112 19008 2176 19012
rect 2192 19068 2256 19072
rect 2192 19012 2196 19068
rect 2196 19012 2252 19068
rect 2252 19012 2256 19068
rect 2192 19008 2256 19012
rect 6952 19068 7016 19072
rect 6952 19012 6956 19068
rect 6956 19012 7012 19068
rect 7012 19012 7016 19068
rect 6952 19008 7016 19012
rect 7032 19068 7096 19072
rect 7032 19012 7036 19068
rect 7036 19012 7092 19068
rect 7092 19012 7096 19068
rect 7032 19008 7096 19012
rect 7112 19068 7176 19072
rect 7112 19012 7116 19068
rect 7116 19012 7172 19068
rect 7172 19012 7176 19068
rect 7112 19008 7176 19012
rect 7192 19068 7256 19072
rect 7192 19012 7196 19068
rect 7196 19012 7252 19068
rect 7252 19012 7256 19068
rect 7192 19008 7256 19012
rect 11952 19068 12016 19072
rect 11952 19012 11956 19068
rect 11956 19012 12012 19068
rect 12012 19012 12016 19068
rect 11952 19008 12016 19012
rect 12032 19068 12096 19072
rect 12032 19012 12036 19068
rect 12036 19012 12092 19068
rect 12092 19012 12096 19068
rect 12032 19008 12096 19012
rect 12112 19068 12176 19072
rect 12112 19012 12116 19068
rect 12116 19012 12172 19068
rect 12172 19012 12176 19068
rect 12112 19008 12176 19012
rect 12192 19068 12256 19072
rect 12192 19012 12196 19068
rect 12196 19012 12252 19068
rect 12252 19012 12256 19068
rect 12192 19008 12256 19012
rect 16952 19068 17016 19072
rect 16952 19012 16956 19068
rect 16956 19012 17012 19068
rect 17012 19012 17016 19068
rect 16952 19008 17016 19012
rect 17032 19068 17096 19072
rect 17032 19012 17036 19068
rect 17036 19012 17092 19068
rect 17092 19012 17096 19068
rect 17032 19008 17096 19012
rect 17112 19068 17176 19072
rect 17112 19012 17116 19068
rect 17116 19012 17172 19068
rect 17172 19012 17176 19068
rect 17112 19008 17176 19012
rect 17192 19068 17256 19072
rect 17192 19012 17196 19068
rect 17196 19012 17252 19068
rect 17252 19012 17256 19068
rect 17192 19008 17256 19012
rect 21952 19068 22016 19072
rect 21952 19012 21956 19068
rect 21956 19012 22012 19068
rect 22012 19012 22016 19068
rect 21952 19008 22016 19012
rect 22032 19068 22096 19072
rect 22032 19012 22036 19068
rect 22036 19012 22092 19068
rect 22092 19012 22096 19068
rect 22032 19008 22096 19012
rect 22112 19068 22176 19072
rect 22112 19012 22116 19068
rect 22116 19012 22172 19068
rect 22172 19012 22176 19068
rect 22112 19008 22176 19012
rect 22192 19068 22256 19072
rect 22192 19012 22196 19068
rect 22196 19012 22252 19068
rect 22252 19012 22256 19068
rect 22192 19008 22256 19012
rect 26952 19068 27016 19072
rect 26952 19012 26956 19068
rect 26956 19012 27012 19068
rect 27012 19012 27016 19068
rect 26952 19008 27016 19012
rect 27032 19068 27096 19072
rect 27032 19012 27036 19068
rect 27036 19012 27092 19068
rect 27092 19012 27096 19068
rect 27032 19008 27096 19012
rect 27112 19068 27176 19072
rect 27112 19012 27116 19068
rect 27116 19012 27172 19068
rect 27172 19012 27176 19068
rect 27112 19008 27176 19012
rect 27192 19068 27256 19072
rect 27192 19012 27196 19068
rect 27196 19012 27252 19068
rect 27252 19012 27256 19068
rect 27192 19008 27256 19012
rect 31952 19068 32016 19072
rect 31952 19012 31956 19068
rect 31956 19012 32012 19068
rect 32012 19012 32016 19068
rect 31952 19008 32016 19012
rect 32032 19068 32096 19072
rect 32032 19012 32036 19068
rect 32036 19012 32092 19068
rect 32092 19012 32096 19068
rect 32032 19008 32096 19012
rect 32112 19068 32176 19072
rect 32112 19012 32116 19068
rect 32116 19012 32172 19068
rect 32172 19012 32176 19068
rect 32112 19008 32176 19012
rect 32192 19068 32256 19072
rect 32192 19012 32196 19068
rect 32196 19012 32252 19068
rect 32252 19012 32256 19068
rect 32192 19008 32256 19012
rect 36952 19068 37016 19072
rect 36952 19012 36956 19068
rect 36956 19012 37012 19068
rect 37012 19012 37016 19068
rect 36952 19008 37016 19012
rect 37032 19068 37096 19072
rect 37032 19012 37036 19068
rect 37036 19012 37092 19068
rect 37092 19012 37096 19068
rect 37032 19008 37096 19012
rect 37112 19068 37176 19072
rect 37112 19012 37116 19068
rect 37116 19012 37172 19068
rect 37172 19012 37176 19068
rect 37112 19008 37176 19012
rect 37192 19068 37256 19072
rect 37192 19012 37196 19068
rect 37196 19012 37252 19068
rect 37252 19012 37256 19068
rect 37192 19008 37256 19012
rect 2612 18524 2676 18528
rect 2612 18468 2616 18524
rect 2616 18468 2672 18524
rect 2672 18468 2676 18524
rect 2612 18464 2676 18468
rect 2692 18524 2756 18528
rect 2692 18468 2696 18524
rect 2696 18468 2752 18524
rect 2752 18468 2756 18524
rect 2692 18464 2756 18468
rect 2772 18524 2836 18528
rect 2772 18468 2776 18524
rect 2776 18468 2832 18524
rect 2832 18468 2836 18524
rect 2772 18464 2836 18468
rect 2852 18524 2916 18528
rect 2852 18468 2856 18524
rect 2856 18468 2912 18524
rect 2912 18468 2916 18524
rect 2852 18464 2916 18468
rect 7612 18524 7676 18528
rect 7612 18468 7616 18524
rect 7616 18468 7672 18524
rect 7672 18468 7676 18524
rect 7612 18464 7676 18468
rect 7692 18524 7756 18528
rect 7692 18468 7696 18524
rect 7696 18468 7752 18524
rect 7752 18468 7756 18524
rect 7692 18464 7756 18468
rect 7772 18524 7836 18528
rect 7772 18468 7776 18524
rect 7776 18468 7832 18524
rect 7832 18468 7836 18524
rect 7772 18464 7836 18468
rect 7852 18524 7916 18528
rect 7852 18468 7856 18524
rect 7856 18468 7912 18524
rect 7912 18468 7916 18524
rect 7852 18464 7916 18468
rect 12612 18524 12676 18528
rect 12612 18468 12616 18524
rect 12616 18468 12672 18524
rect 12672 18468 12676 18524
rect 12612 18464 12676 18468
rect 12692 18524 12756 18528
rect 12692 18468 12696 18524
rect 12696 18468 12752 18524
rect 12752 18468 12756 18524
rect 12692 18464 12756 18468
rect 12772 18524 12836 18528
rect 12772 18468 12776 18524
rect 12776 18468 12832 18524
rect 12832 18468 12836 18524
rect 12772 18464 12836 18468
rect 12852 18524 12916 18528
rect 12852 18468 12856 18524
rect 12856 18468 12912 18524
rect 12912 18468 12916 18524
rect 12852 18464 12916 18468
rect 17612 18524 17676 18528
rect 17612 18468 17616 18524
rect 17616 18468 17672 18524
rect 17672 18468 17676 18524
rect 17612 18464 17676 18468
rect 17692 18524 17756 18528
rect 17692 18468 17696 18524
rect 17696 18468 17752 18524
rect 17752 18468 17756 18524
rect 17692 18464 17756 18468
rect 17772 18524 17836 18528
rect 17772 18468 17776 18524
rect 17776 18468 17832 18524
rect 17832 18468 17836 18524
rect 17772 18464 17836 18468
rect 17852 18524 17916 18528
rect 17852 18468 17856 18524
rect 17856 18468 17912 18524
rect 17912 18468 17916 18524
rect 17852 18464 17916 18468
rect 22612 18524 22676 18528
rect 22612 18468 22616 18524
rect 22616 18468 22672 18524
rect 22672 18468 22676 18524
rect 22612 18464 22676 18468
rect 22692 18524 22756 18528
rect 22692 18468 22696 18524
rect 22696 18468 22752 18524
rect 22752 18468 22756 18524
rect 22692 18464 22756 18468
rect 22772 18524 22836 18528
rect 22772 18468 22776 18524
rect 22776 18468 22832 18524
rect 22832 18468 22836 18524
rect 22772 18464 22836 18468
rect 22852 18524 22916 18528
rect 22852 18468 22856 18524
rect 22856 18468 22912 18524
rect 22912 18468 22916 18524
rect 22852 18464 22916 18468
rect 27612 18524 27676 18528
rect 27612 18468 27616 18524
rect 27616 18468 27672 18524
rect 27672 18468 27676 18524
rect 27612 18464 27676 18468
rect 27692 18524 27756 18528
rect 27692 18468 27696 18524
rect 27696 18468 27752 18524
rect 27752 18468 27756 18524
rect 27692 18464 27756 18468
rect 27772 18524 27836 18528
rect 27772 18468 27776 18524
rect 27776 18468 27832 18524
rect 27832 18468 27836 18524
rect 27772 18464 27836 18468
rect 27852 18524 27916 18528
rect 27852 18468 27856 18524
rect 27856 18468 27912 18524
rect 27912 18468 27916 18524
rect 27852 18464 27916 18468
rect 32612 18524 32676 18528
rect 32612 18468 32616 18524
rect 32616 18468 32672 18524
rect 32672 18468 32676 18524
rect 32612 18464 32676 18468
rect 32692 18524 32756 18528
rect 32692 18468 32696 18524
rect 32696 18468 32752 18524
rect 32752 18468 32756 18524
rect 32692 18464 32756 18468
rect 32772 18524 32836 18528
rect 32772 18468 32776 18524
rect 32776 18468 32832 18524
rect 32832 18468 32836 18524
rect 32772 18464 32836 18468
rect 32852 18524 32916 18528
rect 32852 18468 32856 18524
rect 32856 18468 32912 18524
rect 32912 18468 32916 18524
rect 32852 18464 32916 18468
rect 37612 18524 37676 18528
rect 37612 18468 37616 18524
rect 37616 18468 37672 18524
rect 37672 18468 37676 18524
rect 37612 18464 37676 18468
rect 37692 18524 37756 18528
rect 37692 18468 37696 18524
rect 37696 18468 37752 18524
rect 37752 18468 37756 18524
rect 37692 18464 37756 18468
rect 37772 18524 37836 18528
rect 37772 18468 37776 18524
rect 37776 18468 37832 18524
rect 37832 18468 37836 18524
rect 37772 18464 37836 18468
rect 37852 18524 37916 18528
rect 37852 18468 37856 18524
rect 37856 18468 37912 18524
rect 37912 18468 37916 18524
rect 37852 18464 37916 18468
rect 1952 17980 2016 17984
rect 1952 17924 1956 17980
rect 1956 17924 2012 17980
rect 2012 17924 2016 17980
rect 1952 17920 2016 17924
rect 2032 17980 2096 17984
rect 2032 17924 2036 17980
rect 2036 17924 2092 17980
rect 2092 17924 2096 17980
rect 2032 17920 2096 17924
rect 2112 17980 2176 17984
rect 2112 17924 2116 17980
rect 2116 17924 2172 17980
rect 2172 17924 2176 17980
rect 2112 17920 2176 17924
rect 2192 17980 2256 17984
rect 2192 17924 2196 17980
rect 2196 17924 2252 17980
rect 2252 17924 2256 17980
rect 2192 17920 2256 17924
rect 6952 17980 7016 17984
rect 6952 17924 6956 17980
rect 6956 17924 7012 17980
rect 7012 17924 7016 17980
rect 6952 17920 7016 17924
rect 7032 17980 7096 17984
rect 7032 17924 7036 17980
rect 7036 17924 7092 17980
rect 7092 17924 7096 17980
rect 7032 17920 7096 17924
rect 7112 17980 7176 17984
rect 7112 17924 7116 17980
rect 7116 17924 7172 17980
rect 7172 17924 7176 17980
rect 7112 17920 7176 17924
rect 7192 17980 7256 17984
rect 7192 17924 7196 17980
rect 7196 17924 7252 17980
rect 7252 17924 7256 17980
rect 7192 17920 7256 17924
rect 11952 17980 12016 17984
rect 11952 17924 11956 17980
rect 11956 17924 12012 17980
rect 12012 17924 12016 17980
rect 11952 17920 12016 17924
rect 12032 17980 12096 17984
rect 12032 17924 12036 17980
rect 12036 17924 12092 17980
rect 12092 17924 12096 17980
rect 12032 17920 12096 17924
rect 12112 17980 12176 17984
rect 12112 17924 12116 17980
rect 12116 17924 12172 17980
rect 12172 17924 12176 17980
rect 12112 17920 12176 17924
rect 12192 17980 12256 17984
rect 12192 17924 12196 17980
rect 12196 17924 12252 17980
rect 12252 17924 12256 17980
rect 12192 17920 12256 17924
rect 16952 17980 17016 17984
rect 16952 17924 16956 17980
rect 16956 17924 17012 17980
rect 17012 17924 17016 17980
rect 16952 17920 17016 17924
rect 17032 17980 17096 17984
rect 17032 17924 17036 17980
rect 17036 17924 17092 17980
rect 17092 17924 17096 17980
rect 17032 17920 17096 17924
rect 17112 17980 17176 17984
rect 17112 17924 17116 17980
rect 17116 17924 17172 17980
rect 17172 17924 17176 17980
rect 17112 17920 17176 17924
rect 17192 17980 17256 17984
rect 17192 17924 17196 17980
rect 17196 17924 17252 17980
rect 17252 17924 17256 17980
rect 17192 17920 17256 17924
rect 21952 17980 22016 17984
rect 21952 17924 21956 17980
rect 21956 17924 22012 17980
rect 22012 17924 22016 17980
rect 21952 17920 22016 17924
rect 22032 17980 22096 17984
rect 22032 17924 22036 17980
rect 22036 17924 22092 17980
rect 22092 17924 22096 17980
rect 22032 17920 22096 17924
rect 22112 17980 22176 17984
rect 22112 17924 22116 17980
rect 22116 17924 22172 17980
rect 22172 17924 22176 17980
rect 22112 17920 22176 17924
rect 22192 17980 22256 17984
rect 22192 17924 22196 17980
rect 22196 17924 22252 17980
rect 22252 17924 22256 17980
rect 22192 17920 22256 17924
rect 26952 17980 27016 17984
rect 26952 17924 26956 17980
rect 26956 17924 27012 17980
rect 27012 17924 27016 17980
rect 26952 17920 27016 17924
rect 27032 17980 27096 17984
rect 27032 17924 27036 17980
rect 27036 17924 27092 17980
rect 27092 17924 27096 17980
rect 27032 17920 27096 17924
rect 27112 17980 27176 17984
rect 27112 17924 27116 17980
rect 27116 17924 27172 17980
rect 27172 17924 27176 17980
rect 27112 17920 27176 17924
rect 27192 17980 27256 17984
rect 27192 17924 27196 17980
rect 27196 17924 27252 17980
rect 27252 17924 27256 17980
rect 27192 17920 27256 17924
rect 31952 17980 32016 17984
rect 31952 17924 31956 17980
rect 31956 17924 32012 17980
rect 32012 17924 32016 17980
rect 31952 17920 32016 17924
rect 32032 17980 32096 17984
rect 32032 17924 32036 17980
rect 32036 17924 32092 17980
rect 32092 17924 32096 17980
rect 32032 17920 32096 17924
rect 32112 17980 32176 17984
rect 32112 17924 32116 17980
rect 32116 17924 32172 17980
rect 32172 17924 32176 17980
rect 32112 17920 32176 17924
rect 32192 17980 32256 17984
rect 32192 17924 32196 17980
rect 32196 17924 32252 17980
rect 32252 17924 32256 17980
rect 32192 17920 32256 17924
rect 36952 17980 37016 17984
rect 36952 17924 36956 17980
rect 36956 17924 37012 17980
rect 37012 17924 37016 17980
rect 36952 17920 37016 17924
rect 37032 17980 37096 17984
rect 37032 17924 37036 17980
rect 37036 17924 37092 17980
rect 37092 17924 37096 17980
rect 37032 17920 37096 17924
rect 37112 17980 37176 17984
rect 37112 17924 37116 17980
rect 37116 17924 37172 17980
rect 37172 17924 37176 17980
rect 37112 17920 37176 17924
rect 37192 17980 37256 17984
rect 37192 17924 37196 17980
rect 37196 17924 37252 17980
rect 37252 17924 37256 17980
rect 37192 17920 37256 17924
rect 2612 17436 2676 17440
rect 2612 17380 2616 17436
rect 2616 17380 2672 17436
rect 2672 17380 2676 17436
rect 2612 17376 2676 17380
rect 2692 17436 2756 17440
rect 2692 17380 2696 17436
rect 2696 17380 2752 17436
rect 2752 17380 2756 17436
rect 2692 17376 2756 17380
rect 2772 17436 2836 17440
rect 2772 17380 2776 17436
rect 2776 17380 2832 17436
rect 2832 17380 2836 17436
rect 2772 17376 2836 17380
rect 2852 17436 2916 17440
rect 2852 17380 2856 17436
rect 2856 17380 2912 17436
rect 2912 17380 2916 17436
rect 2852 17376 2916 17380
rect 7612 17436 7676 17440
rect 7612 17380 7616 17436
rect 7616 17380 7672 17436
rect 7672 17380 7676 17436
rect 7612 17376 7676 17380
rect 7692 17436 7756 17440
rect 7692 17380 7696 17436
rect 7696 17380 7752 17436
rect 7752 17380 7756 17436
rect 7692 17376 7756 17380
rect 7772 17436 7836 17440
rect 7772 17380 7776 17436
rect 7776 17380 7832 17436
rect 7832 17380 7836 17436
rect 7772 17376 7836 17380
rect 7852 17436 7916 17440
rect 7852 17380 7856 17436
rect 7856 17380 7912 17436
rect 7912 17380 7916 17436
rect 7852 17376 7916 17380
rect 12612 17436 12676 17440
rect 12612 17380 12616 17436
rect 12616 17380 12672 17436
rect 12672 17380 12676 17436
rect 12612 17376 12676 17380
rect 12692 17436 12756 17440
rect 12692 17380 12696 17436
rect 12696 17380 12752 17436
rect 12752 17380 12756 17436
rect 12692 17376 12756 17380
rect 12772 17436 12836 17440
rect 12772 17380 12776 17436
rect 12776 17380 12832 17436
rect 12832 17380 12836 17436
rect 12772 17376 12836 17380
rect 12852 17436 12916 17440
rect 12852 17380 12856 17436
rect 12856 17380 12912 17436
rect 12912 17380 12916 17436
rect 12852 17376 12916 17380
rect 17612 17436 17676 17440
rect 17612 17380 17616 17436
rect 17616 17380 17672 17436
rect 17672 17380 17676 17436
rect 17612 17376 17676 17380
rect 17692 17436 17756 17440
rect 17692 17380 17696 17436
rect 17696 17380 17752 17436
rect 17752 17380 17756 17436
rect 17692 17376 17756 17380
rect 17772 17436 17836 17440
rect 17772 17380 17776 17436
rect 17776 17380 17832 17436
rect 17832 17380 17836 17436
rect 17772 17376 17836 17380
rect 17852 17436 17916 17440
rect 17852 17380 17856 17436
rect 17856 17380 17912 17436
rect 17912 17380 17916 17436
rect 17852 17376 17916 17380
rect 22612 17436 22676 17440
rect 22612 17380 22616 17436
rect 22616 17380 22672 17436
rect 22672 17380 22676 17436
rect 22612 17376 22676 17380
rect 22692 17436 22756 17440
rect 22692 17380 22696 17436
rect 22696 17380 22752 17436
rect 22752 17380 22756 17436
rect 22692 17376 22756 17380
rect 22772 17436 22836 17440
rect 22772 17380 22776 17436
rect 22776 17380 22832 17436
rect 22832 17380 22836 17436
rect 22772 17376 22836 17380
rect 22852 17436 22916 17440
rect 22852 17380 22856 17436
rect 22856 17380 22912 17436
rect 22912 17380 22916 17436
rect 22852 17376 22916 17380
rect 27612 17436 27676 17440
rect 27612 17380 27616 17436
rect 27616 17380 27672 17436
rect 27672 17380 27676 17436
rect 27612 17376 27676 17380
rect 27692 17436 27756 17440
rect 27692 17380 27696 17436
rect 27696 17380 27752 17436
rect 27752 17380 27756 17436
rect 27692 17376 27756 17380
rect 27772 17436 27836 17440
rect 27772 17380 27776 17436
rect 27776 17380 27832 17436
rect 27832 17380 27836 17436
rect 27772 17376 27836 17380
rect 27852 17436 27916 17440
rect 27852 17380 27856 17436
rect 27856 17380 27912 17436
rect 27912 17380 27916 17436
rect 27852 17376 27916 17380
rect 32612 17436 32676 17440
rect 32612 17380 32616 17436
rect 32616 17380 32672 17436
rect 32672 17380 32676 17436
rect 32612 17376 32676 17380
rect 32692 17436 32756 17440
rect 32692 17380 32696 17436
rect 32696 17380 32752 17436
rect 32752 17380 32756 17436
rect 32692 17376 32756 17380
rect 32772 17436 32836 17440
rect 32772 17380 32776 17436
rect 32776 17380 32832 17436
rect 32832 17380 32836 17436
rect 32772 17376 32836 17380
rect 32852 17436 32916 17440
rect 32852 17380 32856 17436
rect 32856 17380 32912 17436
rect 32912 17380 32916 17436
rect 32852 17376 32916 17380
rect 37612 17436 37676 17440
rect 37612 17380 37616 17436
rect 37616 17380 37672 17436
rect 37672 17380 37676 17436
rect 37612 17376 37676 17380
rect 37692 17436 37756 17440
rect 37692 17380 37696 17436
rect 37696 17380 37752 17436
rect 37752 17380 37756 17436
rect 37692 17376 37756 17380
rect 37772 17436 37836 17440
rect 37772 17380 37776 17436
rect 37776 17380 37832 17436
rect 37832 17380 37836 17436
rect 37772 17376 37836 17380
rect 37852 17436 37916 17440
rect 37852 17380 37856 17436
rect 37856 17380 37912 17436
rect 37912 17380 37916 17436
rect 37852 17376 37916 17380
rect 1952 16892 2016 16896
rect 1952 16836 1956 16892
rect 1956 16836 2012 16892
rect 2012 16836 2016 16892
rect 1952 16832 2016 16836
rect 2032 16892 2096 16896
rect 2032 16836 2036 16892
rect 2036 16836 2092 16892
rect 2092 16836 2096 16892
rect 2032 16832 2096 16836
rect 2112 16892 2176 16896
rect 2112 16836 2116 16892
rect 2116 16836 2172 16892
rect 2172 16836 2176 16892
rect 2112 16832 2176 16836
rect 2192 16892 2256 16896
rect 2192 16836 2196 16892
rect 2196 16836 2252 16892
rect 2252 16836 2256 16892
rect 2192 16832 2256 16836
rect 6952 16892 7016 16896
rect 6952 16836 6956 16892
rect 6956 16836 7012 16892
rect 7012 16836 7016 16892
rect 6952 16832 7016 16836
rect 7032 16892 7096 16896
rect 7032 16836 7036 16892
rect 7036 16836 7092 16892
rect 7092 16836 7096 16892
rect 7032 16832 7096 16836
rect 7112 16892 7176 16896
rect 7112 16836 7116 16892
rect 7116 16836 7172 16892
rect 7172 16836 7176 16892
rect 7112 16832 7176 16836
rect 7192 16892 7256 16896
rect 7192 16836 7196 16892
rect 7196 16836 7252 16892
rect 7252 16836 7256 16892
rect 7192 16832 7256 16836
rect 11952 16892 12016 16896
rect 11952 16836 11956 16892
rect 11956 16836 12012 16892
rect 12012 16836 12016 16892
rect 11952 16832 12016 16836
rect 12032 16892 12096 16896
rect 12032 16836 12036 16892
rect 12036 16836 12092 16892
rect 12092 16836 12096 16892
rect 12032 16832 12096 16836
rect 12112 16892 12176 16896
rect 12112 16836 12116 16892
rect 12116 16836 12172 16892
rect 12172 16836 12176 16892
rect 12112 16832 12176 16836
rect 12192 16892 12256 16896
rect 12192 16836 12196 16892
rect 12196 16836 12252 16892
rect 12252 16836 12256 16892
rect 12192 16832 12256 16836
rect 16952 16892 17016 16896
rect 16952 16836 16956 16892
rect 16956 16836 17012 16892
rect 17012 16836 17016 16892
rect 16952 16832 17016 16836
rect 17032 16892 17096 16896
rect 17032 16836 17036 16892
rect 17036 16836 17092 16892
rect 17092 16836 17096 16892
rect 17032 16832 17096 16836
rect 17112 16892 17176 16896
rect 17112 16836 17116 16892
rect 17116 16836 17172 16892
rect 17172 16836 17176 16892
rect 17112 16832 17176 16836
rect 17192 16892 17256 16896
rect 17192 16836 17196 16892
rect 17196 16836 17252 16892
rect 17252 16836 17256 16892
rect 17192 16832 17256 16836
rect 21952 16892 22016 16896
rect 21952 16836 21956 16892
rect 21956 16836 22012 16892
rect 22012 16836 22016 16892
rect 21952 16832 22016 16836
rect 22032 16892 22096 16896
rect 22032 16836 22036 16892
rect 22036 16836 22092 16892
rect 22092 16836 22096 16892
rect 22032 16832 22096 16836
rect 22112 16892 22176 16896
rect 22112 16836 22116 16892
rect 22116 16836 22172 16892
rect 22172 16836 22176 16892
rect 22112 16832 22176 16836
rect 22192 16892 22256 16896
rect 22192 16836 22196 16892
rect 22196 16836 22252 16892
rect 22252 16836 22256 16892
rect 22192 16832 22256 16836
rect 26952 16892 27016 16896
rect 26952 16836 26956 16892
rect 26956 16836 27012 16892
rect 27012 16836 27016 16892
rect 26952 16832 27016 16836
rect 27032 16892 27096 16896
rect 27032 16836 27036 16892
rect 27036 16836 27092 16892
rect 27092 16836 27096 16892
rect 27032 16832 27096 16836
rect 27112 16892 27176 16896
rect 27112 16836 27116 16892
rect 27116 16836 27172 16892
rect 27172 16836 27176 16892
rect 27112 16832 27176 16836
rect 27192 16892 27256 16896
rect 27192 16836 27196 16892
rect 27196 16836 27252 16892
rect 27252 16836 27256 16892
rect 27192 16832 27256 16836
rect 31952 16892 32016 16896
rect 31952 16836 31956 16892
rect 31956 16836 32012 16892
rect 32012 16836 32016 16892
rect 31952 16832 32016 16836
rect 32032 16892 32096 16896
rect 32032 16836 32036 16892
rect 32036 16836 32092 16892
rect 32092 16836 32096 16892
rect 32032 16832 32096 16836
rect 32112 16892 32176 16896
rect 32112 16836 32116 16892
rect 32116 16836 32172 16892
rect 32172 16836 32176 16892
rect 32112 16832 32176 16836
rect 32192 16892 32256 16896
rect 32192 16836 32196 16892
rect 32196 16836 32252 16892
rect 32252 16836 32256 16892
rect 32192 16832 32256 16836
rect 36952 16892 37016 16896
rect 36952 16836 36956 16892
rect 36956 16836 37012 16892
rect 37012 16836 37016 16892
rect 36952 16832 37016 16836
rect 37032 16892 37096 16896
rect 37032 16836 37036 16892
rect 37036 16836 37092 16892
rect 37092 16836 37096 16892
rect 37032 16832 37096 16836
rect 37112 16892 37176 16896
rect 37112 16836 37116 16892
rect 37116 16836 37172 16892
rect 37172 16836 37176 16892
rect 37112 16832 37176 16836
rect 37192 16892 37256 16896
rect 37192 16836 37196 16892
rect 37196 16836 37252 16892
rect 37252 16836 37256 16892
rect 37192 16832 37256 16836
rect 2612 16348 2676 16352
rect 2612 16292 2616 16348
rect 2616 16292 2672 16348
rect 2672 16292 2676 16348
rect 2612 16288 2676 16292
rect 2692 16348 2756 16352
rect 2692 16292 2696 16348
rect 2696 16292 2752 16348
rect 2752 16292 2756 16348
rect 2692 16288 2756 16292
rect 2772 16348 2836 16352
rect 2772 16292 2776 16348
rect 2776 16292 2832 16348
rect 2832 16292 2836 16348
rect 2772 16288 2836 16292
rect 2852 16348 2916 16352
rect 2852 16292 2856 16348
rect 2856 16292 2912 16348
rect 2912 16292 2916 16348
rect 2852 16288 2916 16292
rect 7612 16348 7676 16352
rect 7612 16292 7616 16348
rect 7616 16292 7672 16348
rect 7672 16292 7676 16348
rect 7612 16288 7676 16292
rect 7692 16348 7756 16352
rect 7692 16292 7696 16348
rect 7696 16292 7752 16348
rect 7752 16292 7756 16348
rect 7692 16288 7756 16292
rect 7772 16348 7836 16352
rect 7772 16292 7776 16348
rect 7776 16292 7832 16348
rect 7832 16292 7836 16348
rect 7772 16288 7836 16292
rect 7852 16348 7916 16352
rect 7852 16292 7856 16348
rect 7856 16292 7912 16348
rect 7912 16292 7916 16348
rect 7852 16288 7916 16292
rect 12612 16348 12676 16352
rect 12612 16292 12616 16348
rect 12616 16292 12672 16348
rect 12672 16292 12676 16348
rect 12612 16288 12676 16292
rect 12692 16348 12756 16352
rect 12692 16292 12696 16348
rect 12696 16292 12752 16348
rect 12752 16292 12756 16348
rect 12692 16288 12756 16292
rect 12772 16348 12836 16352
rect 12772 16292 12776 16348
rect 12776 16292 12832 16348
rect 12832 16292 12836 16348
rect 12772 16288 12836 16292
rect 12852 16348 12916 16352
rect 12852 16292 12856 16348
rect 12856 16292 12912 16348
rect 12912 16292 12916 16348
rect 12852 16288 12916 16292
rect 17612 16348 17676 16352
rect 17612 16292 17616 16348
rect 17616 16292 17672 16348
rect 17672 16292 17676 16348
rect 17612 16288 17676 16292
rect 17692 16348 17756 16352
rect 17692 16292 17696 16348
rect 17696 16292 17752 16348
rect 17752 16292 17756 16348
rect 17692 16288 17756 16292
rect 17772 16348 17836 16352
rect 17772 16292 17776 16348
rect 17776 16292 17832 16348
rect 17832 16292 17836 16348
rect 17772 16288 17836 16292
rect 17852 16348 17916 16352
rect 17852 16292 17856 16348
rect 17856 16292 17912 16348
rect 17912 16292 17916 16348
rect 17852 16288 17916 16292
rect 22612 16348 22676 16352
rect 22612 16292 22616 16348
rect 22616 16292 22672 16348
rect 22672 16292 22676 16348
rect 22612 16288 22676 16292
rect 22692 16348 22756 16352
rect 22692 16292 22696 16348
rect 22696 16292 22752 16348
rect 22752 16292 22756 16348
rect 22692 16288 22756 16292
rect 22772 16348 22836 16352
rect 22772 16292 22776 16348
rect 22776 16292 22832 16348
rect 22832 16292 22836 16348
rect 22772 16288 22836 16292
rect 22852 16348 22916 16352
rect 22852 16292 22856 16348
rect 22856 16292 22912 16348
rect 22912 16292 22916 16348
rect 22852 16288 22916 16292
rect 27612 16348 27676 16352
rect 27612 16292 27616 16348
rect 27616 16292 27672 16348
rect 27672 16292 27676 16348
rect 27612 16288 27676 16292
rect 27692 16348 27756 16352
rect 27692 16292 27696 16348
rect 27696 16292 27752 16348
rect 27752 16292 27756 16348
rect 27692 16288 27756 16292
rect 27772 16348 27836 16352
rect 27772 16292 27776 16348
rect 27776 16292 27832 16348
rect 27832 16292 27836 16348
rect 27772 16288 27836 16292
rect 27852 16348 27916 16352
rect 27852 16292 27856 16348
rect 27856 16292 27912 16348
rect 27912 16292 27916 16348
rect 27852 16288 27916 16292
rect 32612 16348 32676 16352
rect 32612 16292 32616 16348
rect 32616 16292 32672 16348
rect 32672 16292 32676 16348
rect 32612 16288 32676 16292
rect 32692 16348 32756 16352
rect 32692 16292 32696 16348
rect 32696 16292 32752 16348
rect 32752 16292 32756 16348
rect 32692 16288 32756 16292
rect 32772 16348 32836 16352
rect 32772 16292 32776 16348
rect 32776 16292 32832 16348
rect 32832 16292 32836 16348
rect 32772 16288 32836 16292
rect 32852 16348 32916 16352
rect 32852 16292 32856 16348
rect 32856 16292 32912 16348
rect 32912 16292 32916 16348
rect 32852 16288 32916 16292
rect 37612 16348 37676 16352
rect 37612 16292 37616 16348
rect 37616 16292 37672 16348
rect 37672 16292 37676 16348
rect 37612 16288 37676 16292
rect 37692 16348 37756 16352
rect 37692 16292 37696 16348
rect 37696 16292 37752 16348
rect 37752 16292 37756 16348
rect 37692 16288 37756 16292
rect 37772 16348 37836 16352
rect 37772 16292 37776 16348
rect 37776 16292 37832 16348
rect 37832 16292 37836 16348
rect 37772 16288 37836 16292
rect 37852 16348 37916 16352
rect 37852 16292 37856 16348
rect 37856 16292 37912 16348
rect 37912 16292 37916 16348
rect 37852 16288 37916 16292
rect 1952 15804 2016 15808
rect 1952 15748 1956 15804
rect 1956 15748 2012 15804
rect 2012 15748 2016 15804
rect 1952 15744 2016 15748
rect 2032 15804 2096 15808
rect 2032 15748 2036 15804
rect 2036 15748 2092 15804
rect 2092 15748 2096 15804
rect 2032 15744 2096 15748
rect 2112 15804 2176 15808
rect 2112 15748 2116 15804
rect 2116 15748 2172 15804
rect 2172 15748 2176 15804
rect 2112 15744 2176 15748
rect 2192 15804 2256 15808
rect 2192 15748 2196 15804
rect 2196 15748 2252 15804
rect 2252 15748 2256 15804
rect 2192 15744 2256 15748
rect 6952 15804 7016 15808
rect 6952 15748 6956 15804
rect 6956 15748 7012 15804
rect 7012 15748 7016 15804
rect 6952 15744 7016 15748
rect 7032 15804 7096 15808
rect 7032 15748 7036 15804
rect 7036 15748 7092 15804
rect 7092 15748 7096 15804
rect 7032 15744 7096 15748
rect 7112 15804 7176 15808
rect 7112 15748 7116 15804
rect 7116 15748 7172 15804
rect 7172 15748 7176 15804
rect 7112 15744 7176 15748
rect 7192 15804 7256 15808
rect 7192 15748 7196 15804
rect 7196 15748 7252 15804
rect 7252 15748 7256 15804
rect 7192 15744 7256 15748
rect 11952 15804 12016 15808
rect 11952 15748 11956 15804
rect 11956 15748 12012 15804
rect 12012 15748 12016 15804
rect 11952 15744 12016 15748
rect 12032 15804 12096 15808
rect 12032 15748 12036 15804
rect 12036 15748 12092 15804
rect 12092 15748 12096 15804
rect 12032 15744 12096 15748
rect 12112 15804 12176 15808
rect 12112 15748 12116 15804
rect 12116 15748 12172 15804
rect 12172 15748 12176 15804
rect 12112 15744 12176 15748
rect 12192 15804 12256 15808
rect 12192 15748 12196 15804
rect 12196 15748 12252 15804
rect 12252 15748 12256 15804
rect 12192 15744 12256 15748
rect 16952 15804 17016 15808
rect 16952 15748 16956 15804
rect 16956 15748 17012 15804
rect 17012 15748 17016 15804
rect 16952 15744 17016 15748
rect 17032 15804 17096 15808
rect 17032 15748 17036 15804
rect 17036 15748 17092 15804
rect 17092 15748 17096 15804
rect 17032 15744 17096 15748
rect 17112 15804 17176 15808
rect 17112 15748 17116 15804
rect 17116 15748 17172 15804
rect 17172 15748 17176 15804
rect 17112 15744 17176 15748
rect 17192 15804 17256 15808
rect 17192 15748 17196 15804
rect 17196 15748 17252 15804
rect 17252 15748 17256 15804
rect 17192 15744 17256 15748
rect 21952 15804 22016 15808
rect 21952 15748 21956 15804
rect 21956 15748 22012 15804
rect 22012 15748 22016 15804
rect 21952 15744 22016 15748
rect 22032 15804 22096 15808
rect 22032 15748 22036 15804
rect 22036 15748 22092 15804
rect 22092 15748 22096 15804
rect 22032 15744 22096 15748
rect 22112 15804 22176 15808
rect 22112 15748 22116 15804
rect 22116 15748 22172 15804
rect 22172 15748 22176 15804
rect 22112 15744 22176 15748
rect 22192 15804 22256 15808
rect 22192 15748 22196 15804
rect 22196 15748 22252 15804
rect 22252 15748 22256 15804
rect 22192 15744 22256 15748
rect 26952 15804 27016 15808
rect 26952 15748 26956 15804
rect 26956 15748 27012 15804
rect 27012 15748 27016 15804
rect 26952 15744 27016 15748
rect 27032 15804 27096 15808
rect 27032 15748 27036 15804
rect 27036 15748 27092 15804
rect 27092 15748 27096 15804
rect 27032 15744 27096 15748
rect 27112 15804 27176 15808
rect 27112 15748 27116 15804
rect 27116 15748 27172 15804
rect 27172 15748 27176 15804
rect 27112 15744 27176 15748
rect 27192 15804 27256 15808
rect 27192 15748 27196 15804
rect 27196 15748 27252 15804
rect 27252 15748 27256 15804
rect 27192 15744 27256 15748
rect 31952 15804 32016 15808
rect 31952 15748 31956 15804
rect 31956 15748 32012 15804
rect 32012 15748 32016 15804
rect 31952 15744 32016 15748
rect 32032 15804 32096 15808
rect 32032 15748 32036 15804
rect 32036 15748 32092 15804
rect 32092 15748 32096 15804
rect 32032 15744 32096 15748
rect 32112 15804 32176 15808
rect 32112 15748 32116 15804
rect 32116 15748 32172 15804
rect 32172 15748 32176 15804
rect 32112 15744 32176 15748
rect 32192 15804 32256 15808
rect 32192 15748 32196 15804
rect 32196 15748 32252 15804
rect 32252 15748 32256 15804
rect 32192 15744 32256 15748
rect 36952 15804 37016 15808
rect 36952 15748 36956 15804
rect 36956 15748 37012 15804
rect 37012 15748 37016 15804
rect 36952 15744 37016 15748
rect 37032 15804 37096 15808
rect 37032 15748 37036 15804
rect 37036 15748 37092 15804
rect 37092 15748 37096 15804
rect 37032 15744 37096 15748
rect 37112 15804 37176 15808
rect 37112 15748 37116 15804
rect 37116 15748 37172 15804
rect 37172 15748 37176 15804
rect 37112 15744 37176 15748
rect 37192 15804 37256 15808
rect 37192 15748 37196 15804
rect 37196 15748 37252 15804
rect 37252 15748 37256 15804
rect 37192 15744 37256 15748
rect 2612 15260 2676 15264
rect 2612 15204 2616 15260
rect 2616 15204 2672 15260
rect 2672 15204 2676 15260
rect 2612 15200 2676 15204
rect 2692 15260 2756 15264
rect 2692 15204 2696 15260
rect 2696 15204 2752 15260
rect 2752 15204 2756 15260
rect 2692 15200 2756 15204
rect 2772 15260 2836 15264
rect 2772 15204 2776 15260
rect 2776 15204 2832 15260
rect 2832 15204 2836 15260
rect 2772 15200 2836 15204
rect 2852 15260 2916 15264
rect 2852 15204 2856 15260
rect 2856 15204 2912 15260
rect 2912 15204 2916 15260
rect 2852 15200 2916 15204
rect 7612 15260 7676 15264
rect 7612 15204 7616 15260
rect 7616 15204 7672 15260
rect 7672 15204 7676 15260
rect 7612 15200 7676 15204
rect 7692 15260 7756 15264
rect 7692 15204 7696 15260
rect 7696 15204 7752 15260
rect 7752 15204 7756 15260
rect 7692 15200 7756 15204
rect 7772 15260 7836 15264
rect 7772 15204 7776 15260
rect 7776 15204 7832 15260
rect 7832 15204 7836 15260
rect 7772 15200 7836 15204
rect 7852 15260 7916 15264
rect 7852 15204 7856 15260
rect 7856 15204 7912 15260
rect 7912 15204 7916 15260
rect 7852 15200 7916 15204
rect 12612 15260 12676 15264
rect 12612 15204 12616 15260
rect 12616 15204 12672 15260
rect 12672 15204 12676 15260
rect 12612 15200 12676 15204
rect 12692 15260 12756 15264
rect 12692 15204 12696 15260
rect 12696 15204 12752 15260
rect 12752 15204 12756 15260
rect 12692 15200 12756 15204
rect 12772 15260 12836 15264
rect 12772 15204 12776 15260
rect 12776 15204 12832 15260
rect 12832 15204 12836 15260
rect 12772 15200 12836 15204
rect 12852 15260 12916 15264
rect 12852 15204 12856 15260
rect 12856 15204 12912 15260
rect 12912 15204 12916 15260
rect 12852 15200 12916 15204
rect 17612 15260 17676 15264
rect 17612 15204 17616 15260
rect 17616 15204 17672 15260
rect 17672 15204 17676 15260
rect 17612 15200 17676 15204
rect 17692 15260 17756 15264
rect 17692 15204 17696 15260
rect 17696 15204 17752 15260
rect 17752 15204 17756 15260
rect 17692 15200 17756 15204
rect 17772 15260 17836 15264
rect 17772 15204 17776 15260
rect 17776 15204 17832 15260
rect 17832 15204 17836 15260
rect 17772 15200 17836 15204
rect 17852 15260 17916 15264
rect 17852 15204 17856 15260
rect 17856 15204 17912 15260
rect 17912 15204 17916 15260
rect 17852 15200 17916 15204
rect 22612 15260 22676 15264
rect 22612 15204 22616 15260
rect 22616 15204 22672 15260
rect 22672 15204 22676 15260
rect 22612 15200 22676 15204
rect 22692 15260 22756 15264
rect 22692 15204 22696 15260
rect 22696 15204 22752 15260
rect 22752 15204 22756 15260
rect 22692 15200 22756 15204
rect 22772 15260 22836 15264
rect 22772 15204 22776 15260
rect 22776 15204 22832 15260
rect 22832 15204 22836 15260
rect 22772 15200 22836 15204
rect 22852 15260 22916 15264
rect 22852 15204 22856 15260
rect 22856 15204 22912 15260
rect 22912 15204 22916 15260
rect 22852 15200 22916 15204
rect 27612 15260 27676 15264
rect 27612 15204 27616 15260
rect 27616 15204 27672 15260
rect 27672 15204 27676 15260
rect 27612 15200 27676 15204
rect 27692 15260 27756 15264
rect 27692 15204 27696 15260
rect 27696 15204 27752 15260
rect 27752 15204 27756 15260
rect 27692 15200 27756 15204
rect 27772 15260 27836 15264
rect 27772 15204 27776 15260
rect 27776 15204 27832 15260
rect 27832 15204 27836 15260
rect 27772 15200 27836 15204
rect 27852 15260 27916 15264
rect 27852 15204 27856 15260
rect 27856 15204 27912 15260
rect 27912 15204 27916 15260
rect 27852 15200 27916 15204
rect 32612 15260 32676 15264
rect 32612 15204 32616 15260
rect 32616 15204 32672 15260
rect 32672 15204 32676 15260
rect 32612 15200 32676 15204
rect 32692 15260 32756 15264
rect 32692 15204 32696 15260
rect 32696 15204 32752 15260
rect 32752 15204 32756 15260
rect 32692 15200 32756 15204
rect 32772 15260 32836 15264
rect 32772 15204 32776 15260
rect 32776 15204 32832 15260
rect 32832 15204 32836 15260
rect 32772 15200 32836 15204
rect 32852 15260 32916 15264
rect 32852 15204 32856 15260
rect 32856 15204 32912 15260
rect 32912 15204 32916 15260
rect 32852 15200 32916 15204
rect 37612 15260 37676 15264
rect 37612 15204 37616 15260
rect 37616 15204 37672 15260
rect 37672 15204 37676 15260
rect 37612 15200 37676 15204
rect 37692 15260 37756 15264
rect 37692 15204 37696 15260
rect 37696 15204 37752 15260
rect 37752 15204 37756 15260
rect 37692 15200 37756 15204
rect 37772 15260 37836 15264
rect 37772 15204 37776 15260
rect 37776 15204 37832 15260
rect 37832 15204 37836 15260
rect 37772 15200 37836 15204
rect 37852 15260 37916 15264
rect 37852 15204 37856 15260
rect 37856 15204 37912 15260
rect 37912 15204 37916 15260
rect 37852 15200 37916 15204
rect 1952 14716 2016 14720
rect 1952 14660 1956 14716
rect 1956 14660 2012 14716
rect 2012 14660 2016 14716
rect 1952 14656 2016 14660
rect 2032 14716 2096 14720
rect 2032 14660 2036 14716
rect 2036 14660 2092 14716
rect 2092 14660 2096 14716
rect 2032 14656 2096 14660
rect 2112 14716 2176 14720
rect 2112 14660 2116 14716
rect 2116 14660 2172 14716
rect 2172 14660 2176 14716
rect 2112 14656 2176 14660
rect 2192 14716 2256 14720
rect 2192 14660 2196 14716
rect 2196 14660 2252 14716
rect 2252 14660 2256 14716
rect 2192 14656 2256 14660
rect 6952 14716 7016 14720
rect 6952 14660 6956 14716
rect 6956 14660 7012 14716
rect 7012 14660 7016 14716
rect 6952 14656 7016 14660
rect 7032 14716 7096 14720
rect 7032 14660 7036 14716
rect 7036 14660 7092 14716
rect 7092 14660 7096 14716
rect 7032 14656 7096 14660
rect 7112 14716 7176 14720
rect 7112 14660 7116 14716
rect 7116 14660 7172 14716
rect 7172 14660 7176 14716
rect 7112 14656 7176 14660
rect 7192 14716 7256 14720
rect 7192 14660 7196 14716
rect 7196 14660 7252 14716
rect 7252 14660 7256 14716
rect 7192 14656 7256 14660
rect 11952 14716 12016 14720
rect 11952 14660 11956 14716
rect 11956 14660 12012 14716
rect 12012 14660 12016 14716
rect 11952 14656 12016 14660
rect 12032 14716 12096 14720
rect 12032 14660 12036 14716
rect 12036 14660 12092 14716
rect 12092 14660 12096 14716
rect 12032 14656 12096 14660
rect 12112 14716 12176 14720
rect 12112 14660 12116 14716
rect 12116 14660 12172 14716
rect 12172 14660 12176 14716
rect 12112 14656 12176 14660
rect 12192 14716 12256 14720
rect 12192 14660 12196 14716
rect 12196 14660 12252 14716
rect 12252 14660 12256 14716
rect 12192 14656 12256 14660
rect 16952 14716 17016 14720
rect 16952 14660 16956 14716
rect 16956 14660 17012 14716
rect 17012 14660 17016 14716
rect 16952 14656 17016 14660
rect 17032 14716 17096 14720
rect 17032 14660 17036 14716
rect 17036 14660 17092 14716
rect 17092 14660 17096 14716
rect 17032 14656 17096 14660
rect 17112 14716 17176 14720
rect 17112 14660 17116 14716
rect 17116 14660 17172 14716
rect 17172 14660 17176 14716
rect 17112 14656 17176 14660
rect 17192 14716 17256 14720
rect 17192 14660 17196 14716
rect 17196 14660 17252 14716
rect 17252 14660 17256 14716
rect 17192 14656 17256 14660
rect 21952 14716 22016 14720
rect 21952 14660 21956 14716
rect 21956 14660 22012 14716
rect 22012 14660 22016 14716
rect 21952 14656 22016 14660
rect 22032 14716 22096 14720
rect 22032 14660 22036 14716
rect 22036 14660 22092 14716
rect 22092 14660 22096 14716
rect 22032 14656 22096 14660
rect 22112 14716 22176 14720
rect 22112 14660 22116 14716
rect 22116 14660 22172 14716
rect 22172 14660 22176 14716
rect 22112 14656 22176 14660
rect 22192 14716 22256 14720
rect 22192 14660 22196 14716
rect 22196 14660 22252 14716
rect 22252 14660 22256 14716
rect 22192 14656 22256 14660
rect 26952 14716 27016 14720
rect 26952 14660 26956 14716
rect 26956 14660 27012 14716
rect 27012 14660 27016 14716
rect 26952 14656 27016 14660
rect 27032 14716 27096 14720
rect 27032 14660 27036 14716
rect 27036 14660 27092 14716
rect 27092 14660 27096 14716
rect 27032 14656 27096 14660
rect 27112 14716 27176 14720
rect 27112 14660 27116 14716
rect 27116 14660 27172 14716
rect 27172 14660 27176 14716
rect 27112 14656 27176 14660
rect 27192 14716 27256 14720
rect 27192 14660 27196 14716
rect 27196 14660 27252 14716
rect 27252 14660 27256 14716
rect 27192 14656 27256 14660
rect 31952 14716 32016 14720
rect 31952 14660 31956 14716
rect 31956 14660 32012 14716
rect 32012 14660 32016 14716
rect 31952 14656 32016 14660
rect 32032 14716 32096 14720
rect 32032 14660 32036 14716
rect 32036 14660 32092 14716
rect 32092 14660 32096 14716
rect 32032 14656 32096 14660
rect 32112 14716 32176 14720
rect 32112 14660 32116 14716
rect 32116 14660 32172 14716
rect 32172 14660 32176 14716
rect 32112 14656 32176 14660
rect 32192 14716 32256 14720
rect 32192 14660 32196 14716
rect 32196 14660 32252 14716
rect 32252 14660 32256 14716
rect 32192 14656 32256 14660
rect 36952 14716 37016 14720
rect 36952 14660 36956 14716
rect 36956 14660 37012 14716
rect 37012 14660 37016 14716
rect 36952 14656 37016 14660
rect 37032 14716 37096 14720
rect 37032 14660 37036 14716
rect 37036 14660 37092 14716
rect 37092 14660 37096 14716
rect 37032 14656 37096 14660
rect 37112 14716 37176 14720
rect 37112 14660 37116 14716
rect 37116 14660 37172 14716
rect 37172 14660 37176 14716
rect 37112 14656 37176 14660
rect 37192 14716 37256 14720
rect 37192 14660 37196 14716
rect 37196 14660 37252 14716
rect 37252 14660 37256 14716
rect 37192 14656 37256 14660
rect 33916 14316 33980 14380
rect 2612 14172 2676 14176
rect 2612 14116 2616 14172
rect 2616 14116 2672 14172
rect 2672 14116 2676 14172
rect 2612 14112 2676 14116
rect 2692 14172 2756 14176
rect 2692 14116 2696 14172
rect 2696 14116 2752 14172
rect 2752 14116 2756 14172
rect 2692 14112 2756 14116
rect 2772 14172 2836 14176
rect 2772 14116 2776 14172
rect 2776 14116 2832 14172
rect 2832 14116 2836 14172
rect 2772 14112 2836 14116
rect 2852 14172 2916 14176
rect 2852 14116 2856 14172
rect 2856 14116 2912 14172
rect 2912 14116 2916 14172
rect 2852 14112 2916 14116
rect 7612 14172 7676 14176
rect 7612 14116 7616 14172
rect 7616 14116 7672 14172
rect 7672 14116 7676 14172
rect 7612 14112 7676 14116
rect 7692 14172 7756 14176
rect 7692 14116 7696 14172
rect 7696 14116 7752 14172
rect 7752 14116 7756 14172
rect 7692 14112 7756 14116
rect 7772 14172 7836 14176
rect 7772 14116 7776 14172
rect 7776 14116 7832 14172
rect 7832 14116 7836 14172
rect 7772 14112 7836 14116
rect 7852 14172 7916 14176
rect 7852 14116 7856 14172
rect 7856 14116 7912 14172
rect 7912 14116 7916 14172
rect 7852 14112 7916 14116
rect 12612 14172 12676 14176
rect 12612 14116 12616 14172
rect 12616 14116 12672 14172
rect 12672 14116 12676 14172
rect 12612 14112 12676 14116
rect 12692 14172 12756 14176
rect 12692 14116 12696 14172
rect 12696 14116 12752 14172
rect 12752 14116 12756 14172
rect 12692 14112 12756 14116
rect 12772 14172 12836 14176
rect 12772 14116 12776 14172
rect 12776 14116 12832 14172
rect 12832 14116 12836 14172
rect 12772 14112 12836 14116
rect 12852 14172 12916 14176
rect 12852 14116 12856 14172
rect 12856 14116 12912 14172
rect 12912 14116 12916 14172
rect 12852 14112 12916 14116
rect 17612 14172 17676 14176
rect 17612 14116 17616 14172
rect 17616 14116 17672 14172
rect 17672 14116 17676 14172
rect 17612 14112 17676 14116
rect 17692 14172 17756 14176
rect 17692 14116 17696 14172
rect 17696 14116 17752 14172
rect 17752 14116 17756 14172
rect 17692 14112 17756 14116
rect 17772 14172 17836 14176
rect 17772 14116 17776 14172
rect 17776 14116 17832 14172
rect 17832 14116 17836 14172
rect 17772 14112 17836 14116
rect 17852 14172 17916 14176
rect 17852 14116 17856 14172
rect 17856 14116 17912 14172
rect 17912 14116 17916 14172
rect 17852 14112 17916 14116
rect 22612 14172 22676 14176
rect 22612 14116 22616 14172
rect 22616 14116 22672 14172
rect 22672 14116 22676 14172
rect 22612 14112 22676 14116
rect 22692 14172 22756 14176
rect 22692 14116 22696 14172
rect 22696 14116 22752 14172
rect 22752 14116 22756 14172
rect 22692 14112 22756 14116
rect 22772 14172 22836 14176
rect 22772 14116 22776 14172
rect 22776 14116 22832 14172
rect 22832 14116 22836 14172
rect 22772 14112 22836 14116
rect 22852 14172 22916 14176
rect 22852 14116 22856 14172
rect 22856 14116 22912 14172
rect 22912 14116 22916 14172
rect 22852 14112 22916 14116
rect 27612 14172 27676 14176
rect 27612 14116 27616 14172
rect 27616 14116 27672 14172
rect 27672 14116 27676 14172
rect 27612 14112 27676 14116
rect 27692 14172 27756 14176
rect 27692 14116 27696 14172
rect 27696 14116 27752 14172
rect 27752 14116 27756 14172
rect 27692 14112 27756 14116
rect 27772 14172 27836 14176
rect 27772 14116 27776 14172
rect 27776 14116 27832 14172
rect 27832 14116 27836 14172
rect 27772 14112 27836 14116
rect 27852 14172 27916 14176
rect 27852 14116 27856 14172
rect 27856 14116 27912 14172
rect 27912 14116 27916 14172
rect 27852 14112 27916 14116
rect 32612 14172 32676 14176
rect 32612 14116 32616 14172
rect 32616 14116 32672 14172
rect 32672 14116 32676 14172
rect 32612 14112 32676 14116
rect 32692 14172 32756 14176
rect 32692 14116 32696 14172
rect 32696 14116 32752 14172
rect 32752 14116 32756 14172
rect 32692 14112 32756 14116
rect 32772 14172 32836 14176
rect 32772 14116 32776 14172
rect 32776 14116 32832 14172
rect 32832 14116 32836 14172
rect 32772 14112 32836 14116
rect 32852 14172 32916 14176
rect 32852 14116 32856 14172
rect 32856 14116 32912 14172
rect 32912 14116 32916 14172
rect 32852 14112 32916 14116
rect 37612 14172 37676 14176
rect 37612 14116 37616 14172
rect 37616 14116 37672 14172
rect 37672 14116 37676 14172
rect 37612 14112 37676 14116
rect 37692 14172 37756 14176
rect 37692 14116 37696 14172
rect 37696 14116 37752 14172
rect 37752 14116 37756 14172
rect 37692 14112 37756 14116
rect 37772 14172 37836 14176
rect 37772 14116 37776 14172
rect 37776 14116 37832 14172
rect 37832 14116 37836 14172
rect 37772 14112 37836 14116
rect 37852 14172 37916 14176
rect 37852 14116 37856 14172
rect 37856 14116 37912 14172
rect 37912 14116 37916 14172
rect 37852 14112 37916 14116
rect 1952 13628 2016 13632
rect 1952 13572 1956 13628
rect 1956 13572 2012 13628
rect 2012 13572 2016 13628
rect 1952 13568 2016 13572
rect 2032 13628 2096 13632
rect 2032 13572 2036 13628
rect 2036 13572 2092 13628
rect 2092 13572 2096 13628
rect 2032 13568 2096 13572
rect 2112 13628 2176 13632
rect 2112 13572 2116 13628
rect 2116 13572 2172 13628
rect 2172 13572 2176 13628
rect 2112 13568 2176 13572
rect 2192 13628 2256 13632
rect 2192 13572 2196 13628
rect 2196 13572 2252 13628
rect 2252 13572 2256 13628
rect 2192 13568 2256 13572
rect 6952 13628 7016 13632
rect 6952 13572 6956 13628
rect 6956 13572 7012 13628
rect 7012 13572 7016 13628
rect 6952 13568 7016 13572
rect 7032 13628 7096 13632
rect 7032 13572 7036 13628
rect 7036 13572 7092 13628
rect 7092 13572 7096 13628
rect 7032 13568 7096 13572
rect 7112 13628 7176 13632
rect 7112 13572 7116 13628
rect 7116 13572 7172 13628
rect 7172 13572 7176 13628
rect 7112 13568 7176 13572
rect 7192 13628 7256 13632
rect 7192 13572 7196 13628
rect 7196 13572 7252 13628
rect 7252 13572 7256 13628
rect 7192 13568 7256 13572
rect 11952 13628 12016 13632
rect 11952 13572 11956 13628
rect 11956 13572 12012 13628
rect 12012 13572 12016 13628
rect 11952 13568 12016 13572
rect 12032 13628 12096 13632
rect 12032 13572 12036 13628
rect 12036 13572 12092 13628
rect 12092 13572 12096 13628
rect 12032 13568 12096 13572
rect 12112 13628 12176 13632
rect 12112 13572 12116 13628
rect 12116 13572 12172 13628
rect 12172 13572 12176 13628
rect 12112 13568 12176 13572
rect 12192 13628 12256 13632
rect 12192 13572 12196 13628
rect 12196 13572 12252 13628
rect 12252 13572 12256 13628
rect 12192 13568 12256 13572
rect 16952 13628 17016 13632
rect 16952 13572 16956 13628
rect 16956 13572 17012 13628
rect 17012 13572 17016 13628
rect 16952 13568 17016 13572
rect 17032 13628 17096 13632
rect 17032 13572 17036 13628
rect 17036 13572 17092 13628
rect 17092 13572 17096 13628
rect 17032 13568 17096 13572
rect 17112 13628 17176 13632
rect 17112 13572 17116 13628
rect 17116 13572 17172 13628
rect 17172 13572 17176 13628
rect 17112 13568 17176 13572
rect 17192 13628 17256 13632
rect 17192 13572 17196 13628
rect 17196 13572 17252 13628
rect 17252 13572 17256 13628
rect 17192 13568 17256 13572
rect 21952 13628 22016 13632
rect 21952 13572 21956 13628
rect 21956 13572 22012 13628
rect 22012 13572 22016 13628
rect 21952 13568 22016 13572
rect 22032 13628 22096 13632
rect 22032 13572 22036 13628
rect 22036 13572 22092 13628
rect 22092 13572 22096 13628
rect 22032 13568 22096 13572
rect 22112 13628 22176 13632
rect 22112 13572 22116 13628
rect 22116 13572 22172 13628
rect 22172 13572 22176 13628
rect 22112 13568 22176 13572
rect 22192 13628 22256 13632
rect 22192 13572 22196 13628
rect 22196 13572 22252 13628
rect 22252 13572 22256 13628
rect 22192 13568 22256 13572
rect 26952 13628 27016 13632
rect 26952 13572 26956 13628
rect 26956 13572 27012 13628
rect 27012 13572 27016 13628
rect 26952 13568 27016 13572
rect 27032 13628 27096 13632
rect 27032 13572 27036 13628
rect 27036 13572 27092 13628
rect 27092 13572 27096 13628
rect 27032 13568 27096 13572
rect 27112 13628 27176 13632
rect 27112 13572 27116 13628
rect 27116 13572 27172 13628
rect 27172 13572 27176 13628
rect 27112 13568 27176 13572
rect 27192 13628 27256 13632
rect 27192 13572 27196 13628
rect 27196 13572 27252 13628
rect 27252 13572 27256 13628
rect 27192 13568 27256 13572
rect 31952 13628 32016 13632
rect 31952 13572 31956 13628
rect 31956 13572 32012 13628
rect 32012 13572 32016 13628
rect 31952 13568 32016 13572
rect 32032 13628 32096 13632
rect 32032 13572 32036 13628
rect 32036 13572 32092 13628
rect 32092 13572 32096 13628
rect 32032 13568 32096 13572
rect 32112 13628 32176 13632
rect 32112 13572 32116 13628
rect 32116 13572 32172 13628
rect 32172 13572 32176 13628
rect 32112 13568 32176 13572
rect 32192 13628 32256 13632
rect 32192 13572 32196 13628
rect 32196 13572 32252 13628
rect 32252 13572 32256 13628
rect 32192 13568 32256 13572
rect 36952 13628 37016 13632
rect 36952 13572 36956 13628
rect 36956 13572 37012 13628
rect 37012 13572 37016 13628
rect 36952 13568 37016 13572
rect 37032 13628 37096 13632
rect 37032 13572 37036 13628
rect 37036 13572 37092 13628
rect 37092 13572 37096 13628
rect 37032 13568 37096 13572
rect 37112 13628 37176 13632
rect 37112 13572 37116 13628
rect 37116 13572 37172 13628
rect 37172 13572 37176 13628
rect 37112 13568 37176 13572
rect 37192 13628 37256 13632
rect 37192 13572 37196 13628
rect 37196 13572 37252 13628
rect 37252 13572 37256 13628
rect 37192 13568 37256 13572
rect 2612 13084 2676 13088
rect 2612 13028 2616 13084
rect 2616 13028 2672 13084
rect 2672 13028 2676 13084
rect 2612 13024 2676 13028
rect 2692 13084 2756 13088
rect 2692 13028 2696 13084
rect 2696 13028 2752 13084
rect 2752 13028 2756 13084
rect 2692 13024 2756 13028
rect 2772 13084 2836 13088
rect 2772 13028 2776 13084
rect 2776 13028 2832 13084
rect 2832 13028 2836 13084
rect 2772 13024 2836 13028
rect 2852 13084 2916 13088
rect 2852 13028 2856 13084
rect 2856 13028 2912 13084
rect 2912 13028 2916 13084
rect 2852 13024 2916 13028
rect 7612 13084 7676 13088
rect 7612 13028 7616 13084
rect 7616 13028 7672 13084
rect 7672 13028 7676 13084
rect 7612 13024 7676 13028
rect 7692 13084 7756 13088
rect 7692 13028 7696 13084
rect 7696 13028 7752 13084
rect 7752 13028 7756 13084
rect 7692 13024 7756 13028
rect 7772 13084 7836 13088
rect 7772 13028 7776 13084
rect 7776 13028 7832 13084
rect 7832 13028 7836 13084
rect 7772 13024 7836 13028
rect 7852 13084 7916 13088
rect 7852 13028 7856 13084
rect 7856 13028 7912 13084
rect 7912 13028 7916 13084
rect 7852 13024 7916 13028
rect 12612 13084 12676 13088
rect 12612 13028 12616 13084
rect 12616 13028 12672 13084
rect 12672 13028 12676 13084
rect 12612 13024 12676 13028
rect 12692 13084 12756 13088
rect 12692 13028 12696 13084
rect 12696 13028 12752 13084
rect 12752 13028 12756 13084
rect 12692 13024 12756 13028
rect 12772 13084 12836 13088
rect 12772 13028 12776 13084
rect 12776 13028 12832 13084
rect 12832 13028 12836 13084
rect 12772 13024 12836 13028
rect 12852 13084 12916 13088
rect 12852 13028 12856 13084
rect 12856 13028 12912 13084
rect 12912 13028 12916 13084
rect 12852 13024 12916 13028
rect 17612 13084 17676 13088
rect 17612 13028 17616 13084
rect 17616 13028 17672 13084
rect 17672 13028 17676 13084
rect 17612 13024 17676 13028
rect 17692 13084 17756 13088
rect 17692 13028 17696 13084
rect 17696 13028 17752 13084
rect 17752 13028 17756 13084
rect 17692 13024 17756 13028
rect 17772 13084 17836 13088
rect 17772 13028 17776 13084
rect 17776 13028 17832 13084
rect 17832 13028 17836 13084
rect 17772 13024 17836 13028
rect 17852 13084 17916 13088
rect 17852 13028 17856 13084
rect 17856 13028 17912 13084
rect 17912 13028 17916 13084
rect 17852 13024 17916 13028
rect 22612 13084 22676 13088
rect 22612 13028 22616 13084
rect 22616 13028 22672 13084
rect 22672 13028 22676 13084
rect 22612 13024 22676 13028
rect 22692 13084 22756 13088
rect 22692 13028 22696 13084
rect 22696 13028 22752 13084
rect 22752 13028 22756 13084
rect 22692 13024 22756 13028
rect 22772 13084 22836 13088
rect 22772 13028 22776 13084
rect 22776 13028 22832 13084
rect 22832 13028 22836 13084
rect 22772 13024 22836 13028
rect 22852 13084 22916 13088
rect 22852 13028 22856 13084
rect 22856 13028 22912 13084
rect 22912 13028 22916 13084
rect 22852 13024 22916 13028
rect 27612 13084 27676 13088
rect 27612 13028 27616 13084
rect 27616 13028 27672 13084
rect 27672 13028 27676 13084
rect 27612 13024 27676 13028
rect 27692 13084 27756 13088
rect 27692 13028 27696 13084
rect 27696 13028 27752 13084
rect 27752 13028 27756 13084
rect 27692 13024 27756 13028
rect 27772 13084 27836 13088
rect 27772 13028 27776 13084
rect 27776 13028 27832 13084
rect 27832 13028 27836 13084
rect 27772 13024 27836 13028
rect 27852 13084 27916 13088
rect 27852 13028 27856 13084
rect 27856 13028 27912 13084
rect 27912 13028 27916 13084
rect 27852 13024 27916 13028
rect 32612 13084 32676 13088
rect 32612 13028 32616 13084
rect 32616 13028 32672 13084
rect 32672 13028 32676 13084
rect 32612 13024 32676 13028
rect 32692 13084 32756 13088
rect 32692 13028 32696 13084
rect 32696 13028 32752 13084
rect 32752 13028 32756 13084
rect 32692 13024 32756 13028
rect 32772 13084 32836 13088
rect 32772 13028 32776 13084
rect 32776 13028 32832 13084
rect 32832 13028 32836 13084
rect 32772 13024 32836 13028
rect 32852 13084 32916 13088
rect 32852 13028 32856 13084
rect 32856 13028 32912 13084
rect 32912 13028 32916 13084
rect 32852 13024 32916 13028
rect 37612 13084 37676 13088
rect 37612 13028 37616 13084
rect 37616 13028 37672 13084
rect 37672 13028 37676 13084
rect 37612 13024 37676 13028
rect 37692 13084 37756 13088
rect 37692 13028 37696 13084
rect 37696 13028 37752 13084
rect 37752 13028 37756 13084
rect 37692 13024 37756 13028
rect 37772 13084 37836 13088
rect 37772 13028 37776 13084
rect 37776 13028 37832 13084
rect 37832 13028 37836 13084
rect 37772 13024 37836 13028
rect 37852 13084 37916 13088
rect 37852 13028 37856 13084
rect 37856 13028 37912 13084
rect 37912 13028 37916 13084
rect 37852 13024 37916 13028
rect 1952 12540 2016 12544
rect 1952 12484 1956 12540
rect 1956 12484 2012 12540
rect 2012 12484 2016 12540
rect 1952 12480 2016 12484
rect 2032 12540 2096 12544
rect 2032 12484 2036 12540
rect 2036 12484 2092 12540
rect 2092 12484 2096 12540
rect 2032 12480 2096 12484
rect 2112 12540 2176 12544
rect 2112 12484 2116 12540
rect 2116 12484 2172 12540
rect 2172 12484 2176 12540
rect 2112 12480 2176 12484
rect 2192 12540 2256 12544
rect 2192 12484 2196 12540
rect 2196 12484 2252 12540
rect 2252 12484 2256 12540
rect 2192 12480 2256 12484
rect 6952 12540 7016 12544
rect 6952 12484 6956 12540
rect 6956 12484 7012 12540
rect 7012 12484 7016 12540
rect 6952 12480 7016 12484
rect 7032 12540 7096 12544
rect 7032 12484 7036 12540
rect 7036 12484 7092 12540
rect 7092 12484 7096 12540
rect 7032 12480 7096 12484
rect 7112 12540 7176 12544
rect 7112 12484 7116 12540
rect 7116 12484 7172 12540
rect 7172 12484 7176 12540
rect 7112 12480 7176 12484
rect 7192 12540 7256 12544
rect 7192 12484 7196 12540
rect 7196 12484 7252 12540
rect 7252 12484 7256 12540
rect 7192 12480 7256 12484
rect 11952 12540 12016 12544
rect 11952 12484 11956 12540
rect 11956 12484 12012 12540
rect 12012 12484 12016 12540
rect 11952 12480 12016 12484
rect 12032 12540 12096 12544
rect 12032 12484 12036 12540
rect 12036 12484 12092 12540
rect 12092 12484 12096 12540
rect 12032 12480 12096 12484
rect 12112 12540 12176 12544
rect 12112 12484 12116 12540
rect 12116 12484 12172 12540
rect 12172 12484 12176 12540
rect 12112 12480 12176 12484
rect 12192 12540 12256 12544
rect 12192 12484 12196 12540
rect 12196 12484 12252 12540
rect 12252 12484 12256 12540
rect 12192 12480 12256 12484
rect 16952 12540 17016 12544
rect 16952 12484 16956 12540
rect 16956 12484 17012 12540
rect 17012 12484 17016 12540
rect 16952 12480 17016 12484
rect 17032 12540 17096 12544
rect 17032 12484 17036 12540
rect 17036 12484 17092 12540
rect 17092 12484 17096 12540
rect 17032 12480 17096 12484
rect 17112 12540 17176 12544
rect 17112 12484 17116 12540
rect 17116 12484 17172 12540
rect 17172 12484 17176 12540
rect 17112 12480 17176 12484
rect 17192 12540 17256 12544
rect 17192 12484 17196 12540
rect 17196 12484 17252 12540
rect 17252 12484 17256 12540
rect 17192 12480 17256 12484
rect 21952 12540 22016 12544
rect 21952 12484 21956 12540
rect 21956 12484 22012 12540
rect 22012 12484 22016 12540
rect 21952 12480 22016 12484
rect 22032 12540 22096 12544
rect 22032 12484 22036 12540
rect 22036 12484 22092 12540
rect 22092 12484 22096 12540
rect 22032 12480 22096 12484
rect 22112 12540 22176 12544
rect 22112 12484 22116 12540
rect 22116 12484 22172 12540
rect 22172 12484 22176 12540
rect 22112 12480 22176 12484
rect 22192 12540 22256 12544
rect 22192 12484 22196 12540
rect 22196 12484 22252 12540
rect 22252 12484 22256 12540
rect 22192 12480 22256 12484
rect 26952 12540 27016 12544
rect 26952 12484 26956 12540
rect 26956 12484 27012 12540
rect 27012 12484 27016 12540
rect 26952 12480 27016 12484
rect 27032 12540 27096 12544
rect 27032 12484 27036 12540
rect 27036 12484 27092 12540
rect 27092 12484 27096 12540
rect 27032 12480 27096 12484
rect 27112 12540 27176 12544
rect 27112 12484 27116 12540
rect 27116 12484 27172 12540
rect 27172 12484 27176 12540
rect 27112 12480 27176 12484
rect 27192 12540 27256 12544
rect 27192 12484 27196 12540
rect 27196 12484 27252 12540
rect 27252 12484 27256 12540
rect 27192 12480 27256 12484
rect 31952 12540 32016 12544
rect 31952 12484 31956 12540
rect 31956 12484 32012 12540
rect 32012 12484 32016 12540
rect 31952 12480 32016 12484
rect 32032 12540 32096 12544
rect 32032 12484 32036 12540
rect 32036 12484 32092 12540
rect 32092 12484 32096 12540
rect 32032 12480 32096 12484
rect 32112 12540 32176 12544
rect 32112 12484 32116 12540
rect 32116 12484 32172 12540
rect 32172 12484 32176 12540
rect 32112 12480 32176 12484
rect 32192 12540 32256 12544
rect 32192 12484 32196 12540
rect 32196 12484 32252 12540
rect 32252 12484 32256 12540
rect 32192 12480 32256 12484
rect 36952 12540 37016 12544
rect 36952 12484 36956 12540
rect 36956 12484 37012 12540
rect 37012 12484 37016 12540
rect 36952 12480 37016 12484
rect 37032 12540 37096 12544
rect 37032 12484 37036 12540
rect 37036 12484 37092 12540
rect 37092 12484 37096 12540
rect 37032 12480 37096 12484
rect 37112 12540 37176 12544
rect 37112 12484 37116 12540
rect 37116 12484 37172 12540
rect 37172 12484 37176 12540
rect 37112 12480 37176 12484
rect 37192 12540 37256 12544
rect 37192 12484 37196 12540
rect 37196 12484 37252 12540
rect 37252 12484 37256 12540
rect 37192 12480 37256 12484
rect 2612 11996 2676 12000
rect 2612 11940 2616 11996
rect 2616 11940 2672 11996
rect 2672 11940 2676 11996
rect 2612 11936 2676 11940
rect 2692 11996 2756 12000
rect 2692 11940 2696 11996
rect 2696 11940 2752 11996
rect 2752 11940 2756 11996
rect 2692 11936 2756 11940
rect 2772 11996 2836 12000
rect 2772 11940 2776 11996
rect 2776 11940 2832 11996
rect 2832 11940 2836 11996
rect 2772 11936 2836 11940
rect 2852 11996 2916 12000
rect 2852 11940 2856 11996
rect 2856 11940 2912 11996
rect 2912 11940 2916 11996
rect 2852 11936 2916 11940
rect 7612 11996 7676 12000
rect 7612 11940 7616 11996
rect 7616 11940 7672 11996
rect 7672 11940 7676 11996
rect 7612 11936 7676 11940
rect 7692 11996 7756 12000
rect 7692 11940 7696 11996
rect 7696 11940 7752 11996
rect 7752 11940 7756 11996
rect 7692 11936 7756 11940
rect 7772 11996 7836 12000
rect 7772 11940 7776 11996
rect 7776 11940 7832 11996
rect 7832 11940 7836 11996
rect 7772 11936 7836 11940
rect 7852 11996 7916 12000
rect 7852 11940 7856 11996
rect 7856 11940 7912 11996
rect 7912 11940 7916 11996
rect 7852 11936 7916 11940
rect 12612 11996 12676 12000
rect 12612 11940 12616 11996
rect 12616 11940 12672 11996
rect 12672 11940 12676 11996
rect 12612 11936 12676 11940
rect 12692 11996 12756 12000
rect 12692 11940 12696 11996
rect 12696 11940 12752 11996
rect 12752 11940 12756 11996
rect 12692 11936 12756 11940
rect 12772 11996 12836 12000
rect 12772 11940 12776 11996
rect 12776 11940 12832 11996
rect 12832 11940 12836 11996
rect 12772 11936 12836 11940
rect 12852 11996 12916 12000
rect 12852 11940 12856 11996
rect 12856 11940 12912 11996
rect 12912 11940 12916 11996
rect 12852 11936 12916 11940
rect 17612 11996 17676 12000
rect 17612 11940 17616 11996
rect 17616 11940 17672 11996
rect 17672 11940 17676 11996
rect 17612 11936 17676 11940
rect 17692 11996 17756 12000
rect 17692 11940 17696 11996
rect 17696 11940 17752 11996
rect 17752 11940 17756 11996
rect 17692 11936 17756 11940
rect 17772 11996 17836 12000
rect 17772 11940 17776 11996
rect 17776 11940 17832 11996
rect 17832 11940 17836 11996
rect 17772 11936 17836 11940
rect 17852 11996 17916 12000
rect 17852 11940 17856 11996
rect 17856 11940 17912 11996
rect 17912 11940 17916 11996
rect 17852 11936 17916 11940
rect 22612 11996 22676 12000
rect 22612 11940 22616 11996
rect 22616 11940 22672 11996
rect 22672 11940 22676 11996
rect 22612 11936 22676 11940
rect 22692 11996 22756 12000
rect 22692 11940 22696 11996
rect 22696 11940 22752 11996
rect 22752 11940 22756 11996
rect 22692 11936 22756 11940
rect 22772 11996 22836 12000
rect 22772 11940 22776 11996
rect 22776 11940 22832 11996
rect 22832 11940 22836 11996
rect 22772 11936 22836 11940
rect 22852 11996 22916 12000
rect 22852 11940 22856 11996
rect 22856 11940 22912 11996
rect 22912 11940 22916 11996
rect 22852 11936 22916 11940
rect 27612 11996 27676 12000
rect 27612 11940 27616 11996
rect 27616 11940 27672 11996
rect 27672 11940 27676 11996
rect 27612 11936 27676 11940
rect 27692 11996 27756 12000
rect 27692 11940 27696 11996
rect 27696 11940 27752 11996
rect 27752 11940 27756 11996
rect 27692 11936 27756 11940
rect 27772 11996 27836 12000
rect 27772 11940 27776 11996
rect 27776 11940 27832 11996
rect 27832 11940 27836 11996
rect 27772 11936 27836 11940
rect 27852 11996 27916 12000
rect 27852 11940 27856 11996
rect 27856 11940 27912 11996
rect 27912 11940 27916 11996
rect 27852 11936 27916 11940
rect 32612 11996 32676 12000
rect 32612 11940 32616 11996
rect 32616 11940 32672 11996
rect 32672 11940 32676 11996
rect 32612 11936 32676 11940
rect 32692 11996 32756 12000
rect 32692 11940 32696 11996
rect 32696 11940 32752 11996
rect 32752 11940 32756 11996
rect 32692 11936 32756 11940
rect 32772 11996 32836 12000
rect 32772 11940 32776 11996
rect 32776 11940 32832 11996
rect 32832 11940 32836 11996
rect 32772 11936 32836 11940
rect 32852 11996 32916 12000
rect 32852 11940 32856 11996
rect 32856 11940 32912 11996
rect 32912 11940 32916 11996
rect 32852 11936 32916 11940
rect 37612 11996 37676 12000
rect 37612 11940 37616 11996
rect 37616 11940 37672 11996
rect 37672 11940 37676 11996
rect 37612 11936 37676 11940
rect 37692 11996 37756 12000
rect 37692 11940 37696 11996
rect 37696 11940 37752 11996
rect 37752 11940 37756 11996
rect 37692 11936 37756 11940
rect 37772 11996 37836 12000
rect 37772 11940 37776 11996
rect 37776 11940 37832 11996
rect 37832 11940 37836 11996
rect 37772 11936 37836 11940
rect 37852 11996 37916 12000
rect 37852 11940 37856 11996
rect 37856 11940 37912 11996
rect 37912 11940 37916 11996
rect 37852 11936 37916 11940
rect 1952 11452 2016 11456
rect 1952 11396 1956 11452
rect 1956 11396 2012 11452
rect 2012 11396 2016 11452
rect 1952 11392 2016 11396
rect 2032 11452 2096 11456
rect 2032 11396 2036 11452
rect 2036 11396 2092 11452
rect 2092 11396 2096 11452
rect 2032 11392 2096 11396
rect 2112 11452 2176 11456
rect 2112 11396 2116 11452
rect 2116 11396 2172 11452
rect 2172 11396 2176 11452
rect 2112 11392 2176 11396
rect 2192 11452 2256 11456
rect 2192 11396 2196 11452
rect 2196 11396 2252 11452
rect 2252 11396 2256 11452
rect 2192 11392 2256 11396
rect 6952 11452 7016 11456
rect 6952 11396 6956 11452
rect 6956 11396 7012 11452
rect 7012 11396 7016 11452
rect 6952 11392 7016 11396
rect 7032 11452 7096 11456
rect 7032 11396 7036 11452
rect 7036 11396 7092 11452
rect 7092 11396 7096 11452
rect 7032 11392 7096 11396
rect 7112 11452 7176 11456
rect 7112 11396 7116 11452
rect 7116 11396 7172 11452
rect 7172 11396 7176 11452
rect 7112 11392 7176 11396
rect 7192 11452 7256 11456
rect 7192 11396 7196 11452
rect 7196 11396 7252 11452
rect 7252 11396 7256 11452
rect 7192 11392 7256 11396
rect 11952 11452 12016 11456
rect 11952 11396 11956 11452
rect 11956 11396 12012 11452
rect 12012 11396 12016 11452
rect 11952 11392 12016 11396
rect 12032 11452 12096 11456
rect 12032 11396 12036 11452
rect 12036 11396 12092 11452
rect 12092 11396 12096 11452
rect 12032 11392 12096 11396
rect 12112 11452 12176 11456
rect 12112 11396 12116 11452
rect 12116 11396 12172 11452
rect 12172 11396 12176 11452
rect 12112 11392 12176 11396
rect 12192 11452 12256 11456
rect 12192 11396 12196 11452
rect 12196 11396 12252 11452
rect 12252 11396 12256 11452
rect 12192 11392 12256 11396
rect 16952 11452 17016 11456
rect 16952 11396 16956 11452
rect 16956 11396 17012 11452
rect 17012 11396 17016 11452
rect 16952 11392 17016 11396
rect 17032 11452 17096 11456
rect 17032 11396 17036 11452
rect 17036 11396 17092 11452
rect 17092 11396 17096 11452
rect 17032 11392 17096 11396
rect 17112 11452 17176 11456
rect 17112 11396 17116 11452
rect 17116 11396 17172 11452
rect 17172 11396 17176 11452
rect 17112 11392 17176 11396
rect 17192 11452 17256 11456
rect 17192 11396 17196 11452
rect 17196 11396 17252 11452
rect 17252 11396 17256 11452
rect 17192 11392 17256 11396
rect 21952 11452 22016 11456
rect 21952 11396 21956 11452
rect 21956 11396 22012 11452
rect 22012 11396 22016 11452
rect 21952 11392 22016 11396
rect 22032 11452 22096 11456
rect 22032 11396 22036 11452
rect 22036 11396 22092 11452
rect 22092 11396 22096 11452
rect 22032 11392 22096 11396
rect 22112 11452 22176 11456
rect 22112 11396 22116 11452
rect 22116 11396 22172 11452
rect 22172 11396 22176 11452
rect 22112 11392 22176 11396
rect 22192 11452 22256 11456
rect 22192 11396 22196 11452
rect 22196 11396 22252 11452
rect 22252 11396 22256 11452
rect 22192 11392 22256 11396
rect 26952 11452 27016 11456
rect 26952 11396 26956 11452
rect 26956 11396 27012 11452
rect 27012 11396 27016 11452
rect 26952 11392 27016 11396
rect 27032 11452 27096 11456
rect 27032 11396 27036 11452
rect 27036 11396 27092 11452
rect 27092 11396 27096 11452
rect 27032 11392 27096 11396
rect 27112 11452 27176 11456
rect 27112 11396 27116 11452
rect 27116 11396 27172 11452
rect 27172 11396 27176 11452
rect 27112 11392 27176 11396
rect 27192 11452 27256 11456
rect 27192 11396 27196 11452
rect 27196 11396 27252 11452
rect 27252 11396 27256 11452
rect 27192 11392 27256 11396
rect 31952 11452 32016 11456
rect 31952 11396 31956 11452
rect 31956 11396 32012 11452
rect 32012 11396 32016 11452
rect 31952 11392 32016 11396
rect 32032 11452 32096 11456
rect 32032 11396 32036 11452
rect 32036 11396 32092 11452
rect 32092 11396 32096 11452
rect 32032 11392 32096 11396
rect 32112 11452 32176 11456
rect 32112 11396 32116 11452
rect 32116 11396 32172 11452
rect 32172 11396 32176 11452
rect 32112 11392 32176 11396
rect 32192 11452 32256 11456
rect 32192 11396 32196 11452
rect 32196 11396 32252 11452
rect 32252 11396 32256 11452
rect 32192 11392 32256 11396
rect 36952 11452 37016 11456
rect 36952 11396 36956 11452
rect 36956 11396 37012 11452
rect 37012 11396 37016 11452
rect 36952 11392 37016 11396
rect 37032 11452 37096 11456
rect 37032 11396 37036 11452
rect 37036 11396 37092 11452
rect 37092 11396 37096 11452
rect 37032 11392 37096 11396
rect 37112 11452 37176 11456
rect 37112 11396 37116 11452
rect 37116 11396 37172 11452
rect 37172 11396 37176 11452
rect 37112 11392 37176 11396
rect 37192 11452 37256 11456
rect 37192 11396 37196 11452
rect 37196 11396 37252 11452
rect 37252 11396 37256 11452
rect 37192 11392 37256 11396
rect 33180 10976 33244 10980
rect 33180 10920 33194 10976
rect 33194 10920 33244 10976
rect 33180 10916 33244 10920
rect 2612 10908 2676 10912
rect 2612 10852 2616 10908
rect 2616 10852 2672 10908
rect 2672 10852 2676 10908
rect 2612 10848 2676 10852
rect 2692 10908 2756 10912
rect 2692 10852 2696 10908
rect 2696 10852 2752 10908
rect 2752 10852 2756 10908
rect 2692 10848 2756 10852
rect 2772 10908 2836 10912
rect 2772 10852 2776 10908
rect 2776 10852 2832 10908
rect 2832 10852 2836 10908
rect 2772 10848 2836 10852
rect 2852 10908 2916 10912
rect 2852 10852 2856 10908
rect 2856 10852 2912 10908
rect 2912 10852 2916 10908
rect 2852 10848 2916 10852
rect 7612 10908 7676 10912
rect 7612 10852 7616 10908
rect 7616 10852 7672 10908
rect 7672 10852 7676 10908
rect 7612 10848 7676 10852
rect 7692 10908 7756 10912
rect 7692 10852 7696 10908
rect 7696 10852 7752 10908
rect 7752 10852 7756 10908
rect 7692 10848 7756 10852
rect 7772 10908 7836 10912
rect 7772 10852 7776 10908
rect 7776 10852 7832 10908
rect 7832 10852 7836 10908
rect 7772 10848 7836 10852
rect 7852 10908 7916 10912
rect 7852 10852 7856 10908
rect 7856 10852 7912 10908
rect 7912 10852 7916 10908
rect 7852 10848 7916 10852
rect 12612 10908 12676 10912
rect 12612 10852 12616 10908
rect 12616 10852 12672 10908
rect 12672 10852 12676 10908
rect 12612 10848 12676 10852
rect 12692 10908 12756 10912
rect 12692 10852 12696 10908
rect 12696 10852 12752 10908
rect 12752 10852 12756 10908
rect 12692 10848 12756 10852
rect 12772 10908 12836 10912
rect 12772 10852 12776 10908
rect 12776 10852 12832 10908
rect 12832 10852 12836 10908
rect 12772 10848 12836 10852
rect 12852 10908 12916 10912
rect 12852 10852 12856 10908
rect 12856 10852 12912 10908
rect 12912 10852 12916 10908
rect 12852 10848 12916 10852
rect 17612 10908 17676 10912
rect 17612 10852 17616 10908
rect 17616 10852 17672 10908
rect 17672 10852 17676 10908
rect 17612 10848 17676 10852
rect 17692 10908 17756 10912
rect 17692 10852 17696 10908
rect 17696 10852 17752 10908
rect 17752 10852 17756 10908
rect 17692 10848 17756 10852
rect 17772 10908 17836 10912
rect 17772 10852 17776 10908
rect 17776 10852 17832 10908
rect 17832 10852 17836 10908
rect 17772 10848 17836 10852
rect 17852 10908 17916 10912
rect 17852 10852 17856 10908
rect 17856 10852 17912 10908
rect 17912 10852 17916 10908
rect 17852 10848 17916 10852
rect 22612 10908 22676 10912
rect 22612 10852 22616 10908
rect 22616 10852 22672 10908
rect 22672 10852 22676 10908
rect 22612 10848 22676 10852
rect 22692 10908 22756 10912
rect 22692 10852 22696 10908
rect 22696 10852 22752 10908
rect 22752 10852 22756 10908
rect 22692 10848 22756 10852
rect 22772 10908 22836 10912
rect 22772 10852 22776 10908
rect 22776 10852 22832 10908
rect 22832 10852 22836 10908
rect 22772 10848 22836 10852
rect 22852 10908 22916 10912
rect 22852 10852 22856 10908
rect 22856 10852 22912 10908
rect 22912 10852 22916 10908
rect 22852 10848 22916 10852
rect 27612 10908 27676 10912
rect 27612 10852 27616 10908
rect 27616 10852 27672 10908
rect 27672 10852 27676 10908
rect 27612 10848 27676 10852
rect 27692 10908 27756 10912
rect 27692 10852 27696 10908
rect 27696 10852 27752 10908
rect 27752 10852 27756 10908
rect 27692 10848 27756 10852
rect 27772 10908 27836 10912
rect 27772 10852 27776 10908
rect 27776 10852 27832 10908
rect 27832 10852 27836 10908
rect 27772 10848 27836 10852
rect 27852 10908 27916 10912
rect 27852 10852 27856 10908
rect 27856 10852 27912 10908
rect 27912 10852 27916 10908
rect 27852 10848 27916 10852
rect 32612 10908 32676 10912
rect 32612 10852 32616 10908
rect 32616 10852 32672 10908
rect 32672 10852 32676 10908
rect 32612 10848 32676 10852
rect 32692 10908 32756 10912
rect 32692 10852 32696 10908
rect 32696 10852 32752 10908
rect 32752 10852 32756 10908
rect 32692 10848 32756 10852
rect 32772 10908 32836 10912
rect 32772 10852 32776 10908
rect 32776 10852 32832 10908
rect 32832 10852 32836 10908
rect 32772 10848 32836 10852
rect 32852 10908 32916 10912
rect 32852 10852 32856 10908
rect 32856 10852 32912 10908
rect 32912 10852 32916 10908
rect 32852 10848 32916 10852
rect 37612 10908 37676 10912
rect 37612 10852 37616 10908
rect 37616 10852 37672 10908
rect 37672 10852 37676 10908
rect 37612 10848 37676 10852
rect 37692 10908 37756 10912
rect 37692 10852 37696 10908
rect 37696 10852 37752 10908
rect 37752 10852 37756 10908
rect 37692 10848 37756 10852
rect 37772 10908 37836 10912
rect 37772 10852 37776 10908
rect 37776 10852 37832 10908
rect 37832 10852 37836 10908
rect 37772 10848 37836 10852
rect 37852 10908 37916 10912
rect 37852 10852 37856 10908
rect 37856 10852 37912 10908
rect 37912 10852 37916 10908
rect 37852 10848 37916 10852
rect 1952 10364 2016 10368
rect 1952 10308 1956 10364
rect 1956 10308 2012 10364
rect 2012 10308 2016 10364
rect 1952 10304 2016 10308
rect 2032 10364 2096 10368
rect 2032 10308 2036 10364
rect 2036 10308 2092 10364
rect 2092 10308 2096 10364
rect 2032 10304 2096 10308
rect 2112 10364 2176 10368
rect 2112 10308 2116 10364
rect 2116 10308 2172 10364
rect 2172 10308 2176 10364
rect 2112 10304 2176 10308
rect 2192 10364 2256 10368
rect 2192 10308 2196 10364
rect 2196 10308 2252 10364
rect 2252 10308 2256 10364
rect 2192 10304 2256 10308
rect 6952 10364 7016 10368
rect 6952 10308 6956 10364
rect 6956 10308 7012 10364
rect 7012 10308 7016 10364
rect 6952 10304 7016 10308
rect 7032 10364 7096 10368
rect 7032 10308 7036 10364
rect 7036 10308 7092 10364
rect 7092 10308 7096 10364
rect 7032 10304 7096 10308
rect 7112 10364 7176 10368
rect 7112 10308 7116 10364
rect 7116 10308 7172 10364
rect 7172 10308 7176 10364
rect 7112 10304 7176 10308
rect 7192 10364 7256 10368
rect 7192 10308 7196 10364
rect 7196 10308 7252 10364
rect 7252 10308 7256 10364
rect 7192 10304 7256 10308
rect 11952 10364 12016 10368
rect 11952 10308 11956 10364
rect 11956 10308 12012 10364
rect 12012 10308 12016 10364
rect 11952 10304 12016 10308
rect 12032 10364 12096 10368
rect 12032 10308 12036 10364
rect 12036 10308 12092 10364
rect 12092 10308 12096 10364
rect 12032 10304 12096 10308
rect 12112 10364 12176 10368
rect 12112 10308 12116 10364
rect 12116 10308 12172 10364
rect 12172 10308 12176 10364
rect 12112 10304 12176 10308
rect 12192 10364 12256 10368
rect 12192 10308 12196 10364
rect 12196 10308 12252 10364
rect 12252 10308 12256 10364
rect 12192 10304 12256 10308
rect 16952 10364 17016 10368
rect 16952 10308 16956 10364
rect 16956 10308 17012 10364
rect 17012 10308 17016 10364
rect 16952 10304 17016 10308
rect 17032 10364 17096 10368
rect 17032 10308 17036 10364
rect 17036 10308 17092 10364
rect 17092 10308 17096 10364
rect 17032 10304 17096 10308
rect 17112 10364 17176 10368
rect 17112 10308 17116 10364
rect 17116 10308 17172 10364
rect 17172 10308 17176 10364
rect 17112 10304 17176 10308
rect 17192 10364 17256 10368
rect 17192 10308 17196 10364
rect 17196 10308 17252 10364
rect 17252 10308 17256 10364
rect 17192 10304 17256 10308
rect 21952 10364 22016 10368
rect 21952 10308 21956 10364
rect 21956 10308 22012 10364
rect 22012 10308 22016 10364
rect 21952 10304 22016 10308
rect 22032 10364 22096 10368
rect 22032 10308 22036 10364
rect 22036 10308 22092 10364
rect 22092 10308 22096 10364
rect 22032 10304 22096 10308
rect 22112 10364 22176 10368
rect 22112 10308 22116 10364
rect 22116 10308 22172 10364
rect 22172 10308 22176 10364
rect 22112 10304 22176 10308
rect 22192 10364 22256 10368
rect 22192 10308 22196 10364
rect 22196 10308 22252 10364
rect 22252 10308 22256 10364
rect 22192 10304 22256 10308
rect 26952 10364 27016 10368
rect 26952 10308 26956 10364
rect 26956 10308 27012 10364
rect 27012 10308 27016 10364
rect 26952 10304 27016 10308
rect 27032 10364 27096 10368
rect 27032 10308 27036 10364
rect 27036 10308 27092 10364
rect 27092 10308 27096 10364
rect 27032 10304 27096 10308
rect 27112 10364 27176 10368
rect 27112 10308 27116 10364
rect 27116 10308 27172 10364
rect 27172 10308 27176 10364
rect 27112 10304 27176 10308
rect 27192 10364 27256 10368
rect 27192 10308 27196 10364
rect 27196 10308 27252 10364
rect 27252 10308 27256 10364
rect 27192 10304 27256 10308
rect 31952 10364 32016 10368
rect 31952 10308 31956 10364
rect 31956 10308 32012 10364
rect 32012 10308 32016 10364
rect 31952 10304 32016 10308
rect 32032 10364 32096 10368
rect 32032 10308 32036 10364
rect 32036 10308 32092 10364
rect 32092 10308 32096 10364
rect 32032 10304 32096 10308
rect 32112 10364 32176 10368
rect 32112 10308 32116 10364
rect 32116 10308 32172 10364
rect 32172 10308 32176 10364
rect 32112 10304 32176 10308
rect 32192 10364 32256 10368
rect 32192 10308 32196 10364
rect 32196 10308 32252 10364
rect 32252 10308 32256 10364
rect 32192 10304 32256 10308
rect 36952 10364 37016 10368
rect 36952 10308 36956 10364
rect 36956 10308 37012 10364
rect 37012 10308 37016 10364
rect 36952 10304 37016 10308
rect 37032 10364 37096 10368
rect 37032 10308 37036 10364
rect 37036 10308 37092 10364
rect 37092 10308 37096 10364
rect 37032 10304 37096 10308
rect 37112 10364 37176 10368
rect 37112 10308 37116 10364
rect 37116 10308 37172 10364
rect 37172 10308 37176 10364
rect 37112 10304 37176 10308
rect 37192 10364 37256 10368
rect 37192 10308 37196 10364
rect 37196 10308 37252 10364
rect 37252 10308 37256 10364
rect 37192 10304 37256 10308
rect 2612 9820 2676 9824
rect 2612 9764 2616 9820
rect 2616 9764 2672 9820
rect 2672 9764 2676 9820
rect 2612 9760 2676 9764
rect 2692 9820 2756 9824
rect 2692 9764 2696 9820
rect 2696 9764 2752 9820
rect 2752 9764 2756 9820
rect 2692 9760 2756 9764
rect 2772 9820 2836 9824
rect 2772 9764 2776 9820
rect 2776 9764 2832 9820
rect 2832 9764 2836 9820
rect 2772 9760 2836 9764
rect 2852 9820 2916 9824
rect 2852 9764 2856 9820
rect 2856 9764 2912 9820
rect 2912 9764 2916 9820
rect 2852 9760 2916 9764
rect 7612 9820 7676 9824
rect 7612 9764 7616 9820
rect 7616 9764 7672 9820
rect 7672 9764 7676 9820
rect 7612 9760 7676 9764
rect 7692 9820 7756 9824
rect 7692 9764 7696 9820
rect 7696 9764 7752 9820
rect 7752 9764 7756 9820
rect 7692 9760 7756 9764
rect 7772 9820 7836 9824
rect 7772 9764 7776 9820
rect 7776 9764 7832 9820
rect 7832 9764 7836 9820
rect 7772 9760 7836 9764
rect 7852 9820 7916 9824
rect 7852 9764 7856 9820
rect 7856 9764 7912 9820
rect 7912 9764 7916 9820
rect 7852 9760 7916 9764
rect 12612 9820 12676 9824
rect 12612 9764 12616 9820
rect 12616 9764 12672 9820
rect 12672 9764 12676 9820
rect 12612 9760 12676 9764
rect 12692 9820 12756 9824
rect 12692 9764 12696 9820
rect 12696 9764 12752 9820
rect 12752 9764 12756 9820
rect 12692 9760 12756 9764
rect 12772 9820 12836 9824
rect 12772 9764 12776 9820
rect 12776 9764 12832 9820
rect 12832 9764 12836 9820
rect 12772 9760 12836 9764
rect 12852 9820 12916 9824
rect 12852 9764 12856 9820
rect 12856 9764 12912 9820
rect 12912 9764 12916 9820
rect 12852 9760 12916 9764
rect 17612 9820 17676 9824
rect 17612 9764 17616 9820
rect 17616 9764 17672 9820
rect 17672 9764 17676 9820
rect 17612 9760 17676 9764
rect 17692 9820 17756 9824
rect 17692 9764 17696 9820
rect 17696 9764 17752 9820
rect 17752 9764 17756 9820
rect 17692 9760 17756 9764
rect 17772 9820 17836 9824
rect 17772 9764 17776 9820
rect 17776 9764 17832 9820
rect 17832 9764 17836 9820
rect 17772 9760 17836 9764
rect 17852 9820 17916 9824
rect 17852 9764 17856 9820
rect 17856 9764 17912 9820
rect 17912 9764 17916 9820
rect 17852 9760 17916 9764
rect 22612 9820 22676 9824
rect 22612 9764 22616 9820
rect 22616 9764 22672 9820
rect 22672 9764 22676 9820
rect 22612 9760 22676 9764
rect 22692 9820 22756 9824
rect 22692 9764 22696 9820
rect 22696 9764 22752 9820
rect 22752 9764 22756 9820
rect 22692 9760 22756 9764
rect 22772 9820 22836 9824
rect 22772 9764 22776 9820
rect 22776 9764 22832 9820
rect 22832 9764 22836 9820
rect 22772 9760 22836 9764
rect 22852 9820 22916 9824
rect 22852 9764 22856 9820
rect 22856 9764 22912 9820
rect 22912 9764 22916 9820
rect 22852 9760 22916 9764
rect 27612 9820 27676 9824
rect 27612 9764 27616 9820
rect 27616 9764 27672 9820
rect 27672 9764 27676 9820
rect 27612 9760 27676 9764
rect 27692 9820 27756 9824
rect 27692 9764 27696 9820
rect 27696 9764 27752 9820
rect 27752 9764 27756 9820
rect 27692 9760 27756 9764
rect 27772 9820 27836 9824
rect 27772 9764 27776 9820
rect 27776 9764 27832 9820
rect 27832 9764 27836 9820
rect 27772 9760 27836 9764
rect 27852 9820 27916 9824
rect 27852 9764 27856 9820
rect 27856 9764 27912 9820
rect 27912 9764 27916 9820
rect 27852 9760 27916 9764
rect 32612 9820 32676 9824
rect 32612 9764 32616 9820
rect 32616 9764 32672 9820
rect 32672 9764 32676 9820
rect 32612 9760 32676 9764
rect 32692 9820 32756 9824
rect 32692 9764 32696 9820
rect 32696 9764 32752 9820
rect 32752 9764 32756 9820
rect 32692 9760 32756 9764
rect 32772 9820 32836 9824
rect 32772 9764 32776 9820
rect 32776 9764 32832 9820
rect 32832 9764 32836 9820
rect 32772 9760 32836 9764
rect 32852 9820 32916 9824
rect 32852 9764 32856 9820
rect 32856 9764 32912 9820
rect 32912 9764 32916 9820
rect 32852 9760 32916 9764
rect 37612 9820 37676 9824
rect 37612 9764 37616 9820
rect 37616 9764 37672 9820
rect 37672 9764 37676 9820
rect 37612 9760 37676 9764
rect 37692 9820 37756 9824
rect 37692 9764 37696 9820
rect 37696 9764 37752 9820
rect 37752 9764 37756 9820
rect 37692 9760 37756 9764
rect 37772 9820 37836 9824
rect 37772 9764 37776 9820
rect 37776 9764 37832 9820
rect 37832 9764 37836 9820
rect 37772 9760 37836 9764
rect 37852 9820 37916 9824
rect 37852 9764 37856 9820
rect 37856 9764 37912 9820
rect 37912 9764 37916 9820
rect 37852 9760 37916 9764
rect 33364 9556 33428 9620
rect 1952 9276 2016 9280
rect 1952 9220 1956 9276
rect 1956 9220 2012 9276
rect 2012 9220 2016 9276
rect 1952 9216 2016 9220
rect 2032 9276 2096 9280
rect 2032 9220 2036 9276
rect 2036 9220 2092 9276
rect 2092 9220 2096 9276
rect 2032 9216 2096 9220
rect 2112 9276 2176 9280
rect 2112 9220 2116 9276
rect 2116 9220 2172 9276
rect 2172 9220 2176 9276
rect 2112 9216 2176 9220
rect 2192 9276 2256 9280
rect 2192 9220 2196 9276
rect 2196 9220 2252 9276
rect 2252 9220 2256 9276
rect 2192 9216 2256 9220
rect 6952 9276 7016 9280
rect 6952 9220 6956 9276
rect 6956 9220 7012 9276
rect 7012 9220 7016 9276
rect 6952 9216 7016 9220
rect 7032 9276 7096 9280
rect 7032 9220 7036 9276
rect 7036 9220 7092 9276
rect 7092 9220 7096 9276
rect 7032 9216 7096 9220
rect 7112 9276 7176 9280
rect 7112 9220 7116 9276
rect 7116 9220 7172 9276
rect 7172 9220 7176 9276
rect 7112 9216 7176 9220
rect 7192 9276 7256 9280
rect 7192 9220 7196 9276
rect 7196 9220 7252 9276
rect 7252 9220 7256 9276
rect 7192 9216 7256 9220
rect 11952 9276 12016 9280
rect 11952 9220 11956 9276
rect 11956 9220 12012 9276
rect 12012 9220 12016 9276
rect 11952 9216 12016 9220
rect 12032 9276 12096 9280
rect 12032 9220 12036 9276
rect 12036 9220 12092 9276
rect 12092 9220 12096 9276
rect 12032 9216 12096 9220
rect 12112 9276 12176 9280
rect 12112 9220 12116 9276
rect 12116 9220 12172 9276
rect 12172 9220 12176 9276
rect 12112 9216 12176 9220
rect 12192 9276 12256 9280
rect 12192 9220 12196 9276
rect 12196 9220 12252 9276
rect 12252 9220 12256 9276
rect 12192 9216 12256 9220
rect 16952 9276 17016 9280
rect 16952 9220 16956 9276
rect 16956 9220 17012 9276
rect 17012 9220 17016 9276
rect 16952 9216 17016 9220
rect 17032 9276 17096 9280
rect 17032 9220 17036 9276
rect 17036 9220 17092 9276
rect 17092 9220 17096 9276
rect 17032 9216 17096 9220
rect 17112 9276 17176 9280
rect 17112 9220 17116 9276
rect 17116 9220 17172 9276
rect 17172 9220 17176 9276
rect 17112 9216 17176 9220
rect 17192 9276 17256 9280
rect 17192 9220 17196 9276
rect 17196 9220 17252 9276
rect 17252 9220 17256 9276
rect 17192 9216 17256 9220
rect 21952 9276 22016 9280
rect 21952 9220 21956 9276
rect 21956 9220 22012 9276
rect 22012 9220 22016 9276
rect 21952 9216 22016 9220
rect 22032 9276 22096 9280
rect 22032 9220 22036 9276
rect 22036 9220 22092 9276
rect 22092 9220 22096 9276
rect 22032 9216 22096 9220
rect 22112 9276 22176 9280
rect 22112 9220 22116 9276
rect 22116 9220 22172 9276
rect 22172 9220 22176 9276
rect 22112 9216 22176 9220
rect 22192 9276 22256 9280
rect 22192 9220 22196 9276
rect 22196 9220 22252 9276
rect 22252 9220 22256 9276
rect 22192 9216 22256 9220
rect 26952 9276 27016 9280
rect 26952 9220 26956 9276
rect 26956 9220 27012 9276
rect 27012 9220 27016 9276
rect 26952 9216 27016 9220
rect 27032 9276 27096 9280
rect 27032 9220 27036 9276
rect 27036 9220 27092 9276
rect 27092 9220 27096 9276
rect 27032 9216 27096 9220
rect 27112 9276 27176 9280
rect 27112 9220 27116 9276
rect 27116 9220 27172 9276
rect 27172 9220 27176 9276
rect 27112 9216 27176 9220
rect 27192 9276 27256 9280
rect 27192 9220 27196 9276
rect 27196 9220 27252 9276
rect 27252 9220 27256 9276
rect 27192 9216 27256 9220
rect 31952 9276 32016 9280
rect 31952 9220 31956 9276
rect 31956 9220 32012 9276
rect 32012 9220 32016 9276
rect 31952 9216 32016 9220
rect 32032 9276 32096 9280
rect 32032 9220 32036 9276
rect 32036 9220 32092 9276
rect 32092 9220 32096 9276
rect 32032 9216 32096 9220
rect 32112 9276 32176 9280
rect 32112 9220 32116 9276
rect 32116 9220 32172 9276
rect 32172 9220 32176 9276
rect 32112 9216 32176 9220
rect 32192 9276 32256 9280
rect 32192 9220 32196 9276
rect 32196 9220 32252 9276
rect 32252 9220 32256 9276
rect 32192 9216 32256 9220
rect 36952 9276 37016 9280
rect 36952 9220 36956 9276
rect 36956 9220 37012 9276
rect 37012 9220 37016 9276
rect 36952 9216 37016 9220
rect 37032 9276 37096 9280
rect 37032 9220 37036 9276
rect 37036 9220 37092 9276
rect 37092 9220 37096 9276
rect 37032 9216 37096 9220
rect 37112 9276 37176 9280
rect 37112 9220 37116 9276
rect 37116 9220 37172 9276
rect 37172 9220 37176 9276
rect 37112 9216 37176 9220
rect 37192 9276 37256 9280
rect 37192 9220 37196 9276
rect 37196 9220 37252 9276
rect 37252 9220 37256 9276
rect 37192 9216 37256 9220
rect 2612 8732 2676 8736
rect 2612 8676 2616 8732
rect 2616 8676 2672 8732
rect 2672 8676 2676 8732
rect 2612 8672 2676 8676
rect 2692 8732 2756 8736
rect 2692 8676 2696 8732
rect 2696 8676 2752 8732
rect 2752 8676 2756 8732
rect 2692 8672 2756 8676
rect 2772 8732 2836 8736
rect 2772 8676 2776 8732
rect 2776 8676 2832 8732
rect 2832 8676 2836 8732
rect 2772 8672 2836 8676
rect 2852 8732 2916 8736
rect 2852 8676 2856 8732
rect 2856 8676 2912 8732
rect 2912 8676 2916 8732
rect 2852 8672 2916 8676
rect 7612 8732 7676 8736
rect 7612 8676 7616 8732
rect 7616 8676 7672 8732
rect 7672 8676 7676 8732
rect 7612 8672 7676 8676
rect 7692 8732 7756 8736
rect 7692 8676 7696 8732
rect 7696 8676 7752 8732
rect 7752 8676 7756 8732
rect 7692 8672 7756 8676
rect 7772 8732 7836 8736
rect 7772 8676 7776 8732
rect 7776 8676 7832 8732
rect 7832 8676 7836 8732
rect 7772 8672 7836 8676
rect 7852 8732 7916 8736
rect 7852 8676 7856 8732
rect 7856 8676 7912 8732
rect 7912 8676 7916 8732
rect 7852 8672 7916 8676
rect 12612 8732 12676 8736
rect 12612 8676 12616 8732
rect 12616 8676 12672 8732
rect 12672 8676 12676 8732
rect 12612 8672 12676 8676
rect 12692 8732 12756 8736
rect 12692 8676 12696 8732
rect 12696 8676 12752 8732
rect 12752 8676 12756 8732
rect 12692 8672 12756 8676
rect 12772 8732 12836 8736
rect 12772 8676 12776 8732
rect 12776 8676 12832 8732
rect 12832 8676 12836 8732
rect 12772 8672 12836 8676
rect 12852 8732 12916 8736
rect 12852 8676 12856 8732
rect 12856 8676 12912 8732
rect 12912 8676 12916 8732
rect 12852 8672 12916 8676
rect 17612 8732 17676 8736
rect 17612 8676 17616 8732
rect 17616 8676 17672 8732
rect 17672 8676 17676 8732
rect 17612 8672 17676 8676
rect 17692 8732 17756 8736
rect 17692 8676 17696 8732
rect 17696 8676 17752 8732
rect 17752 8676 17756 8732
rect 17692 8672 17756 8676
rect 17772 8732 17836 8736
rect 17772 8676 17776 8732
rect 17776 8676 17832 8732
rect 17832 8676 17836 8732
rect 17772 8672 17836 8676
rect 17852 8732 17916 8736
rect 17852 8676 17856 8732
rect 17856 8676 17912 8732
rect 17912 8676 17916 8732
rect 17852 8672 17916 8676
rect 22612 8732 22676 8736
rect 22612 8676 22616 8732
rect 22616 8676 22672 8732
rect 22672 8676 22676 8732
rect 22612 8672 22676 8676
rect 22692 8732 22756 8736
rect 22692 8676 22696 8732
rect 22696 8676 22752 8732
rect 22752 8676 22756 8732
rect 22692 8672 22756 8676
rect 22772 8732 22836 8736
rect 22772 8676 22776 8732
rect 22776 8676 22832 8732
rect 22832 8676 22836 8732
rect 22772 8672 22836 8676
rect 22852 8732 22916 8736
rect 22852 8676 22856 8732
rect 22856 8676 22912 8732
rect 22912 8676 22916 8732
rect 22852 8672 22916 8676
rect 27612 8732 27676 8736
rect 27612 8676 27616 8732
rect 27616 8676 27672 8732
rect 27672 8676 27676 8732
rect 27612 8672 27676 8676
rect 27692 8732 27756 8736
rect 27692 8676 27696 8732
rect 27696 8676 27752 8732
rect 27752 8676 27756 8732
rect 27692 8672 27756 8676
rect 27772 8732 27836 8736
rect 27772 8676 27776 8732
rect 27776 8676 27832 8732
rect 27832 8676 27836 8732
rect 27772 8672 27836 8676
rect 27852 8732 27916 8736
rect 27852 8676 27856 8732
rect 27856 8676 27912 8732
rect 27912 8676 27916 8732
rect 27852 8672 27916 8676
rect 32612 8732 32676 8736
rect 32612 8676 32616 8732
rect 32616 8676 32672 8732
rect 32672 8676 32676 8732
rect 32612 8672 32676 8676
rect 32692 8732 32756 8736
rect 32692 8676 32696 8732
rect 32696 8676 32752 8732
rect 32752 8676 32756 8732
rect 32692 8672 32756 8676
rect 32772 8732 32836 8736
rect 32772 8676 32776 8732
rect 32776 8676 32832 8732
rect 32832 8676 32836 8732
rect 32772 8672 32836 8676
rect 32852 8732 32916 8736
rect 32852 8676 32856 8732
rect 32856 8676 32912 8732
rect 32912 8676 32916 8732
rect 32852 8672 32916 8676
rect 37612 8732 37676 8736
rect 37612 8676 37616 8732
rect 37616 8676 37672 8732
rect 37672 8676 37676 8732
rect 37612 8672 37676 8676
rect 37692 8732 37756 8736
rect 37692 8676 37696 8732
rect 37696 8676 37752 8732
rect 37752 8676 37756 8732
rect 37692 8672 37756 8676
rect 37772 8732 37836 8736
rect 37772 8676 37776 8732
rect 37776 8676 37832 8732
rect 37832 8676 37836 8732
rect 37772 8672 37836 8676
rect 37852 8732 37916 8736
rect 37852 8676 37856 8732
rect 37856 8676 37912 8732
rect 37912 8676 37916 8732
rect 37852 8672 37916 8676
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 6952 8188 7016 8192
rect 6952 8132 6956 8188
rect 6956 8132 7012 8188
rect 7012 8132 7016 8188
rect 6952 8128 7016 8132
rect 7032 8188 7096 8192
rect 7032 8132 7036 8188
rect 7036 8132 7092 8188
rect 7092 8132 7096 8188
rect 7032 8128 7096 8132
rect 7112 8188 7176 8192
rect 7112 8132 7116 8188
rect 7116 8132 7172 8188
rect 7172 8132 7176 8188
rect 7112 8128 7176 8132
rect 7192 8188 7256 8192
rect 7192 8132 7196 8188
rect 7196 8132 7252 8188
rect 7252 8132 7256 8188
rect 7192 8128 7256 8132
rect 11952 8188 12016 8192
rect 11952 8132 11956 8188
rect 11956 8132 12012 8188
rect 12012 8132 12016 8188
rect 11952 8128 12016 8132
rect 12032 8188 12096 8192
rect 12032 8132 12036 8188
rect 12036 8132 12092 8188
rect 12092 8132 12096 8188
rect 12032 8128 12096 8132
rect 12112 8188 12176 8192
rect 12112 8132 12116 8188
rect 12116 8132 12172 8188
rect 12172 8132 12176 8188
rect 12112 8128 12176 8132
rect 12192 8188 12256 8192
rect 12192 8132 12196 8188
rect 12196 8132 12252 8188
rect 12252 8132 12256 8188
rect 12192 8128 12256 8132
rect 16952 8188 17016 8192
rect 16952 8132 16956 8188
rect 16956 8132 17012 8188
rect 17012 8132 17016 8188
rect 16952 8128 17016 8132
rect 17032 8188 17096 8192
rect 17032 8132 17036 8188
rect 17036 8132 17092 8188
rect 17092 8132 17096 8188
rect 17032 8128 17096 8132
rect 17112 8188 17176 8192
rect 17112 8132 17116 8188
rect 17116 8132 17172 8188
rect 17172 8132 17176 8188
rect 17112 8128 17176 8132
rect 17192 8188 17256 8192
rect 17192 8132 17196 8188
rect 17196 8132 17252 8188
rect 17252 8132 17256 8188
rect 17192 8128 17256 8132
rect 21952 8188 22016 8192
rect 21952 8132 21956 8188
rect 21956 8132 22012 8188
rect 22012 8132 22016 8188
rect 21952 8128 22016 8132
rect 22032 8188 22096 8192
rect 22032 8132 22036 8188
rect 22036 8132 22092 8188
rect 22092 8132 22096 8188
rect 22032 8128 22096 8132
rect 22112 8188 22176 8192
rect 22112 8132 22116 8188
rect 22116 8132 22172 8188
rect 22172 8132 22176 8188
rect 22112 8128 22176 8132
rect 22192 8188 22256 8192
rect 22192 8132 22196 8188
rect 22196 8132 22252 8188
rect 22252 8132 22256 8188
rect 22192 8128 22256 8132
rect 26952 8188 27016 8192
rect 26952 8132 26956 8188
rect 26956 8132 27012 8188
rect 27012 8132 27016 8188
rect 26952 8128 27016 8132
rect 27032 8188 27096 8192
rect 27032 8132 27036 8188
rect 27036 8132 27092 8188
rect 27092 8132 27096 8188
rect 27032 8128 27096 8132
rect 27112 8188 27176 8192
rect 27112 8132 27116 8188
rect 27116 8132 27172 8188
rect 27172 8132 27176 8188
rect 27112 8128 27176 8132
rect 27192 8188 27256 8192
rect 27192 8132 27196 8188
rect 27196 8132 27252 8188
rect 27252 8132 27256 8188
rect 27192 8128 27256 8132
rect 31952 8188 32016 8192
rect 31952 8132 31956 8188
rect 31956 8132 32012 8188
rect 32012 8132 32016 8188
rect 31952 8128 32016 8132
rect 32032 8188 32096 8192
rect 32032 8132 32036 8188
rect 32036 8132 32092 8188
rect 32092 8132 32096 8188
rect 32032 8128 32096 8132
rect 32112 8188 32176 8192
rect 32112 8132 32116 8188
rect 32116 8132 32172 8188
rect 32172 8132 32176 8188
rect 32112 8128 32176 8132
rect 32192 8188 32256 8192
rect 32192 8132 32196 8188
rect 32196 8132 32252 8188
rect 32252 8132 32256 8188
rect 32192 8128 32256 8132
rect 36952 8188 37016 8192
rect 36952 8132 36956 8188
rect 36956 8132 37012 8188
rect 37012 8132 37016 8188
rect 36952 8128 37016 8132
rect 37032 8188 37096 8192
rect 37032 8132 37036 8188
rect 37036 8132 37092 8188
rect 37092 8132 37096 8188
rect 37032 8128 37096 8132
rect 37112 8188 37176 8192
rect 37112 8132 37116 8188
rect 37116 8132 37172 8188
rect 37172 8132 37176 8188
rect 37112 8128 37176 8132
rect 37192 8188 37256 8192
rect 37192 8132 37196 8188
rect 37196 8132 37252 8188
rect 37252 8132 37256 8188
rect 37192 8128 37256 8132
rect 33548 7788 33612 7852
rect 2612 7644 2676 7648
rect 2612 7588 2616 7644
rect 2616 7588 2672 7644
rect 2672 7588 2676 7644
rect 2612 7584 2676 7588
rect 2692 7644 2756 7648
rect 2692 7588 2696 7644
rect 2696 7588 2752 7644
rect 2752 7588 2756 7644
rect 2692 7584 2756 7588
rect 2772 7644 2836 7648
rect 2772 7588 2776 7644
rect 2776 7588 2832 7644
rect 2832 7588 2836 7644
rect 2772 7584 2836 7588
rect 2852 7644 2916 7648
rect 2852 7588 2856 7644
rect 2856 7588 2912 7644
rect 2912 7588 2916 7644
rect 2852 7584 2916 7588
rect 7612 7644 7676 7648
rect 7612 7588 7616 7644
rect 7616 7588 7672 7644
rect 7672 7588 7676 7644
rect 7612 7584 7676 7588
rect 7692 7644 7756 7648
rect 7692 7588 7696 7644
rect 7696 7588 7752 7644
rect 7752 7588 7756 7644
rect 7692 7584 7756 7588
rect 7772 7644 7836 7648
rect 7772 7588 7776 7644
rect 7776 7588 7832 7644
rect 7832 7588 7836 7644
rect 7772 7584 7836 7588
rect 7852 7644 7916 7648
rect 7852 7588 7856 7644
rect 7856 7588 7912 7644
rect 7912 7588 7916 7644
rect 7852 7584 7916 7588
rect 12612 7644 12676 7648
rect 12612 7588 12616 7644
rect 12616 7588 12672 7644
rect 12672 7588 12676 7644
rect 12612 7584 12676 7588
rect 12692 7644 12756 7648
rect 12692 7588 12696 7644
rect 12696 7588 12752 7644
rect 12752 7588 12756 7644
rect 12692 7584 12756 7588
rect 12772 7644 12836 7648
rect 12772 7588 12776 7644
rect 12776 7588 12832 7644
rect 12832 7588 12836 7644
rect 12772 7584 12836 7588
rect 12852 7644 12916 7648
rect 12852 7588 12856 7644
rect 12856 7588 12912 7644
rect 12912 7588 12916 7644
rect 12852 7584 12916 7588
rect 17612 7644 17676 7648
rect 17612 7588 17616 7644
rect 17616 7588 17672 7644
rect 17672 7588 17676 7644
rect 17612 7584 17676 7588
rect 17692 7644 17756 7648
rect 17692 7588 17696 7644
rect 17696 7588 17752 7644
rect 17752 7588 17756 7644
rect 17692 7584 17756 7588
rect 17772 7644 17836 7648
rect 17772 7588 17776 7644
rect 17776 7588 17832 7644
rect 17832 7588 17836 7644
rect 17772 7584 17836 7588
rect 17852 7644 17916 7648
rect 17852 7588 17856 7644
rect 17856 7588 17912 7644
rect 17912 7588 17916 7644
rect 17852 7584 17916 7588
rect 22612 7644 22676 7648
rect 22612 7588 22616 7644
rect 22616 7588 22672 7644
rect 22672 7588 22676 7644
rect 22612 7584 22676 7588
rect 22692 7644 22756 7648
rect 22692 7588 22696 7644
rect 22696 7588 22752 7644
rect 22752 7588 22756 7644
rect 22692 7584 22756 7588
rect 22772 7644 22836 7648
rect 22772 7588 22776 7644
rect 22776 7588 22832 7644
rect 22832 7588 22836 7644
rect 22772 7584 22836 7588
rect 22852 7644 22916 7648
rect 22852 7588 22856 7644
rect 22856 7588 22912 7644
rect 22912 7588 22916 7644
rect 22852 7584 22916 7588
rect 27612 7644 27676 7648
rect 27612 7588 27616 7644
rect 27616 7588 27672 7644
rect 27672 7588 27676 7644
rect 27612 7584 27676 7588
rect 27692 7644 27756 7648
rect 27692 7588 27696 7644
rect 27696 7588 27752 7644
rect 27752 7588 27756 7644
rect 27692 7584 27756 7588
rect 27772 7644 27836 7648
rect 27772 7588 27776 7644
rect 27776 7588 27832 7644
rect 27832 7588 27836 7644
rect 27772 7584 27836 7588
rect 27852 7644 27916 7648
rect 27852 7588 27856 7644
rect 27856 7588 27912 7644
rect 27912 7588 27916 7644
rect 27852 7584 27916 7588
rect 32612 7644 32676 7648
rect 32612 7588 32616 7644
rect 32616 7588 32672 7644
rect 32672 7588 32676 7644
rect 32612 7584 32676 7588
rect 32692 7644 32756 7648
rect 32692 7588 32696 7644
rect 32696 7588 32752 7644
rect 32752 7588 32756 7644
rect 32692 7584 32756 7588
rect 32772 7644 32836 7648
rect 32772 7588 32776 7644
rect 32776 7588 32832 7644
rect 32832 7588 32836 7644
rect 32772 7584 32836 7588
rect 32852 7644 32916 7648
rect 32852 7588 32856 7644
rect 32856 7588 32912 7644
rect 32912 7588 32916 7644
rect 32852 7584 32916 7588
rect 37612 7644 37676 7648
rect 37612 7588 37616 7644
rect 37616 7588 37672 7644
rect 37672 7588 37676 7644
rect 37612 7584 37676 7588
rect 37692 7644 37756 7648
rect 37692 7588 37696 7644
rect 37696 7588 37752 7644
rect 37752 7588 37756 7644
rect 37692 7584 37756 7588
rect 37772 7644 37836 7648
rect 37772 7588 37776 7644
rect 37776 7588 37832 7644
rect 37832 7588 37836 7644
rect 37772 7584 37836 7588
rect 37852 7644 37916 7648
rect 37852 7588 37856 7644
rect 37856 7588 37912 7644
rect 37912 7588 37916 7644
rect 37852 7584 37916 7588
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 6952 7100 7016 7104
rect 6952 7044 6956 7100
rect 6956 7044 7012 7100
rect 7012 7044 7016 7100
rect 6952 7040 7016 7044
rect 7032 7100 7096 7104
rect 7032 7044 7036 7100
rect 7036 7044 7092 7100
rect 7092 7044 7096 7100
rect 7032 7040 7096 7044
rect 7112 7100 7176 7104
rect 7112 7044 7116 7100
rect 7116 7044 7172 7100
rect 7172 7044 7176 7100
rect 7112 7040 7176 7044
rect 7192 7100 7256 7104
rect 7192 7044 7196 7100
rect 7196 7044 7252 7100
rect 7252 7044 7256 7100
rect 7192 7040 7256 7044
rect 11952 7100 12016 7104
rect 11952 7044 11956 7100
rect 11956 7044 12012 7100
rect 12012 7044 12016 7100
rect 11952 7040 12016 7044
rect 12032 7100 12096 7104
rect 12032 7044 12036 7100
rect 12036 7044 12092 7100
rect 12092 7044 12096 7100
rect 12032 7040 12096 7044
rect 12112 7100 12176 7104
rect 12112 7044 12116 7100
rect 12116 7044 12172 7100
rect 12172 7044 12176 7100
rect 12112 7040 12176 7044
rect 12192 7100 12256 7104
rect 12192 7044 12196 7100
rect 12196 7044 12252 7100
rect 12252 7044 12256 7100
rect 12192 7040 12256 7044
rect 16952 7100 17016 7104
rect 16952 7044 16956 7100
rect 16956 7044 17012 7100
rect 17012 7044 17016 7100
rect 16952 7040 17016 7044
rect 17032 7100 17096 7104
rect 17032 7044 17036 7100
rect 17036 7044 17092 7100
rect 17092 7044 17096 7100
rect 17032 7040 17096 7044
rect 17112 7100 17176 7104
rect 17112 7044 17116 7100
rect 17116 7044 17172 7100
rect 17172 7044 17176 7100
rect 17112 7040 17176 7044
rect 17192 7100 17256 7104
rect 17192 7044 17196 7100
rect 17196 7044 17252 7100
rect 17252 7044 17256 7100
rect 17192 7040 17256 7044
rect 21952 7100 22016 7104
rect 21952 7044 21956 7100
rect 21956 7044 22012 7100
rect 22012 7044 22016 7100
rect 21952 7040 22016 7044
rect 22032 7100 22096 7104
rect 22032 7044 22036 7100
rect 22036 7044 22092 7100
rect 22092 7044 22096 7100
rect 22032 7040 22096 7044
rect 22112 7100 22176 7104
rect 22112 7044 22116 7100
rect 22116 7044 22172 7100
rect 22172 7044 22176 7100
rect 22112 7040 22176 7044
rect 22192 7100 22256 7104
rect 22192 7044 22196 7100
rect 22196 7044 22252 7100
rect 22252 7044 22256 7100
rect 22192 7040 22256 7044
rect 26952 7100 27016 7104
rect 26952 7044 26956 7100
rect 26956 7044 27012 7100
rect 27012 7044 27016 7100
rect 26952 7040 27016 7044
rect 27032 7100 27096 7104
rect 27032 7044 27036 7100
rect 27036 7044 27092 7100
rect 27092 7044 27096 7100
rect 27032 7040 27096 7044
rect 27112 7100 27176 7104
rect 27112 7044 27116 7100
rect 27116 7044 27172 7100
rect 27172 7044 27176 7100
rect 27112 7040 27176 7044
rect 27192 7100 27256 7104
rect 27192 7044 27196 7100
rect 27196 7044 27252 7100
rect 27252 7044 27256 7100
rect 27192 7040 27256 7044
rect 31952 7100 32016 7104
rect 31952 7044 31956 7100
rect 31956 7044 32012 7100
rect 32012 7044 32016 7100
rect 31952 7040 32016 7044
rect 32032 7100 32096 7104
rect 32032 7044 32036 7100
rect 32036 7044 32092 7100
rect 32092 7044 32096 7100
rect 32032 7040 32096 7044
rect 32112 7100 32176 7104
rect 32112 7044 32116 7100
rect 32116 7044 32172 7100
rect 32172 7044 32176 7100
rect 32112 7040 32176 7044
rect 32192 7100 32256 7104
rect 32192 7044 32196 7100
rect 32196 7044 32252 7100
rect 32252 7044 32256 7100
rect 32192 7040 32256 7044
rect 36952 7100 37016 7104
rect 36952 7044 36956 7100
rect 36956 7044 37012 7100
rect 37012 7044 37016 7100
rect 36952 7040 37016 7044
rect 37032 7100 37096 7104
rect 37032 7044 37036 7100
rect 37036 7044 37092 7100
rect 37092 7044 37096 7100
rect 37032 7040 37096 7044
rect 37112 7100 37176 7104
rect 37112 7044 37116 7100
rect 37116 7044 37172 7100
rect 37172 7044 37176 7100
rect 37112 7040 37176 7044
rect 37192 7100 37256 7104
rect 37192 7044 37196 7100
rect 37196 7044 37252 7100
rect 37252 7044 37256 7100
rect 37192 7040 37256 7044
rect 2612 6556 2676 6560
rect 2612 6500 2616 6556
rect 2616 6500 2672 6556
rect 2672 6500 2676 6556
rect 2612 6496 2676 6500
rect 2692 6556 2756 6560
rect 2692 6500 2696 6556
rect 2696 6500 2752 6556
rect 2752 6500 2756 6556
rect 2692 6496 2756 6500
rect 2772 6556 2836 6560
rect 2772 6500 2776 6556
rect 2776 6500 2832 6556
rect 2832 6500 2836 6556
rect 2772 6496 2836 6500
rect 2852 6556 2916 6560
rect 2852 6500 2856 6556
rect 2856 6500 2912 6556
rect 2912 6500 2916 6556
rect 2852 6496 2916 6500
rect 7612 6556 7676 6560
rect 7612 6500 7616 6556
rect 7616 6500 7672 6556
rect 7672 6500 7676 6556
rect 7612 6496 7676 6500
rect 7692 6556 7756 6560
rect 7692 6500 7696 6556
rect 7696 6500 7752 6556
rect 7752 6500 7756 6556
rect 7692 6496 7756 6500
rect 7772 6556 7836 6560
rect 7772 6500 7776 6556
rect 7776 6500 7832 6556
rect 7832 6500 7836 6556
rect 7772 6496 7836 6500
rect 7852 6556 7916 6560
rect 7852 6500 7856 6556
rect 7856 6500 7912 6556
rect 7912 6500 7916 6556
rect 7852 6496 7916 6500
rect 12612 6556 12676 6560
rect 12612 6500 12616 6556
rect 12616 6500 12672 6556
rect 12672 6500 12676 6556
rect 12612 6496 12676 6500
rect 12692 6556 12756 6560
rect 12692 6500 12696 6556
rect 12696 6500 12752 6556
rect 12752 6500 12756 6556
rect 12692 6496 12756 6500
rect 12772 6556 12836 6560
rect 12772 6500 12776 6556
rect 12776 6500 12832 6556
rect 12832 6500 12836 6556
rect 12772 6496 12836 6500
rect 12852 6556 12916 6560
rect 12852 6500 12856 6556
rect 12856 6500 12912 6556
rect 12912 6500 12916 6556
rect 12852 6496 12916 6500
rect 17612 6556 17676 6560
rect 17612 6500 17616 6556
rect 17616 6500 17672 6556
rect 17672 6500 17676 6556
rect 17612 6496 17676 6500
rect 17692 6556 17756 6560
rect 17692 6500 17696 6556
rect 17696 6500 17752 6556
rect 17752 6500 17756 6556
rect 17692 6496 17756 6500
rect 17772 6556 17836 6560
rect 17772 6500 17776 6556
rect 17776 6500 17832 6556
rect 17832 6500 17836 6556
rect 17772 6496 17836 6500
rect 17852 6556 17916 6560
rect 17852 6500 17856 6556
rect 17856 6500 17912 6556
rect 17912 6500 17916 6556
rect 17852 6496 17916 6500
rect 22612 6556 22676 6560
rect 22612 6500 22616 6556
rect 22616 6500 22672 6556
rect 22672 6500 22676 6556
rect 22612 6496 22676 6500
rect 22692 6556 22756 6560
rect 22692 6500 22696 6556
rect 22696 6500 22752 6556
rect 22752 6500 22756 6556
rect 22692 6496 22756 6500
rect 22772 6556 22836 6560
rect 22772 6500 22776 6556
rect 22776 6500 22832 6556
rect 22832 6500 22836 6556
rect 22772 6496 22836 6500
rect 22852 6556 22916 6560
rect 22852 6500 22856 6556
rect 22856 6500 22912 6556
rect 22912 6500 22916 6556
rect 22852 6496 22916 6500
rect 27612 6556 27676 6560
rect 27612 6500 27616 6556
rect 27616 6500 27672 6556
rect 27672 6500 27676 6556
rect 27612 6496 27676 6500
rect 27692 6556 27756 6560
rect 27692 6500 27696 6556
rect 27696 6500 27752 6556
rect 27752 6500 27756 6556
rect 27692 6496 27756 6500
rect 27772 6556 27836 6560
rect 27772 6500 27776 6556
rect 27776 6500 27832 6556
rect 27832 6500 27836 6556
rect 27772 6496 27836 6500
rect 27852 6556 27916 6560
rect 27852 6500 27856 6556
rect 27856 6500 27912 6556
rect 27912 6500 27916 6556
rect 27852 6496 27916 6500
rect 32612 6556 32676 6560
rect 32612 6500 32616 6556
rect 32616 6500 32672 6556
rect 32672 6500 32676 6556
rect 32612 6496 32676 6500
rect 32692 6556 32756 6560
rect 32692 6500 32696 6556
rect 32696 6500 32752 6556
rect 32752 6500 32756 6556
rect 32692 6496 32756 6500
rect 32772 6556 32836 6560
rect 32772 6500 32776 6556
rect 32776 6500 32832 6556
rect 32832 6500 32836 6556
rect 32772 6496 32836 6500
rect 32852 6556 32916 6560
rect 32852 6500 32856 6556
rect 32856 6500 32912 6556
rect 32912 6500 32916 6556
rect 32852 6496 32916 6500
rect 37612 6556 37676 6560
rect 37612 6500 37616 6556
rect 37616 6500 37672 6556
rect 37672 6500 37676 6556
rect 37612 6496 37676 6500
rect 37692 6556 37756 6560
rect 37692 6500 37696 6556
rect 37696 6500 37752 6556
rect 37752 6500 37756 6556
rect 37692 6496 37756 6500
rect 37772 6556 37836 6560
rect 37772 6500 37776 6556
rect 37776 6500 37832 6556
rect 37832 6500 37836 6556
rect 37772 6496 37836 6500
rect 37852 6556 37916 6560
rect 37852 6500 37856 6556
rect 37856 6500 37912 6556
rect 37912 6500 37916 6556
rect 37852 6496 37916 6500
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 6952 6012 7016 6016
rect 6952 5956 6956 6012
rect 6956 5956 7012 6012
rect 7012 5956 7016 6012
rect 6952 5952 7016 5956
rect 7032 6012 7096 6016
rect 7032 5956 7036 6012
rect 7036 5956 7092 6012
rect 7092 5956 7096 6012
rect 7032 5952 7096 5956
rect 7112 6012 7176 6016
rect 7112 5956 7116 6012
rect 7116 5956 7172 6012
rect 7172 5956 7176 6012
rect 7112 5952 7176 5956
rect 7192 6012 7256 6016
rect 7192 5956 7196 6012
rect 7196 5956 7252 6012
rect 7252 5956 7256 6012
rect 7192 5952 7256 5956
rect 11952 6012 12016 6016
rect 11952 5956 11956 6012
rect 11956 5956 12012 6012
rect 12012 5956 12016 6012
rect 11952 5952 12016 5956
rect 12032 6012 12096 6016
rect 12032 5956 12036 6012
rect 12036 5956 12092 6012
rect 12092 5956 12096 6012
rect 12032 5952 12096 5956
rect 12112 6012 12176 6016
rect 12112 5956 12116 6012
rect 12116 5956 12172 6012
rect 12172 5956 12176 6012
rect 12112 5952 12176 5956
rect 12192 6012 12256 6016
rect 12192 5956 12196 6012
rect 12196 5956 12252 6012
rect 12252 5956 12256 6012
rect 12192 5952 12256 5956
rect 16952 6012 17016 6016
rect 16952 5956 16956 6012
rect 16956 5956 17012 6012
rect 17012 5956 17016 6012
rect 16952 5952 17016 5956
rect 17032 6012 17096 6016
rect 17032 5956 17036 6012
rect 17036 5956 17092 6012
rect 17092 5956 17096 6012
rect 17032 5952 17096 5956
rect 17112 6012 17176 6016
rect 17112 5956 17116 6012
rect 17116 5956 17172 6012
rect 17172 5956 17176 6012
rect 17112 5952 17176 5956
rect 17192 6012 17256 6016
rect 17192 5956 17196 6012
rect 17196 5956 17252 6012
rect 17252 5956 17256 6012
rect 17192 5952 17256 5956
rect 21952 6012 22016 6016
rect 21952 5956 21956 6012
rect 21956 5956 22012 6012
rect 22012 5956 22016 6012
rect 21952 5952 22016 5956
rect 22032 6012 22096 6016
rect 22032 5956 22036 6012
rect 22036 5956 22092 6012
rect 22092 5956 22096 6012
rect 22032 5952 22096 5956
rect 22112 6012 22176 6016
rect 22112 5956 22116 6012
rect 22116 5956 22172 6012
rect 22172 5956 22176 6012
rect 22112 5952 22176 5956
rect 22192 6012 22256 6016
rect 22192 5956 22196 6012
rect 22196 5956 22252 6012
rect 22252 5956 22256 6012
rect 22192 5952 22256 5956
rect 26952 6012 27016 6016
rect 26952 5956 26956 6012
rect 26956 5956 27012 6012
rect 27012 5956 27016 6012
rect 26952 5952 27016 5956
rect 27032 6012 27096 6016
rect 27032 5956 27036 6012
rect 27036 5956 27092 6012
rect 27092 5956 27096 6012
rect 27032 5952 27096 5956
rect 27112 6012 27176 6016
rect 27112 5956 27116 6012
rect 27116 5956 27172 6012
rect 27172 5956 27176 6012
rect 27112 5952 27176 5956
rect 27192 6012 27256 6016
rect 27192 5956 27196 6012
rect 27196 5956 27252 6012
rect 27252 5956 27256 6012
rect 27192 5952 27256 5956
rect 31952 6012 32016 6016
rect 31952 5956 31956 6012
rect 31956 5956 32012 6012
rect 32012 5956 32016 6012
rect 31952 5952 32016 5956
rect 32032 6012 32096 6016
rect 32032 5956 32036 6012
rect 32036 5956 32092 6012
rect 32092 5956 32096 6012
rect 32032 5952 32096 5956
rect 32112 6012 32176 6016
rect 32112 5956 32116 6012
rect 32116 5956 32172 6012
rect 32172 5956 32176 6012
rect 32112 5952 32176 5956
rect 32192 6012 32256 6016
rect 32192 5956 32196 6012
rect 32196 5956 32252 6012
rect 32252 5956 32256 6012
rect 32192 5952 32256 5956
rect 36952 6012 37016 6016
rect 36952 5956 36956 6012
rect 36956 5956 37012 6012
rect 37012 5956 37016 6012
rect 36952 5952 37016 5956
rect 37032 6012 37096 6016
rect 37032 5956 37036 6012
rect 37036 5956 37092 6012
rect 37092 5956 37096 6012
rect 37032 5952 37096 5956
rect 37112 6012 37176 6016
rect 37112 5956 37116 6012
rect 37116 5956 37172 6012
rect 37172 5956 37176 6012
rect 37112 5952 37176 5956
rect 37192 6012 37256 6016
rect 37192 5956 37196 6012
rect 37196 5956 37252 6012
rect 37252 5956 37256 6012
rect 37192 5952 37256 5956
rect 2612 5468 2676 5472
rect 2612 5412 2616 5468
rect 2616 5412 2672 5468
rect 2672 5412 2676 5468
rect 2612 5408 2676 5412
rect 2692 5468 2756 5472
rect 2692 5412 2696 5468
rect 2696 5412 2752 5468
rect 2752 5412 2756 5468
rect 2692 5408 2756 5412
rect 2772 5468 2836 5472
rect 2772 5412 2776 5468
rect 2776 5412 2832 5468
rect 2832 5412 2836 5468
rect 2772 5408 2836 5412
rect 2852 5468 2916 5472
rect 2852 5412 2856 5468
rect 2856 5412 2912 5468
rect 2912 5412 2916 5468
rect 2852 5408 2916 5412
rect 7612 5468 7676 5472
rect 7612 5412 7616 5468
rect 7616 5412 7672 5468
rect 7672 5412 7676 5468
rect 7612 5408 7676 5412
rect 7692 5468 7756 5472
rect 7692 5412 7696 5468
rect 7696 5412 7752 5468
rect 7752 5412 7756 5468
rect 7692 5408 7756 5412
rect 7772 5468 7836 5472
rect 7772 5412 7776 5468
rect 7776 5412 7832 5468
rect 7832 5412 7836 5468
rect 7772 5408 7836 5412
rect 7852 5468 7916 5472
rect 7852 5412 7856 5468
rect 7856 5412 7912 5468
rect 7912 5412 7916 5468
rect 7852 5408 7916 5412
rect 12612 5468 12676 5472
rect 12612 5412 12616 5468
rect 12616 5412 12672 5468
rect 12672 5412 12676 5468
rect 12612 5408 12676 5412
rect 12692 5468 12756 5472
rect 12692 5412 12696 5468
rect 12696 5412 12752 5468
rect 12752 5412 12756 5468
rect 12692 5408 12756 5412
rect 12772 5468 12836 5472
rect 12772 5412 12776 5468
rect 12776 5412 12832 5468
rect 12832 5412 12836 5468
rect 12772 5408 12836 5412
rect 12852 5468 12916 5472
rect 12852 5412 12856 5468
rect 12856 5412 12912 5468
rect 12912 5412 12916 5468
rect 12852 5408 12916 5412
rect 17612 5468 17676 5472
rect 17612 5412 17616 5468
rect 17616 5412 17672 5468
rect 17672 5412 17676 5468
rect 17612 5408 17676 5412
rect 17692 5468 17756 5472
rect 17692 5412 17696 5468
rect 17696 5412 17752 5468
rect 17752 5412 17756 5468
rect 17692 5408 17756 5412
rect 17772 5468 17836 5472
rect 17772 5412 17776 5468
rect 17776 5412 17832 5468
rect 17832 5412 17836 5468
rect 17772 5408 17836 5412
rect 17852 5468 17916 5472
rect 17852 5412 17856 5468
rect 17856 5412 17912 5468
rect 17912 5412 17916 5468
rect 17852 5408 17916 5412
rect 22612 5468 22676 5472
rect 22612 5412 22616 5468
rect 22616 5412 22672 5468
rect 22672 5412 22676 5468
rect 22612 5408 22676 5412
rect 22692 5468 22756 5472
rect 22692 5412 22696 5468
rect 22696 5412 22752 5468
rect 22752 5412 22756 5468
rect 22692 5408 22756 5412
rect 22772 5468 22836 5472
rect 22772 5412 22776 5468
rect 22776 5412 22832 5468
rect 22832 5412 22836 5468
rect 22772 5408 22836 5412
rect 22852 5468 22916 5472
rect 22852 5412 22856 5468
rect 22856 5412 22912 5468
rect 22912 5412 22916 5468
rect 22852 5408 22916 5412
rect 27612 5468 27676 5472
rect 27612 5412 27616 5468
rect 27616 5412 27672 5468
rect 27672 5412 27676 5468
rect 27612 5408 27676 5412
rect 27692 5468 27756 5472
rect 27692 5412 27696 5468
rect 27696 5412 27752 5468
rect 27752 5412 27756 5468
rect 27692 5408 27756 5412
rect 27772 5468 27836 5472
rect 27772 5412 27776 5468
rect 27776 5412 27832 5468
rect 27832 5412 27836 5468
rect 27772 5408 27836 5412
rect 27852 5468 27916 5472
rect 27852 5412 27856 5468
rect 27856 5412 27912 5468
rect 27912 5412 27916 5468
rect 27852 5408 27916 5412
rect 32612 5468 32676 5472
rect 32612 5412 32616 5468
rect 32616 5412 32672 5468
rect 32672 5412 32676 5468
rect 32612 5408 32676 5412
rect 32692 5468 32756 5472
rect 32692 5412 32696 5468
rect 32696 5412 32752 5468
rect 32752 5412 32756 5468
rect 32692 5408 32756 5412
rect 32772 5468 32836 5472
rect 32772 5412 32776 5468
rect 32776 5412 32832 5468
rect 32832 5412 32836 5468
rect 32772 5408 32836 5412
rect 32852 5468 32916 5472
rect 32852 5412 32856 5468
rect 32856 5412 32912 5468
rect 32912 5412 32916 5468
rect 32852 5408 32916 5412
rect 37612 5468 37676 5472
rect 37612 5412 37616 5468
rect 37616 5412 37672 5468
rect 37672 5412 37676 5468
rect 37612 5408 37676 5412
rect 37692 5468 37756 5472
rect 37692 5412 37696 5468
rect 37696 5412 37752 5468
rect 37752 5412 37756 5468
rect 37692 5408 37756 5412
rect 37772 5468 37836 5472
rect 37772 5412 37776 5468
rect 37776 5412 37832 5468
rect 37832 5412 37836 5468
rect 37772 5408 37836 5412
rect 37852 5468 37916 5472
rect 37852 5412 37856 5468
rect 37856 5412 37912 5468
rect 37912 5412 37916 5468
rect 37852 5408 37916 5412
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 6952 4924 7016 4928
rect 6952 4868 6956 4924
rect 6956 4868 7012 4924
rect 7012 4868 7016 4924
rect 6952 4864 7016 4868
rect 7032 4924 7096 4928
rect 7032 4868 7036 4924
rect 7036 4868 7092 4924
rect 7092 4868 7096 4924
rect 7032 4864 7096 4868
rect 7112 4924 7176 4928
rect 7112 4868 7116 4924
rect 7116 4868 7172 4924
rect 7172 4868 7176 4924
rect 7112 4864 7176 4868
rect 7192 4924 7256 4928
rect 7192 4868 7196 4924
rect 7196 4868 7252 4924
rect 7252 4868 7256 4924
rect 7192 4864 7256 4868
rect 11952 4924 12016 4928
rect 11952 4868 11956 4924
rect 11956 4868 12012 4924
rect 12012 4868 12016 4924
rect 11952 4864 12016 4868
rect 12032 4924 12096 4928
rect 12032 4868 12036 4924
rect 12036 4868 12092 4924
rect 12092 4868 12096 4924
rect 12032 4864 12096 4868
rect 12112 4924 12176 4928
rect 12112 4868 12116 4924
rect 12116 4868 12172 4924
rect 12172 4868 12176 4924
rect 12112 4864 12176 4868
rect 12192 4924 12256 4928
rect 12192 4868 12196 4924
rect 12196 4868 12252 4924
rect 12252 4868 12256 4924
rect 12192 4864 12256 4868
rect 16952 4924 17016 4928
rect 16952 4868 16956 4924
rect 16956 4868 17012 4924
rect 17012 4868 17016 4924
rect 16952 4864 17016 4868
rect 17032 4924 17096 4928
rect 17032 4868 17036 4924
rect 17036 4868 17092 4924
rect 17092 4868 17096 4924
rect 17032 4864 17096 4868
rect 17112 4924 17176 4928
rect 17112 4868 17116 4924
rect 17116 4868 17172 4924
rect 17172 4868 17176 4924
rect 17112 4864 17176 4868
rect 17192 4924 17256 4928
rect 17192 4868 17196 4924
rect 17196 4868 17252 4924
rect 17252 4868 17256 4924
rect 17192 4864 17256 4868
rect 21952 4924 22016 4928
rect 21952 4868 21956 4924
rect 21956 4868 22012 4924
rect 22012 4868 22016 4924
rect 21952 4864 22016 4868
rect 22032 4924 22096 4928
rect 22032 4868 22036 4924
rect 22036 4868 22092 4924
rect 22092 4868 22096 4924
rect 22032 4864 22096 4868
rect 22112 4924 22176 4928
rect 22112 4868 22116 4924
rect 22116 4868 22172 4924
rect 22172 4868 22176 4924
rect 22112 4864 22176 4868
rect 22192 4924 22256 4928
rect 22192 4868 22196 4924
rect 22196 4868 22252 4924
rect 22252 4868 22256 4924
rect 22192 4864 22256 4868
rect 26952 4924 27016 4928
rect 26952 4868 26956 4924
rect 26956 4868 27012 4924
rect 27012 4868 27016 4924
rect 26952 4864 27016 4868
rect 27032 4924 27096 4928
rect 27032 4868 27036 4924
rect 27036 4868 27092 4924
rect 27092 4868 27096 4924
rect 27032 4864 27096 4868
rect 27112 4924 27176 4928
rect 27112 4868 27116 4924
rect 27116 4868 27172 4924
rect 27172 4868 27176 4924
rect 27112 4864 27176 4868
rect 27192 4924 27256 4928
rect 27192 4868 27196 4924
rect 27196 4868 27252 4924
rect 27252 4868 27256 4924
rect 27192 4864 27256 4868
rect 31952 4924 32016 4928
rect 31952 4868 31956 4924
rect 31956 4868 32012 4924
rect 32012 4868 32016 4924
rect 31952 4864 32016 4868
rect 32032 4924 32096 4928
rect 32032 4868 32036 4924
rect 32036 4868 32092 4924
rect 32092 4868 32096 4924
rect 32032 4864 32096 4868
rect 32112 4924 32176 4928
rect 32112 4868 32116 4924
rect 32116 4868 32172 4924
rect 32172 4868 32176 4924
rect 32112 4864 32176 4868
rect 32192 4924 32256 4928
rect 32192 4868 32196 4924
rect 32196 4868 32252 4924
rect 32252 4868 32256 4924
rect 32192 4864 32256 4868
rect 36952 4924 37016 4928
rect 36952 4868 36956 4924
rect 36956 4868 37012 4924
rect 37012 4868 37016 4924
rect 36952 4864 37016 4868
rect 37032 4924 37096 4928
rect 37032 4868 37036 4924
rect 37036 4868 37092 4924
rect 37092 4868 37096 4924
rect 37032 4864 37096 4868
rect 37112 4924 37176 4928
rect 37112 4868 37116 4924
rect 37116 4868 37172 4924
rect 37172 4868 37176 4924
rect 37112 4864 37176 4868
rect 37192 4924 37256 4928
rect 37192 4868 37196 4924
rect 37196 4868 37252 4924
rect 37252 4868 37256 4924
rect 37192 4864 37256 4868
rect 2612 4380 2676 4384
rect 2612 4324 2616 4380
rect 2616 4324 2672 4380
rect 2672 4324 2676 4380
rect 2612 4320 2676 4324
rect 2692 4380 2756 4384
rect 2692 4324 2696 4380
rect 2696 4324 2752 4380
rect 2752 4324 2756 4380
rect 2692 4320 2756 4324
rect 2772 4380 2836 4384
rect 2772 4324 2776 4380
rect 2776 4324 2832 4380
rect 2832 4324 2836 4380
rect 2772 4320 2836 4324
rect 2852 4380 2916 4384
rect 2852 4324 2856 4380
rect 2856 4324 2912 4380
rect 2912 4324 2916 4380
rect 2852 4320 2916 4324
rect 7612 4380 7676 4384
rect 7612 4324 7616 4380
rect 7616 4324 7672 4380
rect 7672 4324 7676 4380
rect 7612 4320 7676 4324
rect 7692 4380 7756 4384
rect 7692 4324 7696 4380
rect 7696 4324 7752 4380
rect 7752 4324 7756 4380
rect 7692 4320 7756 4324
rect 7772 4380 7836 4384
rect 7772 4324 7776 4380
rect 7776 4324 7832 4380
rect 7832 4324 7836 4380
rect 7772 4320 7836 4324
rect 7852 4380 7916 4384
rect 7852 4324 7856 4380
rect 7856 4324 7912 4380
rect 7912 4324 7916 4380
rect 7852 4320 7916 4324
rect 12612 4380 12676 4384
rect 12612 4324 12616 4380
rect 12616 4324 12672 4380
rect 12672 4324 12676 4380
rect 12612 4320 12676 4324
rect 12692 4380 12756 4384
rect 12692 4324 12696 4380
rect 12696 4324 12752 4380
rect 12752 4324 12756 4380
rect 12692 4320 12756 4324
rect 12772 4380 12836 4384
rect 12772 4324 12776 4380
rect 12776 4324 12832 4380
rect 12832 4324 12836 4380
rect 12772 4320 12836 4324
rect 12852 4380 12916 4384
rect 12852 4324 12856 4380
rect 12856 4324 12912 4380
rect 12912 4324 12916 4380
rect 12852 4320 12916 4324
rect 17612 4380 17676 4384
rect 17612 4324 17616 4380
rect 17616 4324 17672 4380
rect 17672 4324 17676 4380
rect 17612 4320 17676 4324
rect 17692 4380 17756 4384
rect 17692 4324 17696 4380
rect 17696 4324 17752 4380
rect 17752 4324 17756 4380
rect 17692 4320 17756 4324
rect 17772 4380 17836 4384
rect 17772 4324 17776 4380
rect 17776 4324 17832 4380
rect 17832 4324 17836 4380
rect 17772 4320 17836 4324
rect 17852 4380 17916 4384
rect 17852 4324 17856 4380
rect 17856 4324 17912 4380
rect 17912 4324 17916 4380
rect 17852 4320 17916 4324
rect 22612 4380 22676 4384
rect 22612 4324 22616 4380
rect 22616 4324 22672 4380
rect 22672 4324 22676 4380
rect 22612 4320 22676 4324
rect 22692 4380 22756 4384
rect 22692 4324 22696 4380
rect 22696 4324 22752 4380
rect 22752 4324 22756 4380
rect 22692 4320 22756 4324
rect 22772 4380 22836 4384
rect 22772 4324 22776 4380
rect 22776 4324 22832 4380
rect 22832 4324 22836 4380
rect 22772 4320 22836 4324
rect 22852 4380 22916 4384
rect 22852 4324 22856 4380
rect 22856 4324 22912 4380
rect 22912 4324 22916 4380
rect 22852 4320 22916 4324
rect 27612 4380 27676 4384
rect 27612 4324 27616 4380
rect 27616 4324 27672 4380
rect 27672 4324 27676 4380
rect 27612 4320 27676 4324
rect 27692 4380 27756 4384
rect 27692 4324 27696 4380
rect 27696 4324 27752 4380
rect 27752 4324 27756 4380
rect 27692 4320 27756 4324
rect 27772 4380 27836 4384
rect 27772 4324 27776 4380
rect 27776 4324 27832 4380
rect 27832 4324 27836 4380
rect 27772 4320 27836 4324
rect 27852 4380 27916 4384
rect 27852 4324 27856 4380
rect 27856 4324 27912 4380
rect 27912 4324 27916 4380
rect 27852 4320 27916 4324
rect 32612 4380 32676 4384
rect 32612 4324 32616 4380
rect 32616 4324 32672 4380
rect 32672 4324 32676 4380
rect 32612 4320 32676 4324
rect 32692 4380 32756 4384
rect 32692 4324 32696 4380
rect 32696 4324 32752 4380
rect 32752 4324 32756 4380
rect 32692 4320 32756 4324
rect 32772 4380 32836 4384
rect 32772 4324 32776 4380
rect 32776 4324 32832 4380
rect 32832 4324 32836 4380
rect 32772 4320 32836 4324
rect 32852 4380 32916 4384
rect 32852 4324 32856 4380
rect 32856 4324 32912 4380
rect 32912 4324 32916 4380
rect 32852 4320 32916 4324
rect 37612 4380 37676 4384
rect 37612 4324 37616 4380
rect 37616 4324 37672 4380
rect 37672 4324 37676 4380
rect 37612 4320 37676 4324
rect 37692 4380 37756 4384
rect 37692 4324 37696 4380
rect 37696 4324 37752 4380
rect 37752 4324 37756 4380
rect 37692 4320 37756 4324
rect 37772 4380 37836 4384
rect 37772 4324 37776 4380
rect 37776 4324 37832 4380
rect 37832 4324 37836 4380
rect 37772 4320 37836 4324
rect 37852 4380 37916 4384
rect 37852 4324 37856 4380
rect 37856 4324 37912 4380
rect 37912 4324 37916 4380
rect 37852 4320 37916 4324
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 6952 3836 7016 3840
rect 6952 3780 6956 3836
rect 6956 3780 7012 3836
rect 7012 3780 7016 3836
rect 6952 3776 7016 3780
rect 7032 3836 7096 3840
rect 7032 3780 7036 3836
rect 7036 3780 7092 3836
rect 7092 3780 7096 3836
rect 7032 3776 7096 3780
rect 7112 3836 7176 3840
rect 7112 3780 7116 3836
rect 7116 3780 7172 3836
rect 7172 3780 7176 3836
rect 7112 3776 7176 3780
rect 7192 3836 7256 3840
rect 7192 3780 7196 3836
rect 7196 3780 7252 3836
rect 7252 3780 7256 3836
rect 7192 3776 7256 3780
rect 11952 3836 12016 3840
rect 11952 3780 11956 3836
rect 11956 3780 12012 3836
rect 12012 3780 12016 3836
rect 11952 3776 12016 3780
rect 12032 3836 12096 3840
rect 12032 3780 12036 3836
rect 12036 3780 12092 3836
rect 12092 3780 12096 3836
rect 12032 3776 12096 3780
rect 12112 3836 12176 3840
rect 12112 3780 12116 3836
rect 12116 3780 12172 3836
rect 12172 3780 12176 3836
rect 12112 3776 12176 3780
rect 12192 3836 12256 3840
rect 12192 3780 12196 3836
rect 12196 3780 12252 3836
rect 12252 3780 12256 3836
rect 12192 3776 12256 3780
rect 16952 3836 17016 3840
rect 16952 3780 16956 3836
rect 16956 3780 17012 3836
rect 17012 3780 17016 3836
rect 16952 3776 17016 3780
rect 17032 3836 17096 3840
rect 17032 3780 17036 3836
rect 17036 3780 17092 3836
rect 17092 3780 17096 3836
rect 17032 3776 17096 3780
rect 17112 3836 17176 3840
rect 17112 3780 17116 3836
rect 17116 3780 17172 3836
rect 17172 3780 17176 3836
rect 17112 3776 17176 3780
rect 17192 3836 17256 3840
rect 17192 3780 17196 3836
rect 17196 3780 17252 3836
rect 17252 3780 17256 3836
rect 17192 3776 17256 3780
rect 21952 3836 22016 3840
rect 21952 3780 21956 3836
rect 21956 3780 22012 3836
rect 22012 3780 22016 3836
rect 21952 3776 22016 3780
rect 22032 3836 22096 3840
rect 22032 3780 22036 3836
rect 22036 3780 22092 3836
rect 22092 3780 22096 3836
rect 22032 3776 22096 3780
rect 22112 3836 22176 3840
rect 22112 3780 22116 3836
rect 22116 3780 22172 3836
rect 22172 3780 22176 3836
rect 22112 3776 22176 3780
rect 22192 3836 22256 3840
rect 22192 3780 22196 3836
rect 22196 3780 22252 3836
rect 22252 3780 22256 3836
rect 22192 3776 22256 3780
rect 26952 3836 27016 3840
rect 26952 3780 26956 3836
rect 26956 3780 27012 3836
rect 27012 3780 27016 3836
rect 26952 3776 27016 3780
rect 27032 3836 27096 3840
rect 27032 3780 27036 3836
rect 27036 3780 27092 3836
rect 27092 3780 27096 3836
rect 27032 3776 27096 3780
rect 27112 3836 27176 3840
rect 27112 3780 27116 3836
rect 27116 3780 27172 3836
rect 27172 3780 27176 3836
rect 27112 3776 27176 3780
rect 27192 3836 27256 3840
rect 27192 3780 27196 3836
rect 27196 3780 27252 3836
rect 27252 3780 27256 3836
rect 27192 3776 27256 3780
rect 31952 3836 32016 3840
rect 31952 3780 31956 3836
rect 31956 3780 32012 3836
rect 32012 3780 32016 3836
rect 31952 3776 32016 3780
rect 32032 3836 32096 3840
rect 32032 3780 32036 3836
rect 32036 3780 32092 3836
rect 32092 3780 32096 3836
rect 32032 3776 32096 3780
rect 32112 3836 32176 3840
rect 32112 3780 32116 3836
rect 32116 3780 32172 3836
rect 32172 3780 32176 3836
rect 32112 3776 32176 3780
rect 32192 3836 32256 3840
rect 32192 3780 32196 3836
rect 32196 3780 32252 3836
rect 32252 3780 32256 3836
rect 32192 3776 32256 3780
rect 36952 3836 37016 3840
rect 36952 3780 36956 3836
rect 36956 3780 37012 3836
rect 37012 3780 37016 3836
rect 36952 3776 37016 3780
rect 37032 3836 37096 3840
rect 37032 3780 37036 3836
rect 37036 3780 37092 3836
rect 37092 3780 37096 3836
rect 37032 3776 37096 3780
rect 37112 3836 37176 3840
rect 37112 3780 37116 3836
rect 37116 3780 37172 3836
rect 37172 3780 37176 3836
rect 37112 3776 37176 3780
rect 37192 3836 37256 3840
rect 37192 3780 37196 3836
rect 37196 3780 37252 3836
rect 37252 3780 37256 3836
rect 37192 3776 37256 3780
rect 2612 3292 2676 3296
rect 2612 3236 2616 3292
rect 2616 3236 2672 3292
rect 2672 3236 2676 3292
rect 2612 3232 2676 3236
rect 2692 3292 2756 3296
rect 2692 3236 2696 3292
rect 2696 3236 2752 3292
rect 2752 3236 2756 3292
rect 2692 3232 2756 3236
rect 2772 3292 2836 3296
rect 2772 3236 2776 3292
rect 2776 3236 2832 3292
rect 2832 3236 2836 3292
rect 2772 3232 2836 3236
rect 2852 3292 2916 3296
rect 2852 3236 2856 3292
rect 2856 3236 2912 3292
rect 2912 3236 2916 3292
rect 2852 3232 2916 3236
rect 7612 3292 7676 3296
rect 7612 3236 7616 3292
rect 7616 3236 7672 3292
rect 7672 3236 7676 3292
rect 7612 3232 7676 3236
rect 7692 3292 7756 3296
rect 7692 3236 7696 3292
rect 7696 3236 7752 3292
rect 7752 3236 7756 3292
rect 7692 3232 7756 3236
rect 7772 3292 7836 3296
rect 7772 3236 7776 3292
rect 7776 3236 7832 3292
rect 7832 3236 7836 3292
rect 7772 3232 7836 3236
rect 7852 3292 7916 3296
rect 7852 3236 7856 3292
rect 7856 3236 7912 3292
rect 7912 3236 7916 3292
rect 7852 3232 7916 3236
rect 12612 3292 12676 3296
rect 12612 3236 12616 3292
rect 12616 3236 12672 3292
rect 12672 3236 12676 3292
rect 12612 3232 12676 3236
rect 12692 3292 12756 3296
rect 12692 3236 12696 3292
rect 12696 3236 12752 3292
rect 12752 3236 12756 3292
rect 12692 3232 12756 3236
rect 12772 3292 12836 3296
rect 12772 3236 12776 3292
rect 12776 3236 12832 3292
rect 12832 3236 12836 3292
rect 12772 3232 12836 3236
rect 12852 3292 12916 3296
rect 12852 3236 12856 3292
rect 12856 3236 12912 3292
rect 12912 3236 12916 3292
rect 12852 3232 12916 3236
rect 17612 3292 17676 3296
rect 17612 3236 17616 3292
rect 17616 3236 17672 3292
rect 17672 3236 17676 3292
rect 17612 3232 17676 3236
rect 17692 3292 17756 3296
rect 17692 3236 17696 3292
rect 17696 3236 17752 3292
rect 17752 3236 17756 3292
rect 17692 3232 17756 3236
rect 17772 3292 17836 3296
rect 17772 3236 17776 3292
rect 17776 3236 17832 3292
rect 17832 3236 17836 3292
rect 17772 3232 17836 3236
rect 17852 3292 17916 3296
rect 17852 3236 17856 3292
rect 17856 3236 17912 3292
rect 17912 3236 17916 3292
rect 17852 3232 17916 3236
rect 22612 3292 22676 3296
rect 22612 3236 22616 3292
rect 22616 3236 22672 3292
rect 22672 3236 22676 3292
rect 22612 3232 22676 3236
rect 22692 3292 22756 3296
rect 22692 3236 22696 3292
rect 22696 3236 22752 3292
rect 22752 3236 22756 3292
rect 22692 3232 22756 3236
rect 22772 3292 22836 3296
rect 22772 3236 22776 3292
rect 22776 3236 22832 3292
rect 22832 3236 22836 3292
rect 22772 3232 22836 3236
rect 22852 3292 22916 3296
rect 22852 3236 22856 3292
rect 22856 3236 22912 3292
rect 22912 3236 22916 3292
rect 22852 3232 22916 3236
rect 27612 3292 27676 3296
rect 27612 3236 27616 3292
rect 27616 3236 27672 3292
rect 27672 3236 27676 3292
rect 27612 3232 27676 3236
rect 27692 3292 27756 3296
rect 27692 3236 27696 3292
rect 27696 3236 27752 3292
rect 27752 3236 27756 3292
rect 27692 3232 27756 3236
rect 27772 3292 27836 3296
rect 27772 3236 27776 3292
rect 27776 3236 27832 3292
rect 27832 3236 27836 3292
rect 27772 3232 27836 3236
rect 27852 3292 27916 3296
rect 27852 3236 27856 3292
rect 27856 3236 27912 3292
rect 27912 3236 27916 3292
rect 27852 3232 27916 3236
rect 32612 3292 32676 3296
rect 32612 3236 32616 3292
rect 32616 3236 32672 3292
rect 32672 3236 32676 3292
rect 32612 3232 32676 3236
rect 32692 3292 32756 3296
rect 32692 3236 32696 3292
rect 32696 3236 32752 3292
rect 32752 3236 32756 3292
rect 32692 3232 32756 3236
rect 32772 3292 32836 3296
rect 32772 3236 32776 3292
rect 32776 3236 32832 3292
rect 32832 3236 32836 3292
rect 32772 3232 32836 3236
rect 32852 3292 32916 3296
rect 32852 3236 32856 3292
rect 32856 3236 32912 3292
rect 32912 3236 32916 3292
rect 32852 3232 32916 3236
rect 37612 3292 37676 3296
rect 37612 3236 37616 3292
rect 37616 3236 37672 3292
rect 37672 3236 37676 3292
rect 37612 3232 37676 3236
rect 37692 3292 37756 3296
rect 37692 3236 37696 3292
rect 37696 3236 37752 3292
rect 37752 3236 37756 3292
rect 37692 3232 37756 3236
rect 37772 3292 37836 3296
rect 37772 3236 37776 3292
rect 37776 3236 37832 3292
rect 37832 3236 37836 3292
rect 37772 3232 37836 3236
rect 37852 3292 37916 3296
rect 37852 3236 37856 3292
rect 37856 3236 37912 3292
rect 37912 3236 37916 3292
rect 37852 3232 37916 3236
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 6952 2748 7016 2752
rect 6952 2692 6956 2748
rect 6956 2692 7012 2748
rect 7012 2692 7016 2748
rect 6952 2688 7016 2692
rect 7032 2748 7096 2752
rect 7032 2692 7036 2748
rect 7036 2692 7092 2748
rect 7092 2692 7096 2748
rect 7032 2688 7096 2692
rect 7112 2748 7176 2752
rect 7112 2692 7116 2748
rect 7116 2692 7172 2748
rect 7172 2692 7176 2748
rect 7112 2688 7176 2692
rect 7192 2748 7256 2752
rect 7192 2692 7196 2748
rect 7196 2692 7252 2748
rect 7252 2692 7256 2748
rect 7192 2688 7256 2692
rect 11952 2748 12016 2752
rect 11952 2692 11956 2748
rect 11956 2692 12012 2748
rect 12012 2692 12016 2748
rect 11952 2688 12016 2692
rect 12032 2748 12096 2752
rect 12032 2692 12036 2748
rect 12036 2692 12092 2748
rect 12092 2692 12096 2748
rect 12032 2688 12096 2692
rect 12112 2748 12176 2752
rect 12112 2692 12116 2748
rect 12116 2692 12172 2748
rect 12172 2692 12176 2748
rect 12112 2688 12176 2692
rect 12192 2748 12256 2752
rect 12192 2692 12196 2748
rect 12196 2692 12252 2748
rect 12252 2692 12256 2748
rect 12192 2688 12256 2692
rect 16952 2748 17016 2752
rect 16952 2692 16956 2748
rect 16956 2692 17012 2748
rect 17012 2692 17016 2748
rect 16952 2688 17016 2692
rect 17032 2748 17096 2752
rect 17032 2692 17036 2748
rect 17036 2692 17092 2748
rect 17092 2692 17096 2748
rect 17032 2688 17096 2692
rect 17112 2748 17176 2752
rect 17112 2692 17116 2748
rect 17116 2692 17172 2748
rect 17172 2692 17176 2748
rect 17112 2688 17176 2692
rect 17192 2748 17256 2752
rect 17192 2692 17196 2748
rect 17196 2692 17252 2748
rect 17252 2692 17256 2748
rect 17192 2688 17256 2692
rect 21952 2748 22016 2752
rect 21952 2692 21956 2748
rect 21956 2692 22012 2748
rect 22012 2692 22016 2748
rect 21952 2688 22016 2692
rect 22032 2748 22096 2752
rect 22032 2692 22036 2748
rect 22036 2692 22092 2748
rect 22092 2692 22096 2748
rect 22032 2688 22096 2692
rect 22112 2748 22176 2752
rect 22112 2692 22116 2748
rect 22116 2692 22172 2748
rect 22172 2692 22176 2748
rect 22112 2688 22176 2692
rect 22192 2748 22256 2752
rect 22192 2692 22196 2748
rect 22196 2692 22252 2748
rect 22252 2692 22256 2748
rect 22192 2688 22256 2692
rect 26952 2748 27016 2752
rect 26952 2692 26956 2748
rect 26956 2692 27012 2748
rect 27012 2692 27016 2748
rect 26952 2688 27016 2692
rect 27032 2748 27096 2752
rect 27032 2692 27036 2748
rect 27036 2692 27092 2748
rect 27092 2692 27096 2748
rect 27032 2688 27096 2692
rect 27112 2748 27176 2752
rect 27112 2692 27116 2748
rect 27116 2692 27172 2748
rect 27172 2692 27176 2748
rect 27112 2688 27176 2692
rect 27192 2748 27256 2752
rect 27192 2692 27196 2748
rect 27196 2692 27252 2748
rect 27252 2692 27256 2748
rect 27192 2688 27256 2692
rect 31952 2748 32016 2752
rect 31952 2692 31956 2748
rect 31956 2692 32012 2748
rect 32012 2692 32016 2748
rect 31952 2688 32016 2692
rect 32032 2748 32096 2752
rect 32032 2692 32036 2748
rect 32036 2692 32092 2748
rect 32092 2692 32096 2748
rect 32032 2688 32096 2692
rect 32112 2748 32176 2752
rect 32112 2692 32116 2748
rect 32116 2692 32172 2748
rect 32172 2692 32176 2748
rect 32112 2688 32176 2692
rect 32192 2748 32256 2752
rect 32192 2692 32196 2748
rect 32196 2692 32252 2748
rect 32252 2692 32256 2748
rect 32192 2688 32256 2692
rect 36952 2748 37016 2752
rect 36952 2692 36956 2748
rect 36956 2692 37012 2748
rect 37012 2692 37016 2748
rect 36952 2688 37016 2692
rect 37032 2748 37096 2752
rect 37032 2692 37036 2748
rect 37036 2692 37092 2748
rect 37092 2692 37096 2748
rect 37032 2688 37096 2692
rect 37112 2748 37176 2752
rect 37112 2692 37116 2748
rect 37116 2692 37172 2748
rect 37172 2692 37176 2748
rect 37112 2688 37176 2692
rect 37192 2748 37256 2752
rect 37192 2692 37196 2748
rect 37196 2692 37252 2748
rect 37252 2692 37256 2748
rect 37192 2688 37256 2692
rect 2612 2204 2676 2208
rect 2612 2148 2616 2204
rect 2616 2148 2672 2204
rect 2672 2148 2676 2204
rect 2612 2144 2676 2148
rect 2692 2204 2756 2208
rect 2692 2148 2696 2204
rect 2696 2148 2752 2204
rect 2752 2148 2756 2204
rect 2692 2144 2756 2148
rect 2772 2204 2836 2208
rect 2772 2148 2776 2204
rect 2776 2148 2832 2204
rect 2832 2148 2836 2204
rect 2772 2144 2836 2148
rect 2852 2204 2916 2208
rect 2852 2148 2856 2204
rect 2856 2148 2912 2204
rect 2912 2148 2916 2204
rect 2852 2144 2916 2148
rect 7612 2204 7676 2208
rect 7612 2148 7616 2204
rect 7616 2148 7672 2204
rect 7672 2148 7676 2204
rect 7612 2144 7676 2148
rect 7692 2204 7756 2208
rect 7692 2148 7696 2204
rect 7696 2148 7752 2204
rect 7752 2148 7756 2204
rect 7692 2144 7756 2148
rect 7772 2204 7836 2208
rect 7772 2148 7776 2204
rect 7776 2148 7832 2204
rect 7832 2148 7836 2204
rect 7772 2144 7836 2148
rect 7852 2204 7916 2208
rect 7852 2148 7856 2204
rect 7856 2148 7912 2204
rect 7912 2148 7916 2204
rect 7852 2144 7916 2148
rect 12612 2204 12676 2208
rect 12612 2148 12616 2204
rect 12616 2148 12672 2204
rect 12672 2148 12676 2204
rect 12612 2144 12676 2148
rect 12692 2204 12756 2208
rect 12692 2148 12696 2204
rect 12696 2148 12752 2204
rect 12752 2148 12756 2204
rect 12692 2144 12756 2148
rect 12772 2204 12836 2208
rect 12772 2148 12776 2204
rect 12776 2148 12832 2204
rect 12832 2148 12836 2204
rect 12772 2144 12836 2148
rect 12852 2204 12916 2208
rect 12852 2148 12856 2204
rect 12856 2148 12912 2204
rect 12912 2148 12916 2204
rect 12852 2144 12916 2148
rect 17612 2204 17676 2208
rect 17612 2148 17616 2204
rect 17616 2148 17672 2204
rect 17672 2148 17676 2204
rect 17612 2144 17676 2148
rect 17692 2204 17756 2208
rect 17692 2148 17696 2204
rect 17696 2148 17752 2204
rect 17752 2148 17756 2204
rect 17692 2144 17756 2148
rect 17772 2204 17836 2208
rect 17772 2148 17776 2204
rect 17776 2148 17832 2204
rect 17832 2148 17836 2204
rect 17772 2144 17836 2148
rect 17852 2204 17916 2208
rect 17852 2148 17856 2204
rect 17856 2148 17912 2204
rect 17912 2148 17916 2204
rect 17852 2144 17916 2148
rect 22612 2204 22676 2208
rect 22612 2148 22616 2204
rect 22616 2148 22672 2204
rect 22672 2148 22676 2204
rect 22612 2144 22676 2148
rect 22692 2204 22756 2208
rect 22692 2148 22696 2204
rect 22696 2148 22752 2204
rect 22752 2148 22756 2204
rect 22692 2144 22756 2148
rect 22772 2204 22836 2208
rect 22772 2148 22776 2204
rect 22776 2148 22832 2204
rect 22832 2148 22836 2204
rect 22772 2144 22836 2148
rect 22852 2204 22916 2208
rect 22852 2148 22856 2204
rect 22856 2148 22912 2204
rect 22912 2148 22916 2204
rect 22852 2144 22916 2148
rect 27612 2204 27676 2208
rect 27612 2148 27616 2204
rect 27616 2148 27672 2204
rect 27672 2148 27676 2204
rect 27612 2144 27676 2148
rect 27692 2204 27756 2208
rect 27692 2148 27696 2204
rect 27696 2148 27752 2204
rect 27752 2148 27756 2204
rect 27692 2144 27756 2148
rect 27772 2204 27836 2208
rect 27772 2148 27776 2204
rect 27776 2148 27832 2204
rect 27832 2148 27836 2204
rect 27772 2144 27836 2148
rect 27852 2204 27916 2208
rect 27852 2148 27856 2204
rect 27856 2148 27912 2204
rect 27912 2148 27916 2204
rect 27852 2144 27916 2148
rect 32612 2204 32676 2208
rect 32612 2148 32616 2204
rect 32616 2148 32672 2204
rect 32672 2148 32676 2204
rect 32612 2144 32676 2148
rect 32692 2204 32756 2208
rect 32692 2148 32696 2204
rect 32696 2148 32752 2204
rect 32752 2148 32756 2204
rect 32692 2144 32756 2148
rect 32772 2204 32836 2208
rect 32772 2148 32776 2204
rect 32776 2148 32832 2204
rect 32832 2148 32836 2204
rect 32772 2144 32836 2148
rect 32852 2204 32916 2208
rect 32852 2148 32856 2204
rect 32856 2148 32912 2204
rect 32912 2148 32916 2204
rect 32852 2144 32916 2148
rect 37612 2204 37676 2208
rect 37612 2148 37616 2204
rect 37616 2148 37672 2204
rect 37672 2148 37676 2204
rect 37612 2144 37676 2148
rect 37692 2204 37756 2208
rect 37692 2148 37696 2204
rect 37696 2148 37752 2204
rect 37752 2148 37756 2204
rect 37692 2144 37756 2148
rect 37772 2204 37836 2208
rect 37772 2148 37776 2204
rect 37776 2148 37832 2204
rect 37832 2148 37836 2204
rect 37772 2144 37836 2148
rect 37852 2204 37916 2208
rect 37852 2148 37856 2204
rect 37856 2148 37912 2204
rect 37912 2148 37916 2204
rect 37852 2144 37916 2148
<< metal4 >>
rect 1944 69120 2264 69680
rect 1944 69056 1952 69120
rect 2016 69056 2032 69120
rect 2096 69056 2112 69120
rect 2176 69056 2192 69120
rect 2256 69056 2264 69120
rect 1944 68294 2264 69056
rect 1944 68058 1986 68294
rect 2222 68058 2264 68294
rect 1944 68032 2264 68058
rect 1944 67968 1952 68032
rect 2016 67968 2032 68032
rect 2096 67968 2112 68032
rect 2176 67968 2192 68032
rect 2256 67968 2264 68032
rect 1944 66944 2264 67968
rect 1944 66880 1952 66944
rect 2016 66880 2032 66944
rect 2096 66880 2112 66944
rect 2176 66880 2192 66944
rect 2256 66880 2264 66944
rect 1944 65856 2264 66880
rect 1944 65792 1952 65856
rect 2016 65792 2032 65856
rect 2096 65792 2112 65856
rect 2176 65792 2192 65856
rect 2256 65792 2264 65856
rect 1944 64768 2264 65792
rect 1944 64704 1952 64768
rect 2016 64704 2032 64768
rect 2096 64704 2112 64768
rect 2176 64704 2192 64768
rect 2256 64704 2264 64768
rect 1944 63680 2264 64704
rect 1944 63616 1952 63680
rect 2016 63616 2032 63680
rect 2096 63616 2112 63680
rect 2176 63616 2192 63680
rect 2256 63616 2264 63680
rect 1944 63294 2264 63616
rect 1944 63058 1986 63294
rect 2222 63058 2264 63294
rect 1944 62592 2264 63058
rect 1944 62528 1952 62592
rect 2016 62528 2032 62592
rect 2096 62528 2112 62592
rect 2176 62528 2192 62592
rect 2256 62528 2264 62592
rect 1944 61504 2264 62528
rect 1944 61440 1952 61504
rect 2016 61440 2032 61504
rect 2096 61440 2112 61504
rect 2176 61440 2192 61504
rect 2256 61440 2264 61504
rect 1944 60416 2264 61440
rect 1944 60352 1952 60416
rect 2016 60352 2032 60416
rect 2096 60352 2112 60416
rect 2176 60352 2192 60416
rect 2256 60352 2264 60416
rect 1944 59328 2264 60352
rect 1944 59264 1952 59328
rect 2016 59264 2032 59328
rect 2096 59264 2112 59328
rect 2176 59264 2192 59328
rect 2256 59264 2264 59328
rect 1944 58294 2264 59264
rect 1944 58240 1986 58294
rect 2222 58240 2264 58294
rect 1944 58176 1952 58240
rect 2256 58176 2264 58240
rect 1944 58058 1986 58176
rect 2222 58058 2264 58176
rect 1944 57152 2264 58058
rect 1944 57088 1952 57152
rect 2016 57088 2032 57152
rect 2096 57088 2112 57152
rect 2176 57088 2192 57152
rect 2256 57088 2264 57152
rect 1944 56064 2264 57088
rect 1944 56000 1952 56064
rect 2016 56000 2032 56064
rect 2096 56000 2112 56064
rect 2176 56000 2192 56064
rect 2256 56000 2264 56064
rect 1944 54976 2264 56000
rect 1944 54912 1952 54976
rect 2016 54912 2032 54976
rect 2096 54912 2112 54976
rect 2176 54912 2192 54976
rect 2256 54912 2264 54976
rect 1944 53888 2264 54912
rect 1944 53824 1952 53888
rect 2016 53824 2032 53888
rect 2096 53824 2112 53888
rect 2176 53824 2192 53888
rect 2256 53824 2264 53888
rect 1944 53294 2264 53824
rect 1944 53058 1986 53294
rect 2222 53058 2264 53294
rect 1944 52800 2264 53058
rect 1944 52736 1952 52800
rect 2016 52736 2032 52800
rect 2096 52736 2112 52800
rect 2176 52736 2192 52800
rect 2256 52736 2264 52800
rect 1944 51712 2264 52736
rect 1944 51648 1952 51712
rect 2016 51648 2032 51712
rect 2096 51648 2112 51712
rect 2176 51648 2192 51712
rect 2256 51648 2264 51712
rect 1944 50624 2264 51648
rect 1944 50560 1952 50624
rect 2016 50560 2032 50624
rect 2096 50560 2112 50624
rect 2176 50560 2192 50624
rect 2256 50560 2264 50624
rect 1944 49536 2264 50560
rect 1944 49472 1952 49536
rect 2016 49472 2032 49536
rect 2096 49472 2112 49536
rect 2176 49472 2192 49536
rect 2256 49472 2264 49536
rect 1944 48448 2264 49472
rect 1944 48384 1952 48448
rect 2016 48384 2032 48448
rect 2096 48384 2112 48448
rect 2176 48384 2192 48448
rect 2256 48384 2264 48448
rect 1944 48294 2264 48384
rect 1944 48058 1986 48294
rect 2222 48058 2264 48294
rect 1944 47360 2264 48058
rect 1944 47296 1952 47360
rect 2016 47296 2032 47360
rect 2096 47296 2112 47360
rect 2176 47296 2192 47360
rect 2256 47296 2264 47360
rect 1944 46272 2264 47296
rect 1944 46208 1952 46272
rect 2016 46208 2032 46272
rect 2096 46208 2112 46272
rect 2176 46208 2192 46272
rect 2256 46208 2264 46272
rect 1944 45184 2264 46208
rect 1944 45120 1952 45184
rect 2016 45120 2032 45184
rect 2096 45120 2112 45184
rect 2176 45120 2192 45184
rect 2256 45120 2264 45184
rect 1944 44096 2264 45120
rect 1944 44032 1952 44096
rect 2016 44032 2032 44096
rect 2096 44032 2112 44096
rect 2176 44032 2192 44096
rect 2256 44032 2264 44096
rect 1944 43294 2264 44032
rect 1944 43058 1986 43294
rect 2222 43058 2264 43294
rect 1944 43008 2264 43058
rect 1944 42944 1952 43008
rect 2016 42944 2032 43008
rect 2096 42944 2112 43008
rect 2176 42944 2192 43008
rect 2256 42944 2264 43008
rect 1944 41920 2264 42944
rect 1944 41856 1952 41920
rect 2016 41856 2032 41920
rect 2096 41856 2112 41920
rect 2176 41856 2192 41920
rect 2256 41856 2264 41920
rect 1944 40832 2264 41856
rect 1944 40768 1952 40832
rect 2016 40768 2032 40832
rect 2096 40768 2112 40832
rect 2176 40768 2192 40832
rect 2256 40768 2264 40832
rect 1944 39744 2264 40768
rect 1944 39680 1952 39744
rect 2016 39680 2032 39744
rect 2096 39680 2112 39744
rect 2176 39680 2192 39744
rect 2256 39680 2264 39744
rect 1944 38656 2264 39680
rect 1944 38592 1952 38656
rect 2016 38592 2032 38656
rect 2096 38592 2112 38656
rect 2176 38592 2192 38656
rect 2256 38592 2264 38656
rect 1944 38294 2264 38592
rect 1944 38058 1986 38294
rect 2222 38058 2264 38294
rect 1944 37568 2264 38058
rect 1944 37504 1952 37568
rect 2016 37504 2032 37568
rect 2096 37504 2112 37568
rect 2176 37504 2192 37568
rect 2256 37504 2264 37568
rect 1944 36480 2264 37504
rect 1944 36416 1952 36480
rect 2016 36416 2032 36480
rect 2096 36416 2112 36480
rect 2176 36416 2192 36480
rect 2256 36416 2264 36480
rect 1944 35392 2264 36416
rect 1944 35328 1952 35392
rect 2016 35328 2032 35392
rect 2096 35328 2112 35392
rect 2176 35328 2192 35392
rect 2256 35328 2264 35392
rect 1944 34304 2264 35328
rect 1944 34240 1952 34304
rect 2016 34240 2032 34304
rect 2096 34240 2112 34304
rect 2176 34240 2192 34304
rect 2256 34240 2264 34304
rect 1944 33294 2264 34240
rect 1944 33216 1986 33294
rect 2222 33216 2264 33294
rect 1944 33152 1952 33216
rect 2256 33152 2264 33216
rect 1944 33058 1986 33152
rect 2222 33058 2264 33152
rect 1944 32128 2264 33058
rect 1944 32064 1952 32128
rect 2016 32064 2032 32128
rect 2096 32064 2112 32128
rect 2176 32064 2192 32128
rect 2256 32064 2264 32128
rect 1944 31040 2264 32064
rect 1944 30976 1952 31040
rect 2016 30976 2032 31040
rect 2096 30976 2112 31040
rect 2176 30976 2192 31040
rect 2256 30976 2264 31040
rect 1944 29952 2264 30976
rect 1944 29888 1952 29952
rect 2016 29888 2032 29952
rect 2096 29888 2112 29952
rect 2176 29888 2192 29952
rect 2256 29888 2264 29952
rect 1944 28864 2264 29888
rect 1944 28800 1952 28864
rect 2016 28800 2032 28864
rect 2096 28800 2112 28864
rect 2176 28800 2192 28864
rect 2256 28800 2264 28864
rect 1944 28294 2264 28800
rect 1944 28058 1986 28294
rect 2222 28058 2264 28294
rect 1944 27776 2264 28058
rect 1944 27712 1952 27776
rect 2016 27712 2032 27776
rect 2096 27712 2112 27776
rect 2176 27712 2192 27776
rect 2256 27712 2264 27776
rect 1944 26688 2264 27712
rect 1944 26624 1952 26688
rect 2016 26624 2032 26688
rect 2096 26624 2112 26688
rect 2176 26624 2192 26688
rect 2256 26624 2264 26688
rect 1944 25600 2264 26624
rect 1944 25536 1952 25600
rect 2016 25536 2032 25600
rect 2096 25536 2112 25600
rect 2176 25536 2192 25600
rect 2256 25536 2264 25600
rect 1944 24512 2264 25536
rect 1944 24448 1952 24512
rect 2016 24448 2032 24512
rect 2096 24448 2112 24512
rect 2176 24448 2192 24512
rect 2256 24448 2264 24512
rect 1944 23424 2264 24448
rect 1944 23360 1952 23424
rect 2016 23360 2032 23424
rect 2096 23360 2112 23424
rect 2176 23360 2192 23424
rect 2256 23360 2264 23424
rect 1944 23294 2264 23360
rect 1944 23058 1986 23294
rect 2222 23058 2264 23294
rect 1944 22336 2264 23058
rect 1944 22272 1952 22336
rect 2016 22272 2032 22336
rect 2096 22272 2112 22336
rect 2176 22272 2192 22336
rect 2256 22272 2264 22336
rect 1944 21248 2264 22272
rect 1944 21184 1952 21248
rect 2016 21184 2032 21248
rect 2096 21184 2112 21248
rect 2176 21184 2192 21248
rect 2256 21184 2264 21248
rect 1944 20160 2264 21184
rect 1944 20096 1952 20160
rect 2016 20096 2032 20160
rect 2096 20096 2112 20160
rect 2176 20096 2192 20160
rect 2256 20096 2264 20160
rect 1944 19072 2264 20096
rect 1944 19008 1952 19072
rect 2016 19008 2032 19072
rect 2096 19008 2112 19072
rect 2176 19008 2192 19072
rect 2256 19008 2264 19072
rect 1944 18294 2264 19008
rect 1944 18058 1986 18294
rect 2222 18058 2264 18294
rect 1944 17984 2264 18058
rect 1944 17920 1952 17984
rect 2016 17920 2032 17984
rect 2096 17920 2112 17984
rect 2176 17920 2192 17984
rect 2256 17920 2264 17984
rect 1944 16896 2264 17920
rect 1944 16832 1952 16896
rect 2016 16832 2032 16896
rect 2096 16832 2112 16896
rect 2176 16832 2192 16896
rect 2256 16832 2264 16896
rect 1944 15808 2264 16832
rect 1944 15744 1952 15808
rect 2016 15744 2032 15808
rect 2096 15744 2112 15808
rect 2176 15744 2192 15808
rect 2256 15744 2264 15808
rect 1944 14720 2264 15744
rect 1944 14656 1952 14720
rect 2016 14656 2032 14720
rect 2096 14656 2112 14720
rect 2176 14656 2192 14720
rect 2256 14656 2264 14720
rect 1944 13632 2264 14656
rect 1944 13568 1952 13632
rect 2016 13568 2032 13632
rect 2096 13568 2112 13632
rect 2176 13568 2192 13632
rect 2256 13568 2264 13632
rect 1944 13294 2264 13568
rect 1944 13058 1986 13294
rect 2222 13058 2264 13294
rect 1944 12544 2264 13058
rect 1944 12480 1952 12544
rect 2016 12480 2032 12544
rect 2096 12480 2112 12544
rect 2176 12480 2192 12544
rect 2256 12480 2264 12544
rect 1944 11456 2264 12480
rect 1944 11392 1952 11456
rect 2016 11392 2032 11456
rect 2096 11392 2112 11456
rect 2176 11392 2192 11456
rect 2256 11392 2264 11456
rect 1944 10368 2264 11392
rect 1944 10304 1952 10368
rect 2016 10304 2032 10368
rect 2096 10304 2112 10368
rect 2176 10304 2192 10368
rect 2256 10304 2264 10368
rect 1944 9280 2264 10304
rect 1944 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2264 9280
rect 1944 8294 2264 9216
rect 1944 8192 1986 8294
rect 2222 8192 2264 8294
rect 1944 8128 1952 8192
rect 2256 8128 2264 8192
rect 1944 8058 1986 8128
rect 2222 8058 2264 8128
rect 1944 7104 2264 8058
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 3294 2264 3776
rect 1944 3058 1986 3294
rect 2222 3058 2264 3294
rect 1944 2752 2264 3058
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 2128 2264 2688
rect 2604 69664 2924 69680
rect 2604 69600 2612 69664
rect 2676 69600 2692 69664
rect 2756 69600 2772 69664
rect 2836 69600 2852 69664
rect 2916 69600 2924 69664
rect 2604 68954 2924 69600
rect 2604 68718 2646 68954
rect 2882 68718 2924 68954
rect 2604 68576 2924 68718
rect 2604 68512 2612 68576
rect 2676 68512 2692 68576
rect 2756 68512 2772 68576
rect 2836 68512 2852 68576
rect 2916 68512 2924 68576
rect 2604 67488 2924 68512
rect 2604 67424 2612 67488
rect 2676 67424 2692 67488
rect 2756 67424 2772 67488
rect 2836 67424 2852 67488
rect 2916 67424 2924 67488
rect 2604 66400 2924 67424
rect 2604 66336 2612 66400
rect 2676 66336 2692 66400
rect 2756 66336 2772 66400
rect 2836 66336 2852 66400
rect 2916 66336 2924 66400
rect 2604 65312 2924 66336
rect 2604 65248 2612 65312
rect 2676 65248 2692 65312
rect 2756 65248 2772 65312
rect 2836 65248 2852 65312
rect 2916 65248 2924 65312
rect 2604 64224 2924 65248
rect 2604 64160 2612 64224
rect 2676 64160 2692 64224
rect 2756 64160 2772 64224
rect 2836 64160 2852 64224
rect 2916 64160 2924 64224
rect 2604 63954 2924 64160
rect 2604 63718 2646 63954
rect 2882 63718 2924 63954
rect 2604 63136 2924 63718
rect 2604 63072 2612 63136
rect 2676 63072 2692 63136
rect 2756 63072 2772 63136
rect 2836 63072 2852 63136
rect 2916 63072 2924 63136
rect 2604 62048 2924 63072
rect 2604 61984 2612 62048
rect 2676 61984 2692 62048
rect 2756 61984 2772 62048
rect 2836 61984 2852 62048
rect 2916 61984 2924 62048
rect 2604 60960 2924 61984
rect 2604 60896 2612 60960
rect 2676 60896 2692 60960
rect 2756 60896 2772 60960
rect 2836 60896 2852 60960
rect 2916 60896 2924 60960
rect 2604 59872 2924 60896
rect 2604 59808 2612 59872
rect 2676 59808 2692 59872
rect 2756 59808 2772 59872
rect 2836 59808 2852 59872
rect 2916 59808 2924 59872
rect 2604 58954 2924 59808
rect 2604 58784 2646 58954
rect 2882 58784 2924 58954
rect 2604 58720 2612 58784
rect 2916 58720 2924 58784
rect 2604 58718 2646 58720
rect 2882 58718 2924 58720
rect 2604 57696 2924 58718
rect 2604 57632 2612 57696
rect 2676 57632 2692 57696
rect 2756 57632 2772 57696
rect 2836 57632 2852 57696
rect 2916 57632 2924 57696
rect 2604 56608 2924 57632
rect 2604 56544 2612 56608
rect 2676 56544 2692 56608
rect 2756 56544 2772 56608
rect 2836 56544 2852 56608
rect 2916 56544 2924 56608
rect 2604 55520 2924 56544
rect 2604 55456 2612 55520
rect 2676 55456 2692 55520
rect 2756 55456 2772 55520
rect 2836 55456 2852 55520
rect 2916 55456 2924 55520
rect 2604 54432 2924 55456
rect 2604 54368 2612 54432
rect 2676 54368 2692 54432
rect 2756 54368 2772 54432
rect 2836 54368 2852 54432
rect 2916 54368 2924 54432
rect 2604 53954 2924 54368
rect 2604 53718 2646 53954
rect 2882 53718 2924 53954
rect 2604 53344 2924 53718
rect 2604 53280 2612 53344
rect 2676 53280 2692 53344
rect 2756 53280 2772 53344
rect 2836 53280 2852 53344
rect 2916 53280 2924 53344
rect 2604 52256 2924 53280
rect 2604 52192 2612 52256
rect 2676 52192 2692 52256
rect 2756 52192 2772 52256
rect 2836 52192 2852 52256
rect 2916 52192 2924 52256
rect 2604 51168 2924 52192
rect 2604 51104 2612 51168
rect 2676 51104 2692 51168
rect 2756 51104 2772 51168
rect 2836 51104 2852 51168
rect 2916 51104 2924 51168
rect 2604 50080 2924 51104
rect 2604 50016 2612 50080
rect 2676 50016 2692 50080
rect 2756 50016 2772 50080
rect 2836 50016 2852 50080
rect 2916 50016 2924 50080
rect 2604 48992 2924 50016
rect 2604 48928 2612 48992
rect 2676 48954 2692 48992
rect 2756 48954 2772 48992
rect 2836 48954 2852 48992
rect 2916 48928 2924 48992
rect 2604 48718 2646 48928
rect 2882 48718 2924 48928
rect 2604 47904 2924 48718
rect 2604 47840 2612 47904
rect 2676 47840 2692 47904
rect 2756 47840 2772 47904
rect 2836 47840 2852 47904
rect 2916 47840 2924 47904
rect 2604 46816 2924 47840
rect 2604 46752 2612 46816
rect 2676 46752 2692 46816
rect 2756 46752 2772 46816
rect 2836 46752 2852 46816
rect 2916 46752 2924 46816
rect 2604 45728 2924 46752
rect 2604 45664 2612 45728
rect 2676 45664 2692 45728
rect 2756 45664 2772 45728
rect 2836 45664 2852 45728
rect 2916 45664 2924 45728
rect 2604 44640 2924 45664
rect 2604 44576 2612 44640
rect 2676 44576 2692 44640
rect 2756 44576 2772 44640
rect 2836 44576 2852 44640
rect 2916 44576 2924 44640
rect 2604 43954 2924 44576
rect 2604 43718 2646 43954
rect 2882 43718 2924 43954
rect 2604 43552 2924 43718
rect 2604 43488 2612 43552
rect 2676 43488 2692 43552
rect 2756 43488 2772 43552
rect 2836 43488 2852 43552
rect 2916 43488 2924 43552
rect 2604 42464 2924 43488
rect 2604 42400 2612 42464
rect 2676 42400 2692 42464
rect 2756 42400 2772 42464
rect 2836 42400 2852 42464
rect 2916 42400 2924 42464
rect 2604 41376 2924 42400
rect 2604 41312 2612 41376
rect 2676 41312 2692 41376
rect 2756 41312 2772 41376
rect 2836 41312 2852 41376
rect 2916 41312 2924 41376
rect 2604 40288 2924 41312
rect 2604 40224 2612 40288
rect 2676 40224 2692 40288
rect 2756 40224 2772 40288
rect 2836 40224 2852 40288
rect 2916 40224 2924 40288
rect 2604 39200 2924 40224
rect 2604 39136 2612 39200
rect 2676 39136 2692 39200
rect 2756 39136 2772 39200
rect 2836 39136 2852 39200
rect 2916 39136 2924 39200
rect 2604 38954 2924 39136
rect 2604 38718 2646 38954
rect 2882 38718 2924 38954
rect 2604 38112 2924 38718
rect 2604 38048 2612 38112
rect 2676 38048 2692 38112
rect 2756 38048 2772 38112
rect 2836 38048 2852 38112
rect 2916 38048 2924 38112
rect 2604 37024 2924 38048
rect 2604 36960 2612 37024
rect 2676 36960 2692 37024
rect 2756 36960 2772 37024
rect 2836 36960 2852 37024
rect 2916 36960 2924 37024
rect 2604 35936 2924 36960
rect 2604 35872 2612 35936
rect 2676 35872 2692 35936
rect 2756 35872 2772 35936
rect 2836 35872 2852 35936
rect 2916 35872 2924 35936
rect 2604 34848 2924 35872
rect 2604 34784 2612 34848
rect 2676 34784 2692 34848
rect 2756 34784 2772 34848
rect 2836 34784 2852 34848
rect 2916 34784 2924 34848
rect 2604 33954 2924 34784
rect 2604 33760 2646 33954
rect 2882 33760 2924 33954
rect 2604 33696 2612 33760
rect 2676 33696 2692 33718
rect 2756 33696 2772 33718
rect 2836 33696 2852 33718
rect 2916 33696 2924 33760
rect 2604 32672 2924 33696
rect 2604 32608 2612 32672
rect 2676 32608 2692 32672
rect 2756 32608 2772 32672
rect 2836 32608 2852 32672
rect 2916 32608 2924 32672
rect 2604 31584 2924 32608
rect 2604 31520 2612 31584
rect 2676 31520 2692 31584
rect 2756 31520 2772 31584
rect 2836 31520 2852 31584
rect 2916 31520 2924 31584
rect 2604 30496 2924 31520
rect 2604 30432 2612 30496
rect 2676 30432 2692 30496
rect 2756 30432 2772 30496
rect 2836 30432 2852 30496
rect 2916 30432 2924 30496
rect 2604 29408 2924 30432
rect 2604 29344 2612 29408
rect 2676 29344 2692 29408
rect 2756 29344 2772 29408
rect 2836 29344 2852 29408
rect 2916 29344 2924 29408
rect 2604 28954 2924 29344
rect 2604 28718 2646 28954
rect 2882 28718 2924 28954
rect 2604 28320 2924 28718
rect 2604 28256 2612 28320
rect 2676 28256 2692 28320
rect 2756 28256 2772 28320
rect 2836 28256 2852 28320
rect 2916 28256 2924 28320
rect 2604 27232 2924 28256
rect 2604 27168 2612 27232
rect 2676 27168 2692 27232
rect 2756 27168 2772 27232
rect 2836 27168 2852 27232
rect 2916 27168 2924 27232
rect 2604 26144 2924 27168
rect 2604 26080 2612 26144
rect 2676 26080 2692 26144
rect 2756 26080 2772 26144
rect 2836 26080 2852 26144
rect 2916 26080 2924 26144
rect 2604 25056 2924 26080
rect 2604 24992 2612 25056
rect 2676 24992 2692 25056
rect 2756 24992 2772 25056
rect 2836 24992 2852 25056
rect 2916 24992 2924 25056
rect 2604 23968 2924 24992
rect 2604 23904 2612 23968
rect 2676 23954 2692 23968
rect 2756 23954 2772 23968
rect 2836 23954 2852 23968
rect 2916 23904 2924 23968
rect 2604 23718 2646 23904
rect 2882 23718 2924 23904
rect 2604 22880 2924 23718
rect 2604 22816 2612 22880
rect 2676 22816 2692 22880
rect 2756 22816 2772 22880
rect 2836 22816 2852 22880
rect 2916 22816 2924 22880
rect 2604 21792 2924 22816
rect 2604 21728 2612 21792
rect 2676 21728 2692 21792
rect 2756 21728 2772 21792
rect 2836 21728 2852 21792
rect 2916 21728 2924 21792
rect 2604 20704 2924 21728
rect 2604 20640 2612 20704
rect 2676 20640 2692 20704
rect 2756 20640 2772 20704
rect 2836 20640 2852 20704
rect 2916 20640 2924 20704
rect 2604 19616 2924 20640
rect 2604 19552 2612 19616
rect 2676 19552 2692 19616
rect 2756 19552 2772 19616
rect 2836 19552 2852 19616
rect 2916 19552 2924 19616
rect 2604 18954 2924 19552
rect 2604 18718 2646 18954
rect 2882 18718 2924 18954
rect 2604 18528 2924 18718
rect 2604 18464 2612 18528
rect 2676 18464 2692 18528
rect 2756 18464 2772 18528
rect 2836 18464 2852 18528
rect 2916 18464 2924 18528
rect 2604 17440 2924 18464
rect 2604 17376 2612 17440
rect 2676 17376 2692 17440
rect 2756 17376 2772 17440
rect 2836 17376 2852 17440
rect 2916 17376 2924 17440
rect 2604 16352 2924 17376
rect 2604 16288 2612 16352
rect 2676 16288 2692 16352
rect 2756 16288 2772 16352
rect 2836 16288 2852 16352
rect 2916 16288 2924 16352
rect 2604 15264 2924 16288
rect 2604 15200 2612 15264
rect 2676 15200 2692 15264
rect 2756 15200 2772 15264
rect 2836 15200 2852 15264
rect 2916 15200 2924 15264
rect 2604 14176 2924 15200
rect 2604 14112 2612 14176
rect 2676 14112 2692 14176
rect 2756 14112 2772 14176
rect 2836 14112 2852 14176
rect 2916 14112 2924 14176
rect 2604 13954 2924 14112
rect 2604 13718 2646 13954
rect 2882 13718 2924 13954
rect 2604 13088 2924 13718
rect 2604 13024 2612 13088
rect 2676 13024 2692 13088
rect 2756 13024 2772 13088
rect 2836 13024 2852 13088
rect 2916 13024 2924 13088
rect 2604 12000 2924 13024
rect 2604 11936 2612 12000
rect 2676 11936 2692 12000
rect 2756 11936 2772 12000
rect 2836 11936 2852 12000
rect 2916 11936 2924 12000
rect 2604 10912 2924 11936
rect 2604 10848 2612 10912
rect 2676 10848 2692 10912
rect 2756 10848 2772 10912
rect 2836 10848 2852 10912
rect 2916 10848 2924 10912
rect 2604 9824 2924 10848
rect 2604 9760 2612 9824
rect 2676 9760 2692 9824
rect 2756 9760 2772 9824
rect 2836 9760 2852 9824
rect 2916 9760 2924 9824
rect 2604 8954 2924 9760
rect 2604 8736 2646 8954
rect 2882 8736 2924 8954
rect 2604 8672 2612 8736
rect 2676 8672 2692 8718
rect 2756 8672 2772 8718
rect 2836 8672 2852 8718
rect 2916 8672 2924 8736
rect 2604 7648 2924 8672
rect 2604 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2924 7648
rect 2604 6560 2924 7584
rect 2604 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2924 6560
rect 2604 5472 2924 6496
rect 2604 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2924 5472
rect 2604 4384 2924 5408
rect 2604 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2924 4384
rect 2604 3954 2924 4320
rect 2604 3718 2646 3954
rect 2882 3718 2924 3954
rect 2604 3296 2924 3718
rect 2604 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2924 3296
rect 2604 2208 2924 3232
rect 2604 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2924 2208
rect 2604 2128 2924 2144
rect 6944 69120 7264 69680
rect 6944 69056 6952 69120
rect 7016 69056 7032 69120
rect 7096 69056 7112 69120
rect 7176 69056 7192 69120
rect 7256 69056 7264 69120
rect 6944 68294 7264 69056
rect 6944 68058 6986 68294
rect 7222 68058 7264 68294
rect 6944 68032 7264 68058
rect 6944 67968 6952 68032
rect 7016 67968 7032 68032
rect 7096 67968 7112 68032
rect 7176 67968 7192 68032
rect 7256 67968 7264 68032
rect 6944 66944 7264 67968
rect 6944 66880 6952 66944
rect 7016 66880 7032 66944
rect 7096 66880 7112 66944
rect 7176 66880 7192 66944
rect 7256 66880 7264 66944
rect 6944 65856 7264 66880
rect 6944 65792 6952 65856
rect 7016 65792 7032 65856
rect 7096 65792 7112 65856
rect 7176 65792 7192 65856
rect 7256 65792 7264 65856
rect 6944 64768 7264 65792
rect 6944 64704 6952 64768
rect 7016 64704 7032 64768
rect 7096 64704 7112 64768
rect 7176 64704 7192 64768
rect 7256 64704 7264 64768
rect 6944 63680 7264 64704
rect 6944 63616 6952 63680
rect 7016 63616 7032 63680
rect 7096 63616 7112 63680
rect 7176 63616 7192 63680
rect 7256 63616 7264 63680
rect 6944 63294 7264 63616
rect 6944 63058 6986 63294
rect 7222 63058 7264 63294
rect 6944 62592 7264 63058
rect 6944 62528 6952 62592
rect 7016 62528 7032 62592
rect 7096 62528 7112 62592
rect 7176 62528 7192 62592
rect 7256 62528 7264 62592
rect 6944 61504 7264 62528
rect 6944 61440 6952 61504
rect 7016 61440 7032 61504
rect 7096 61440 7112 61504
rect 7176 61440 7192 61504
rect 7256 61440 7264 61504
rect 6944 60416 7264 61440
rect 6944 60352 6952 60416
rect 7016 60352 7032 60416
rect 7096 60352 7112 60416
rect 7176 60352 7192 60416
rect 7256 60352 7264 60416
rect 6944 59328 7264 60352
rect 6944 59264 6952 59328
rect 7016 59264 7032 59328
rect 7096 59264 7112 59328
rect 7176 59264 7192 59328
rect 7256 59264 7264 59328
rect 6944 58294 7264 59264
rect 6944 58240 6986 58294
rect 7222 58240 7264 58294
rect 6944 58176 6952 58240
rect 7256 58176 7264 58240
rect 6944 58058 6986 58176
rect 7222 58058 7264 58176
rect 6944 57152 7264 58058
rect 6944 57088 6952 57152
rect 7016 57088 7032 57152
rect 7096 57088 7112 57152
rect 7176 57088 7192 57152
rect 7256 57088 7264 57152
rect 6944 56064 7264 57088
rect 6944 56000 6952 56064
rect 7016 56000 7032 56064
rect 7096 56000 7112 56064
rect 7176 56000 7192 56064
rect 7256 56000 7264 56064
rect 6944 54976 7264 56000
rect 6944 54912 6952 54976
rect 7016 54912 7032 54976
rect 7096 54912 7112 54976
rect 7176 54912 7192 54976
rect 7256 54912 7264 54976
rect 6944 53888 7264 54912
rect 6944 53824 6952 53888
rect 7016 53824 7032 53888
rect 7096 53824 7112 53888
rect 7176 53824 7192 53888
rect 7256 53824 7264 53888
rect 6944 53294 7264 53824
rect 6944 53058 6986 53294
rect 7222 53058 7264 53294
rect 6944 52800 7264 53058
rect 6944 52736 6952 52800
rect 7016 52736 7032 52800
rect 7096 52736 7112 52800
rect 7176 52736 7192 52800
rect 7256 52736 7264 52800
rect 6944 51712 7264 52736
rect 6944 51648 6952 51712
rect 7016 51648 7032 51712
rect 7096 51648 7112 51712
rect 7176 51648 7192 51712
rect 7256 51648 7264 51712
rect 6944 50624 7264 51648
rect 6944 50560 6952 50624
rect 7016 50560 7032 50624
rect 7096 50560 7112 50624
rect 7176 50560 7192 50624
rect 7256 50560 7264 50624
rect 6944 49536 7264 50560
rect 6944 49472 6952 49536
rect 7016 49472 7032 49536
rect 7096 49472 7112 49536
rect 7176 49472 7192 49536
rect 7256 49472 7264 49536
rect 6944 48448 7264 49472
rect 6944 48384 6952 48448
rect 7016 48384 7032 48448
rect 7096 48384 7112 48448
rect 7176 48384 7192 48448
rect 7256 48384 7264 48448
rect 6944 48294 7264 48384
rect 6944 48058 6986 48294
rect 7222 48058 7264 48294
rect 6944 47360 7264 48058
rect 6944 47296 6952 47360
rect 7016 47296 7032 47360
rect 7096 47296 7112 47360
rect 7176 47296 7192 47360
rect 7256 47296 7264 47360
rect 6944 46272 7264 47296
rect 6944 46208 6952 46272
rect 7016 46208 7032 46272
rect 7096 46208 7112 46272
rect 7176 46208 7192 46272
rect 7256 46208 7264 46272
rect 6944 45184 7264 46208
rect 6944 45120 6952 45184
rect 7016 45120 7032 45184
rect 7096 45120 7112 45184
rect 7176 45120 7192 45184
rect 7256 45120 7264 45184
rect 6944 44096 7264 45120
rect 6944 44032 6952 44096
rect 7016 44032 7032 44096
rect 7096 44032 7112 44096
rect 7176 44032 7192 44096
rect 7256 44032 7264 44096
rect 6944 43294 7264 44032
rect 6944 43058 6986 43294
rect 7222 43058 7264 43294
rect 6944 43008 7264 43058
rect 6944 42944 6952 43008
rect 7016 42944 7032 43008
rect 7096 42944 7112 43008
rect 7176 42944 7192 43008
rect 7256 42944 7264 43008
rect 6944 41920 7264 42944
rect 6944 41856 6952 41920
rect 7016 41856 7032 41920
rect 7096 41856 7112 41920
rect 7176 41856 7192 41920
rect 7256 41856 7264 41920
rect 6944 40832 7264 41856
rect 6944 40768 6952 40832
rect 7016 40768 7032 40832
rect 7096 40768 7112 40832
rect 7176 40768 7192 40832
rect 7256 40768 7264 40832
rect 6944 39744 7264 40768
rect 6944 39680 6952 39744
rect 7016 39680 7032 39744
rect 7096 39680 7112 39744
rect 7176 39680 7192 39744
rect 7256 39680 7264 39744
rect 6944 38656 7264 39680
rect 6944 38592 6952 38656
rect 7016 38592 7032 38656
rect 7096 38592 7112 38656
rect 7176 38592 7192 38656
rect 7256 38592 7264 38656
rect 6944 38294 7264 38592
rect 6944 38058 6986 38294
rect 7222 38058 7264 38294
rect 6944 37568 7264 38058
rect 6944 37504 6952 37568
rect 7016 37504 7032 37568
rect 7096 37504 7112 37568
rect 7176 37504 7192 37568
rect 7256 37504 7264 37568
rect 6944 36480 7264 37504
rect 6944 36416 6952 36480
rect 7016 36416 7032 36480
rect 7096 36416 7112 36480
rect 7176 36416 7192 36480
rect 7256 36416 7264 36480
rect 6944 35392 7264 36416
rect 6944 35328 6952 35392
rect 7016 35328 7032 35392
rect 7096 35328 7112 35392
rect 7176 35328 7192 35392
rect 7256 35328 7264 35392
rect 6944 34304 7264 35328
rect 6944 34240 6952 34304
rect 7016 34240 7032 34304
rect 7096 34240 7112 34304
rect 7176 34240 7192 34304
rect 7256 34240 7264 34304
rect 6944 33294 7264 34240
rect 6944 33216 6986 33294
rect 7222 33216 7264 33294
rect 6944 33152 6952 33216
rect 7256 33152 7264 33216
rect 6944 33058 6986 33152
rect 7222 33058 7264 33152
rect 6944 32128 7264 33058
rect 6944 32064 6952 32128
rect 7016 32064 7032 32128
rect 7096 32064 7112 32128
rect 7176 32064 7192 32128
rect 7256 32064 7264 32128
rect 6944 31040 7264 32064
rect 6944 30976 6952 31040
rect 7016 30976 7032 31040
rect 7096 30976 7112 31040
rect 7176 30976 7192 31040
rect 7256 30976 7264 31040
rect 6944 29952 7264 30976
rect 6944 29888 6952 29952
rect 7016 29888 7032 29952
rect 7096 29888 7112 29952
rect 7176 29888 7192 29952
rect 7256 29888 7264 29952
rect 6944 28864 7264 29888
rect 6944 28800 6952 28864
rect 7016 28800 7032 28864
rect 7096 28800 7112 28864
rect 7176 28800 7192 28864
rect 7256 28800 7264 28864
rect 6944 28294 7264 28800
rect 6944 28058 6986 28294
rect 7222 28058 7264 28294
rect 6944 27776 7264 28058
rect 6944 27712 6952 27776
rect 7016 27712 7032 27776
rect 7096 27712 7112 27776
rect 7176 27712 7192 27776
rect 7256 27712 7264 27776
rect 6944 26688 7264 27712
rect 6944 26624 6952 26688
rect 7016 26624 7032 26688
rect 7096 26624 7112 26688
rect 7176 26624 7192 26688
rect 7256 26624 7264 26688
rect 6944 25600 7264 26624
rect 6944 25536 6952 25600
rect 7016 25536 7032 25600
rect 7096 25536 7112 25600
rect 7176 25536 7192 25600
rect 7256 25536 7264 25600
rect 6944 24512 7264 25536
rect 6944 24448 6952 24512
rect 7016 24448 7032 24512
rect 7096 24448 7112 24512
rect 7176 24448 7192 24512
rect 7256 24448 7264 24512
rect 6944 23424 7264 24448
rect 6944 23360 6952 23424
rect 7016 23360 7032 23424
rect 7096 23360 7112 23424
rect 7176 23360 7192 23424
rect 7256 23360 7264 23424
rect 6944 23294 7264 23360
rect 6944 23058 6986 23294
rect 7222 23058 7264 23294
rect 6944 22336 7264 23058
rect 6944 22272 6952 22336
rect 7016 22272 7032 22336
rect 7096 22272 7112 22336
rect 7176 22272 7192 22336
rect 7256 22272 7264 22336
rect 6944 21248 7264 22272
rect 6944 21184 6952 21248
rect 7016 21184 7032 21248
rect 7096 21184 7112 21248
rect 7176 21184 7192 21248
rect 7256 21184 7264 21248
rect 6944 20160 7264 21184
rect 6944 20096 6952 20160
rect 7016 20096 7032 20160
rect 7096 20096 7112 20160
rect 7176 20096 7192 20160
rect 7256 20096 7264 20160
rect 6944 19072 7264 20096
rect 6944 19008 6952 19072
rect 7016 19008 7032 19072
rect 7096 19008 7112 19072
rect 7176 19008 7192 19072
rect 7256 19008 7264 19072
rect 6944 18294 7264 19008
rect 6944 18058 6986 18294
rect 7222 18058 7264 18294
rect 6944 17984 7264 18058
rect 6944 17920 6952 17984
rect 7016 17920 7032 17984
rect 7096 17920 7112 17984
rect 7176 17920 7192 17984
rect 7256 17920 7264 17984
rect 6944 16896 7264 17920
rect 6944 16832 6952 16896
rect 7016 16832 7032 16896
rect 7096 16832 7112 16896
rect 7176 16832 7192 16896
rect 7256 16832 7264 16896
rect 6944 15808 7264 16832
rect 6944 15744 6952 15808
rect 7016 15744 7032 15808
rect 7096 15744 7112 15808
rect 7176 15744 7192 15808
rect 7256 15744 7264 15808
rect 6944 14720 7264 15744
rect 6944 14656 6952 14720
rect 7016 14656 7032 14720
rect 7096 14656 7112 14720
rect 7176 14656 7192 14720
rect 7256 14656 7264 14720
rect 6944 13632 7264 14656
rect 6944 13568 6952 13632
rect 7016 13568 7032 13632
rect 7096 13568 7112 13632
rect 7176 13568 7192 13632
rect 7256 13568 7264 13632
rect 6944 13294 7264 13568
rect 6944 13058 6986 13294
rect 7222 13058 7264 13294
rect 6944 12544 7264 13058
rect 6944 12480 6952 12544
rect 7016 12480 7032 12544
rect 7096 12480 7112 12544
rect 7176 12480 7192 12544
rect 7256 12480 7264 12544
rect 6944 11456 7264 12480
rect 6944 11392 6952 11456
rect 7016 11392 7032 11456
rect 7096 11392 7112 11456
rect 7176 11392 7192 11456
rect 7256 11392 7264 11456
rect 6944 10368 7264 11392
rect 6944 10304 6952 10368
rect 7016 10304 7032 10368
rect 7096 10304 7112 10368
rect 7176 10304 7192 10368
rect 7256 10304 7264 10368
rect 6944 9280 7264 10304
rect 6944 9216 6952 9280
rect 7016 9216 7032 9280
rect 7096 9216 7112 9280
rect 7176 9216 7192 9280
rect 7256 9216 7264 9280
rect 6944 8294 7264 9216
rect 6944 8192 6986 8294
rect 7222 8192 7264 8294
rect 6944 8128 6952 8192
rect 7256 8128 7264 8192
rect 6944 8058 6986 8128
rect 7222 8058 7264 8128
rect 6944 7104 7264 8058
rect 6944 7040 6952 7104
rect 7016 7040 7032 7104
rect 7096 7040 7112 7104
rect 7176 7040 7192 7104
rect 7256 7040 7264 7104
rect 6944 6016 7264 7040
rect 6944 5952 6952 6016
rect 7016 5952 7032 6016
rect 7096 5952 7112 6016
rect 7176 5952 7192 6016
rect 7256 5952 7264 6016
rect 6944 4928 7264 5952
rect 6944 4864 6952 4928
rect 7016 4864 7032 4928
rect 7096 4864 7112 4928
rect 7176 4864 7192 4928
rect 7256 4864 7264 4928
rect 6944 3840 7264 4864
rect 6944 3776 6952 3840
rect 7016 3776 7032 3840
rect 7096 3776 7112 3840
rect 7176 3776 7192 3840
rect 7256 3776 7264 3840
rect 6944 3294 7264 3776
rect 6944 3058 6986 3294
rect 7222 3058 7264 3294
rect 6944 2752 7264 3058
rect 6944 2688 6952 2752
rect 7016 2688 7032 2752
rect 7096 2688 7112 2752
rect 7176 2688 7192 2752
rect 7256 2688 7264 2752
rect 6944 2128 7264 2688
rect 7604 69664 7924 69680
rect 7604 69600 7612 69664
rect 7676 69600 7692 69664
rect 7756 69600 7772 69664
rect 7836 69600 7852 69664
rect 7916 69600 7924 69664
rect 7604 68954 7924 69600
rect 7604 68718 7646 68954
rect 7882 68718 7924 68954
rect 7604 68576 7924 68718
rect 7604 68512 7612 68576
rect 7676 68512 7692 68576
rect 7756 68512 7772 68576
rect 7836 68512 7852 68576
rect 7916 68512 7924 68576
rect 7604 67488 7924 68512
rect 7604 67424 7612 67488
rect 7676 67424 7692 67488
rect 7756 67424 7772 67488
rect 7836 67424 7852 67488
rect 7916 67424 7924 67488
rect 7604 66400 7924 67424
rect 7604 66336 7612 66400
rect 7676 66336 7692 66400
rect 7756 66336 7772 66400
rect 7836 66336 7852 66400
rect 7916 66336 7924 66400
rect 7604 65312 7924 66336
rect 7604 65248 7612 65312
rect 7676 65248 7692 65312
rect 7756 65248 7772 65312
rect 7836 65248 7852 65312
rect 7916 65248 7924 65312
rect 7604 64224 7924 65248
rect 7604 64160 7612 64224
rect 7676 64160 7692 64224
rect 7756 64160 7772 64224
rect 7836 64160 7852 64224
rect 7916 64160 7924 64224
rect 7604 63954 7924 64160
rect 7604 63718 7646 63954
rect 7882 63718 7924 63954
rect 7604 63136 7924 63718
rect 7604 63072 7612 63136
rect 7676 63072 7692 63136
rect 7756 63072 7772 63136
rect 7836 63072 7852 63136
rect 7916 63072 7924 63136
rect 7604 62048 7924 63072
rect 7604 61984 7612 62048
rect 7676 61984 7692 62048
rect 7756 61984 7772 62048
rect 7836 61984 7852 62048
rect 7916 61984 7924 62048
rect 7604 60960 7924 61984
rect 7604 60896 7612 60960
rect 7676 60896 7692 60960
rect 7756 60896 7772 60960
rect 7836 60896 7852 60960
rect 7916 60896 7924 60960
rect 7604 59872 7924 60896
rect 7604 59808 7612 59872
rect 7676 59808 7692 59872
rect 7756 59808 7772 59872
rect 7836 59808 7852 59872
rect 7916 59808 7924 59872
rect 7604 58954 7924 59808
rect 7604 58784 7646 58954
rect 7882 58784 7924 58954
rect 7604 58720 7612 58784
rect 7916 58720 7924 58784
rect 7604 58718 7646 58720
rect 7882 58718 7924 58720
rect 7604 57696 7924 58718
rect 7604 57632 7612 57696
rect 7676 57632 7692 57696
rect 7756 57632 7772 57696
rect 7836 57632 7852 57696
rect 7916 57632 7924 57696
rect 7604 56608 7924 57632
rect 7604 56544 7612 56608
rect 7676 56544 7692 56608
rect 7756 56544 7772 56608
rect 7836 56544 7852 56608
rect 7916 56544 7924 56608
rect 7604 55520 7924 56544
rect 7604 55456 7612 55520
rect 7676 55456 7692 55520
rect 7756 55456 7772 55520
rect 7836 55456 7852 55520
rect 7916 55456 7924 55520
rect 7604 54432 7924 55456
rect 7604 54368 7612 54432
rect 7676 54368 7692 54432
rect 7756 54368 7772 54432
rect 7836 54368 7852 54432
rect 7916 54368 7924 54432
rect 7604 53954 7924 54368
rect 7604 53718 7646 53954
rect 7882 53718 7924 53954
rect 7604 53344 7924 53718
rect 7604 53280 7612 53344
rect 7676 53280 7692 53344
rect 7756 53280 7772 53344
rect 7836 53280 7852 53344
rect 7916 53280 7924 53344
rect 7604 52256 7924 53280
rect 7604 52192 7612 52256
rect 7676 52192 7692 52256
rect 7756 52192 7772 52256
rect 7836 52192 7852 52256
rect 7916 52192 7924 52256
rect 7604 51168 7924 52192
rect 7604 51104 7612 51168
rect 7676 51104 7692 51168
rect 7756 51104 7772 51168
rect 7836 51104 7852 51168
rect 7916 51104 7924 51168
rect 7604 50080 7924 51104
rect 7604 50016 7612 50080
rect 7676 50016 7692 50080
rect 7756 50016 7772 50080
rect 7836 50016 7852 50080
rect 7916 50016 7924 50080
rect 7604 48992 7924 50016
rect 7604 48928 7612 48992
rect 7676 48954 7692 48992
rect 7756 48954 7772 48992
rect 7836 48954 7852 48992
rect 7916 48928 7924 48992
rect 7604 48718 7646 48928
rect 7882 48718 7924 48928
rect 7604 47904 7924 48718
rect 7604 47840 7612 47904
rect 7676 47840 7692 47904
rect 7756 47840 7772 47904
rect 7836 47840 7852 47904
rect 7916 47840 7924 47904
rect 7604 46816 7924 47840
rect 7604 46752 7612 46816
rect 7676 46752 7692 46816
rect 7756 46752 7772 46816
rect 7836 46752 7852 46816
rect 7916 46752 7924 46816
rect 7604 45728 7924 46752
rect 7604 45664 7612 45728
rect 7676 45664 7692 45728
rect 7756 45664 7772 45728
rect 7836 45664 7852 45728
rect 7916 45664 7924 45728
rect 7604 44640 7924 45664
rect 7604 44576 7612 44640
rect 7676 44576 7692 44640
rect 7756 44576 7772 44640
rect 7836 44576 7852 44640
rect 7916 44576 7924 44640
rect 7604 43954 7924 44576
rect 7604 43718 7646 43954
rect 7882 43718 7924 43954
rect 7604 43552 7924 43718
rect 7604 43488 7612 43552
rect 7676 43488 7692 43552
rect 7756 43488 7772 43552
rect 7836 43488 7852 43552
rect 7916 43488 7924 43552
rect 7604 42464 7924 43488
rect 7604 42400 7612 42464
rect 7676 42400 7692 42464
rect 7756 42400 7772 42464
rect 7836 42400 7852 42464
rect 7916 42400 7924 42464
rect 7604 41376 7924 42400
rect 7604 41312 7612 41376
rect 7676 41312 7692 41376
rect 7756 41312 7772 41376
rect 7836 41312 7852 41376
rect 7916 41312 7924 41376
rect 7604 40288 7924 41312
rect 7604 40224 7612 40288
rect 7676 40224 7692 40288
rect 7756 40224 7772 40288
rect 7836 40224 7852 40288
rect 7916 40224 7924 40288
rect 7604 39200 7924 40224
rect 7604 39136 7612 39200
rect 7676 39136 7692 39200
rect 7756 39136 7772 39200
rect 7836 39136 7852 39200
rect 7916 39136 7924 39200
rect 7604 38954 7924 39136
rect 7604 38718 7646 38954
rect 7882 38718 7924 38954
rect 7604 38112 7924 38718
rect 7604 38048 7612 38112
rect 7676 38048 7692 38112
rect 7756 38048 7772 38112
rect 7836 38048 7852 38112
rect 7916 38048 7924 38112
rect 7604 37024 7924 38048
rect 7604 36960 7612 37024
rect 7676 36960 7692 37024
rect 7756 36960 7772 37024
rect 7836 36960 7852 37024
rect 7916 36960 7924 37024
rect 7604 35936 7924 36960
rect 7604 35872 7612 35936
rect 7676 35872 7692 35936
rect 7756 35872 7772 35936
rect 7836 35872 7852 35936
rect 7916 35872 7924 35936
rect 7604 34848 7924 35872
rect 7604 34784 7612 34848
rect 7676 34784 7692 34848
rect 7756 34784 7772 34848
rect 7836 34784 7852 34848
rect 7916 34784 7924 34848
rect 7604 33954 7924 34784
rect 7604 33760 7646 33954
rect 7882 33760 7924 33954
rect 7604 33696 7612 33760
rect 7676 33696 7692 33718
rect 7756 33696 7772 33718
rect 7836 33696 7852 33718
rect 7916 33696 7924 33760
rect 7604 32672 7924 33696
rect 7604 32608 7612 32672
rect 7676 32608 7692 32672
rect 7756 32608 7772 32672
rect 7836 32608 7852 32672
rect 7916 32608 7924 32672
rect 7604 31584 7924 32608
rect 7604 31520 7612 31584
rect 7676 31520 7692 31584
rect 7756 31520 7772 31584
rect 7836 31520 7852 31584
rect 7916 31520 7924 31584
rect 7604 30496 7924 31520
rect 7604 30432 7612 30496
rect 7676 30432 7692 30496
rect 7756 30432 7772 30496
rect 7836 30432 7852 30496
rect 7916 30432 7924 30496
rect 7604 29408 7924 30432
rect 7604 29344 7612 29408
rect 7676 29344 7692 29408
rect 7756 29344 7772 29408
rect 7836 29344 7852 29408
rect 7916 29344 7924 29408
rect 7604 28954 7924 29344
rect 7604 28718 7646 28954
rect 7882 28718 7924 28954
rect 7604 28320 7924 28718
rect 7604 28256 7612 28320
rect 7676 28256 7692 28320
rect 7756 28256 7772 28320
rect 7836 28256 7852 28320
rect 7916 28256 7924 28320
rect 7604 27232 7924 28256
rect 7604 27168 7612 27232
rect 7676 27168 7692 27232
rect 7756 27168 7772 27232
rect 7836 27168 7852 27232
rect 7916 27168 7924 27232
rect 7604 26144 7924 27168
rect 7604 26080 7612 26144
rect 7676 26080 7692 26144
rect 7756 26080 7772 26144
rect 7836 26080 7852 26144
rect 7916 26080 7924 26144
rect 7604 25056 7924 26080
rect 7604 24992 7612 25056
rect 7676 24992 7692 25056
rect 7756 24992 7772 25056
rect 7836 24992 7852 25056
rect 7916 24992 7924 25056
rect 7604 23968 7924 24992
rect 7604 23904 7612 23968
rect 7676 23954 7692 23968
rect 7756 23954 7772 23968
rect 7836 23954 7852 23968
rect 7916 23904 7924 23968
rect 7604 23718 7646 23904
rect 7882 23718 7924 23904
rect 7604 22880 7924 23718
rect 7604 22816 7612 22880
rect 7676 22816 7692 22880
rect 7756 22816 7772 22880
rect 7836 22816 7852 22880
rect 7916 22816 7924 22880
rect 7604 21792 7924 22816
rect 7604 21728 7612 21792
rect 7676 21728 7692 21792
rect 7756 21728 7772 21792
rect 7836 21728 7852 21792
rect 7916 21728 7924 21792
rect 7604 20704 7924 21728
rect 7604 20640 7612 20704
rect 7676 20640 7692 20704
rect 7756 20640 7772 20704
rect 7836 20640 7852 20704
rect 7916 20640 7924 20704
rect 7604 19616 7924 20640
rect 7604 19552 7612 19616
rect 7676 19552 7692 19616
rect 7756 19552 7772 19616
rect 7836 19552 7852 19616
rect 7916 19552 7924 19616
rect 7604 18954 7924 19552
rect 7604 18718 7646 18954
rect 7882 18718 7924 18954
rect 7604 18528 7924 18718
rect 7604 18464 7612 18528
rect 7676 18464 7692 18528
rect 7756 18464 7772 18528
rect 7836 18464 7852 18528
rect 7916 18464 7924 18528
rect 7604 17440 7924 18464
rect 7604 17376 7612 17440
rect 7676 17376 7692 17440
rect 7756 17376 7772 17440
rect 7836 17376 7852 17440
rect 7916 17376 7924 17440
rect 7604 16352 7924 17376
rect 7604 16288 7612 16352
rect 7676 16288 7692 16352
rect 7756 16288 7772 16352
rect 7836 16288 7852 16352
rect 7916 16288 7924 16352
rect 7604 15264 7924 16288
rect 7604 15200 7612 15264
rect 7676 15200 7692 15264
rect 7756 15200 7772 15264
rect 7836 15200 7852 15264
rect 7916 15200 7924 15264
rect 7604 14176 7924 15200
rect 7604 14112 7612 14176
rect 7676 14112 7692 14176
rect 7756 14112 7772 14176
rect 7836 14112 7852 14176
rect 7916 14112 7924 14176
rect 7604 13954 7924 14112
rect 7604 13718 7646 13954
rect 7882 13718 7924 13954
rect 7604 13088 7924 13718
rect 7604 13024 7612 13088
rect 7676 13024 7692 13088
rect 7756 13024 7772 13088
rect 7836 13024 7852 13088
rect 7916 13024 7924 13088
rect 7604 12000 7924 13024
rect 7604 11936 7612 12000
rect 7676 11936 7692 12000
rect 7756 11936 7772 12000
rect 7836 11936 7852 12000
rect 7916 11936 7924 12000
rect 7604 10912 7924 11936
rect 7604 10848 7612 10912
rect 7676 10848 7692 10912
rect 7756 10848 7772 10912
rect 7836 10848 7852 10912
rect 7916 10848 7924 10912
rect 7604 9824 7924 10848
rect 7604 9760 7612 9824
rect 7676 9760 7692 9824
rect 7756 9760 7772 9824
rect 7836 9760 7852 9824
rect 7916 9760 7924 9824
rect 7604 8954 7924 9760
rect 7604 8736 7646 8954
rect 7882 8736 7924 8954
rect 7604 8672 7612 8736
rect 7676 8672 7692 8718
rect 7756 8672 7772 8718
rect 7836 8672 7852 8718
rect 7916 8672 7924 8736
rect 7604 7648 7924 8672
rect 7604 7584 7612 7648
rect 7676 7584 7692 7648
rect 7756 7584 7772 7648
rect 7836 7584 7852 7648
rect 7916 7584 7924 7648
rect 7604 6560 7924 7584
rect 7604 6496 7612 6560
rect 7676 6496 7692 6560
rect 7756 6496 7772 6560
rect 7836 6496 7852 6560
rect 7916 6496 7924 6560
rect 7604 5472 7924 6496
rect 7604 5408 7612 5472
rect 7676 5408 7692 5472
rect 7756 5408 7772 5472
rect 7836 5408 7852 5472
rect 7916 5408 7924 5472
rect 7604 4384 7924 5408
rect 7604 4320 7612 4384
rect 7676 4320 7692 4384
rect 7756 4320 7772 4384
rect 7836 4320 7852 4384
rect 7916 4320 7924 4384
rect 7604 3954 7924 4320
rect 7604 3718 7646 3954
rect 7882 3718 7924 3954
rect 7604 3296 7924 3718
rect 7604 3232 7612 3296
rect 7676 3232 7692 3296
rect 7756 3232 7772 3296
rect 7836 3232 7852 3296
rect 7916 3232 7924 3296
rect 7604 2208 7924 3232
rect 7604 2144 7612 2208
rect 7676 2144 7692 2208
rect 7756 2144 7772 2208
rect 7836 2144 7852 2208
rect 7916 2144 7924 2208
rect 7604 2128 7924 2144
rect 11944 69120 12264 69680
rect 11944 69056 11952 69120
rect 12016 69056 12032 69120
rect 12096 69056 12112 69120
rect 12176 69056 12192 69120
rect 12256 69056 12264 69120
rect 11944 68294 12264 69056
rect 11944 68058 11986 68294
rect 12222 68058 12264 68294
rect 11944 68032 12264 68058
rect 11944 67968 11952 68032
rect 12016 67968 12032 68032
rect 12096 67968 12112 68032
rect 12176 67968 12192 68032
rect 12256 67968 12264 68032
rect 11944 66944 12264 67968
rect 11944 66880 11952 66944
rect 12016 66880 12032 66944
rect 12096 66880 12112 66944
rect 12176 66880 12192 66944
rect 12256 66880 12264 66944
rect 11944 65856 12264 66880
rect 11944 65792 11952 65856
rect 12016 65792 12032 65856
rect 12096 65792 12112 65856
rect 12176 65792 12192 65856
rect 12256 65792 12264 65856
rect 11944 64768 12264 65792
rect 11944 64704 11952 64768
rect 12016 64704 12032 64768
rect 12096 64704 12112 64768
rect 12176 64704 12192 64768
rect 12256 64704 12264 64768
rect 11944 63680 12264 64704
rect 11944 63616 11952 63680
rect 12016 63616 12032 63680
rect 12096 63616 12112 63680
rect 12176 63616 12192 63680
rect 12256 63616 12264 63680
rect 11944 63294 12264 63616
rect 11944 63058 11986 63294
rect 12222 63058 12264 63294
rect 11944 62592 12264 63058
rect 11944 62528 11952 62592
rect 12016 62528 12032 62592
rect 12096 62528 12112 62592
rect 12176 62528 12192 62592
rect 12256 62528 12264 62592
rect 11944 61504 12264 62528
rect 11944 61440 11952 61504
rect 12016 61440 12032 61504
rect 12096 61440 12112 61504
rect 12176 61440 12192 61504
rect 12256 61440 12264 61504
rect 11944 60416 12264 61440
rect 11944 60352 11952 60416
rect 12016 60352 12032 60416
rect 12096 60352 12112 60416
rect 12176 60352 12192 60416
rect 12256 60352 12264 60416
rect 11944 59328 12264 60352
rect 11944 59264 11952 59328
rect 12016 59264 12032 59328
rect 12096 59264 12112 59328
rect 12176 59264 12192 59328
rect 12256 59264 12264 59328
rect 11944 58294 12264 59264
rect 11944 58240 11986 58294
rect 12222 58240 12264 58294
rect 11944 58176 11952 58240
rect 12256 58176 12264 58240
rect 11944 58058 11986 58176
rect 12222 58058 12264 58176
rect 11944 57152 12264 58058
rect 11944 57088 11952 57152
rect 12016 57088 12032 57152
rect 12096 57088 12112 57152
rect 12176 57088 12192 57152
rect 12256 57088 12264 57152
rect 11944 56064 12264 57088
rect 11944 56000 11952 56064
rect 12016 56000 12032 56064
rect 12096 56000 12112 56064
rect 12176 56000 12192 56064
rect 12256 56000 12264 56064
rect 11944 54976 12264 56000
rect 11944 54912 11952 54976
rect 12016 54912 12032 54976
rect 12096 54912 12112 54976
rect 12176 54912 12192 54976
rect 12256 54912 12264 54976
rect 11944 53888 12264 54912
rect 11944 53824 11952 53888
rect 12016 53824 12032 53888
rect 12096 53824 12112 53888
rect 12176 53824 12192 53888
rect 12256 53824 12264 53888
rect 11944 53294 12264 53824
rect 11944 53058 11986 53294
rect 12222 53058 12264 53294
rect 11944 52800 12264 53058
rect 11944 52736 11952 52800
rect 12016 52736 12032 52800
rect 12096 52736 12112 52800
rect 12176 52736 12192 52800
rect 12256 52736 12264 52800
rect 11944 51712 12264 52736
rect 11944 51648 11952 51712
rect 12016 51648 12032 51712
rect 12096 51648 12112 51712
rect 12176 51648 12192 51712
rect 12256 51648 12264 51712
rect 11944 50624 12264 51648
rect 11944 50560 11952 50624
rect 12016 50560 12032 50624
rect 12096 50560 12112 50624
rect 12176 50560 12192 50624
rect 12256 50560 12264 50624
rect 11944 49536 12264 50560
rect 11944 49472 11952 49536
rect 12016 49472 12032 49536
rect 12096 49472 12112 49536
rect 12176 49472 12192 49536
rect 12256 49472 12264 49536
rect 11944 48448 12264 49472
rect 11944 48384 11952 48448
rect 12016 48384 12032 48448
rect 12096 48384 12112 48448
rect 12176 48384 12192 48448
rect 12256 48384 12264 48448
rect 11944 48294 12264 48384
rect 11944 48058 11986 48294
rect 12222 48058 12264 48294
rect 11944 47360 12264 48058
rect 11944 47296 11952 47360
rect 12016 47296 12032 47360
rect 12096 47296 12112 47360
rect 12176 47296 12192 47360
rect 12256 47296 12264 47360
rect 11944 46272 12264 47296
rect 11944 46208 11952 46272
rect 12016 46208 12032 46272
rect 12096 46208 12112 46272
rect 12176 46208 12192 46272
rect 12256 46208 12264 46272
rect 11944 45184 12264 46208
rect 11944 45120 11952 45184
rect 12016 45120 12032 45184
rect 12096 45120 12112 45184
rect 12176 45120 12192 45184
rect 12256 45120 12264 45184
rect 11944 44096 12264 45120
rect 11944 44032 11952 44096
rect 12016 44032 12032 44096
rect 12096 44032 12112 44096
rect 12176 44032 12192 44096
rect 12256 44032 12264 44096
rect 11944 43294 12264 44032
rect 11944 43058 11986 43294
rect 12222 43058 12264 43294
rect 11944 43008 12264 43058
rect 11944 42944 11952 43008
rect 12016 42944 12032 43008
rect 12096 42944 12112 43008
rect 12176 42944 12192 43008
rect 12256 42944 12264 43008
rect 11944 41920 12264 42944
rect 11944 41856 11952 41920
rect 12016 41856 12032 41920
rect 12096 41856 12112 41920
rect 12176 41856 12192 41920
rect 12256 41856 12264 41920
rect 11944 40832 12264 41856
rect 11944 40768 11952 40832
rect 12016 40768 12032 40832
rect 12096 40768 12112 40832
rect 12176 40768 12192 40832
rect 12256 40768 12264 40832
rect 11944 39744 12264 40768
rect 11944 39680 11952 39744
rect 12016 39680 12032 39744
rect 12096 39680 12112 39744
rect 12176 39680 12192 39744
rect 12256 39680 12264 39744
rect 11944 38656 12264 39680
rect 11944 38592 11952 38656
rect 12016 38592 12032 38656
rect 12096 38592 12112 38656
rect 12176 38592 12192 38656
rect 12256 38592 12264 38656
rect 11944 38294 12264 38592
rect 11944 38058 11986 38294
rect 12222 38058 12264 38294
rect 11944 37568 12264 38058
rect 11944 37504 11952 37568
rect 12016 37504 12032 37568
rect 12096 37504 12112 37568
rect 12176 37504 12192 37568
rect 12256 37504 12264 37568
rect 11944 36480 12264 37504
rect 11944 36416 11952 36480
rect 12016 36416 12032 36480
rect 12096 36416 12112 36480
rect 12176 36416 12192 36480
rect 12256 36416 12264 36480
rect 11944 35392 12264 36416
rect 11944 35328 11952 35392
rect 12016 35328 12032 35392
rect 12096 35328 12112 35392
rect 12176 35328 12192 35392
rect 12256 35328 12264 35392
rect 11944 34304 12264 35328
rect 11944 34240 11952 34304
rect 12016 34240 12032 34304
rect 12096 34240 12112 34304
rect 12176 34240 12192 34304
rect 12256 34240 12264 34304
rect 11944 33294 12264 34240
rect 11944 33216 11986 33294
rect 12222 33216 12264 33294
rect 11944 33152 11952 33216
rect 12256 33152 12264 33216
rect 11944 33058 11986 33152
rect 12222 33058 12264 33152
rect 11944 32128 12264 33058
rect 11944 32064 11952 32128
rect 12016 32064 12032 32128
rect 12096 32064 12112 32128
rect 12176 32064 12192 32128
rect 12256 32064 12264 32128
rect 11944 31040 12264 32064
rect 11944 30976 11952 31040
rect 12016 30976 12032 31040
rect 12096 30976 12112 31040
rect 12176 30976 12192 31040
rect 12256 30976 12264 31040
rect 11944 29952 12264 30976
rect 11944 29888 11952 29952
rect 12016 29888 12032 29952
rect 12096 29888 12112 29952
rect 12176 29888 12192 29952
rect 12256 29888 12264 29952
rect 11944 28864 12264 29888
rect 11944 28800 11952 28864
rect 12016 28800 12032 28864
rect 12096 28800 12112 28864
rect 12176 28800 12192 28864
rect 12256 28800 12264 28864
rect 11944 28294 12264 28800
rect 11944 28058 11986 28294
rect 12222 28058 12264 28294
rect 11944 27776 12264 28058
rect 11944 27712 11952 27776
rect 12016 27712 12032 27776
rect 12096 27712 12112 27776
rect 12176 27712 12192 27776
rect 12256 27712 12264 27776
rect 11944 26688 12264 27712
rect 11944 26624 11952 26688
rect 12016 26624 12032 26688
rect 12096 26624 12112 26688
rect 12176 26624 12192 26688
rect 12256 26624 12264 26688
rect 11944 25600 12264 26624
rect 11944 25536 11952 25600
rect 12016 25536 12032 25600
rect 12096 25536 12112 25600
rect 12176 25536 12192 25600
rect 12256 25536 12264 25600
rect 11944 24512 12264 25536
rect 11944 24448 11952 24512
rect 12016 24448 12032 24512
rect 12096 24448 12112 24512
rect 12176 24448 12192 24512
rect 12256 24448 12264 24512
rect 11944 23424 12264 24448
rect 11944 23360 11952 23424
rect 12016 23360 12032 23424
rect 12096 23360 12112 23424
rect 12176 23360 12192 23424
rect 12256 23360 12264 23424
rect 11944 23294 12264 23360
rect 11944 23058 11986 23294
rect 12222 23058 12264 23294
rect 11944 22336 12264 23058
rect 11944 22272 11952 22336
rect 12016 22272 12032 22336
rect 12096 22272 12112 22336
rect 12176 22272 12192 22336
rect 12256 22272 12264 22336
rect 11944 21248 12264 22272
rect 11944 21184 11952 21248
rect 12016 21184 12032 21248
rect 12096 21184 12112 21248
rect 12176 21184 12192 21248
rect 12256 21184 12264 21248
rect 11944 20160 12264 21184
rect 11944 20096 11952 20160
rect 12016 20096 12032 20160
rect 12096 20096 12112 20160
rect 12176 20096 12192 20160
rect 12256 20096 12264 20160
rect 11944 19072 12264 20096
rect 11944 19008 11952 19072
rect 12016 19008 12032 19072
rect 12096 19008 12112 19072
rect 12176 19008 12192 19072
rect 12256 19008 12264 19072
rect 11944 18294 12264 19008
rect 11944 18058 11986 18294
rect 12222 18058 12264 18294
rect 11944 17984 12264 18058
rect 11944 17920 11952 17984
rect 12016 17920 12032 17984
rect 12096 17920 12112 17984
rect 12176 17920 12192 17984
rect 12256 17920 12264 17984
rect 11944 16896 12264 17920
rect 11944 16832 11952 16896
rect 12016 16832 12032 16896
rect 12096 16832 12112 16896
rect 12176 16832 12192 16896
rect 12256 16832 12264 16896
rect 11944 15808 12264 16832
rect 11944 15744 11952 15808
rect 12016 15744 12032 15808
rect 12096 15744 12112 15808
rect 12176 15744 12192 15808
rect 12256 15744 12264 15808
rect 11944 14720 12264 15744
rect 11944 14656 11952 14720
rect 12016 14656 12032 14720
rect 12096 14656 12112 14720
rect 12176 14656 12192 14720
rect 12256 14656 12264 14720
rect 11944 13632 12264 14656
rect 11944 13568 11952 13632
rect 12016 13568 12032 13632
rect 12096 13568 12112 13632
rect 12176 13568 12192 13632
rect 12256 13568 12264 13632
rect 11944 13294 12264 13568
rect 11944 13058 11986 13294
rect 12222 13058 12264 13294
rect 11944 12544 12264 13058
rect 11944 12480 11952 12544
rect 12016 12480 12032 12544
rect 12096 12480 12112 12544
rect 12176 12480 12192 12544
rect 12256 12480 12264 12544
rect 11944 11456 12264 12480
rect 11944 11392 11952 11456
rect 12016 11392 12032 11456
rect 12096 11392 12112 11456
rect 12176 11392 12192 11456
rect 12256 11392 12264 11456
rect 11944 10368 12264 11392
rect 11944 10304 11952 10368
rect 12016 10304 12032 10368
rect 12096 10304 12112 10368
rect 12176 10304 12192 10368
rect 12256 10304 12264 10368
rect 11944 9280 12264 10304
rect 11944 9216 11952 9280
rect 12016 9216 12032 9280
rect 12096 9216 12112 9280
rect 12176 9216 12192 9280
rect 12256 9216 12264 9280
rect 11944 8294 12264 9216
rect 11944 8192 11986 8294
rect 12222 8192 12264 8294
rect 11944 8128 11952 8192
rect 12256 8128 12264 8192
rect 11944 8058 11986 8128
rect 12222 8058 12264 8128
rect 11944 7104 12264 8058
rect 11944 7040 11952 7104
rect 12016 7040 12032 7104
rect 12096 7040 12112 7104
rect 12176 7040 12192 7104
rect 12256 7040 12264 7104
rect 11944 6016 12264 7040
rect 11944 5952 11952 6016
rect 12016 5952 12032 6016
rect 12096 5952 12112 6016
rect 12176 5952 12192 6016
rect 12256 5952 12264 6016
rect 11944 4928 12264 5952
rect 11944 4864 11952 4928
rect 12016 4864 12032 4928
rect 12096 4864 12112 4928
rect 12176 4864 12192 4928
rect 12256 4864 12264 4928
rect 11944 3840 12264 4864
rect 11944 3776 11952 3840
rect 12016 3776 12032 3840
rect 12096 3776 12112 3840
rect 12176 3776 12192 3840
rect 12256 3776 12264 3840
rect 11944 3294 12264 3776
rect 11944 3058 11986 3294
rect 12222 3058 12264 3294
rect 11944 2752 12264 3058
rect 11944 2688 11952 2752
rect 12016 2688 12032 2752
rect 12096 2688 12112 2752
rect 12176 2688 12192 2752
rect 12256 2688 12264 2752
rect 11944 2128 12264 2688
rect 12604 69664 12924 69680
rect 12604 69600 12612 69664
rect 12676 69600 12692 69664
rect 12756 69600 12772 69664
rect 12836 69600 12852 69664
rect 12916 69600 12924 69664
rect 12604 68954 12924 69600
rect 12604 68718 12646 68954
rect 12882 68718 12924 68954
rect 12604 68576 12924 68718
rect 12604 68512 12612 68576
rect 12676 68512 12692 68576
rect 12756 68512 12772 68576
rect 12836 68512 12852 68576
rect 12916 68512 12924 68576
rect 12604 67488 12924 68512
rect 12604 67424 12612 67488
rect 12676 67424 12692 67488
rect 12756 67424 12772 67488
rect 12836 67424 12852 67488
rect 12916 67424 12924 67488
rect 12604 66400 12924 67424
rect 12604 66336 12612 66400
rect 12676 66336 12692 66400
rect 12756 66336 12772 66400
rect 12836 66336 12852 66400
rect 12916 66336 12924 66400
rect 12604 65312 12924 66336
rect 12604 65248 12612 65312
rect 12676 65248 12692 65312
rect 12756 65248 12772 65312
rect 12836 65248 12852 65312
rect 12916 65248 12924 65312
rect 12604 64224 12924 65248
rect 12604 64160 12612 64224
rect 12676 64160 12692 64224
rect 12756 64160 12772 64224
rect 12836 64160 12852 64224
rect 12916 64160 12924 64224
rect 12604 63954 12924 64160
rect 12604 63718 12646 63954
rect 12882 63718 12924 63954
rect 12604 63136 12924 63718
rect 12604 63072 12612 63136
rect 12676 63072 12692 63136
rect 12756 63072 12772 63136
rect 12836 63072 12852 63136
rect 12916 63072 12924 63136
rect 12604 62048 12924 63072
rect 12604 61984 12612 62048
rect 12676 61984 12692 62048
rect 12756 61984 12772 62048
rect 12836 61984 12852 62048
rect 12916 61984 12924 62048
rect 12604 60960 12924 61984
rect 12604 60896 12612 60960
rect 12676 60896 12692 60960
rect 12756 60896 12772 60960
rect 12836 60896 12852 60960
rect 12916 60896 12924 60960
rect 12604 59872 12924 60896
rect 12604 59808 12612 59872
rect 12676 59808 12692 59872
rect 12756 59808 12772 59872
rect 12836 59808 12852 59872
rect 12916 59808 12924 59872
rect 12604 58954 12924 59808
rect 12604 58784 12646 58954
rect 12882 58784 12924 58954
rect 12604 58720 12612 58784
rect 12916 58720 12924 58784
rect 12604 58718 12646 58720
rect 12882 58718 12924 58720
rect 12604 57696 12924 58718
rect 12604 57632 12612 57696
rect 12676 57632 12692 57696
rect 12756 57632 12772 57696
rect 12836 57632 12852 57696
rect 12916 57632 12924 57696
rect 12604 56608 12924 57632
rect 12604 56544 12612 56608
rect 12676 56544 12692 56608
rect 12756 56544 12772 56608
rect 12836 56544 12852 56608
rect 12916 56544 12924 56608
rect 12604 55520 12924 56544
rect 12604 55456 12612 55520
rect 12676 55456 12692 55520
rect 12756 55456 12772 55520
rect 12836 55456 12852 55520
rect 12916 55456 12924 55520
rect 12604 54432 12924 55456
rect 12604 54368 12612 54432
rect 12676 54368 12692 54432
rect 12756 54368 12772 54432
rect 12836 54368 12852 54432
rect 12916 54368 12924 54432
rect 12604 53954 12924 54368
rect 12604 53718 12646 53954
rect 12882 53718 12924 53954
rect 12604 53344 12924 53718
rect 12604 53280 12612 53344
rect 12676 53280 12692 53344
rect 12756 53280 12772 53344
rect 12836 53280 12852 53344
rect 12916 53280 12924 53344
rect 12604 52256 12924 53280
rect 12604 52192 12612 52256
rect 12676 52192 12692 52256
rect 12756 52192 12772 52256
rect 12836 52192 12852 52256
rect 12916 52192 12924 52256
rect 12604 51168 12924 52192
rect 12604 51104 12612 51168
rect 12676 51104 12692 51168
rect 12756 51104 12772 51168
rect 12836 51104 12852 51168
rect 12916 51104 12924 51168
rect 12604 50080 12924 51104
rect 12604 50016 12612 50080
rect 12676 50016 12692 50080
rect 12756 50016 12772 50080
rect 12836 50016 12852 50080
rect 12916 50016 12924 50080
rect 12604 48992 12924 50016
rect 12604 48928 12612 48992
rect 12676 48954 12692 48992
rect 12756 48954 12772 48992
rect 12836 48954 12852 48992
rect 12916 48928 12924 48992
rect 12604 48718 12646 48928
rect 12882 48718 12924 48928
rect 12604 47904 12924 48718
rect 12604 47840 12612 47904
rect 12676 47840 12692 47904
rect 12756 47840 12772 47904
rect 12836 47840 12852 47904
rect 12916 47840 12924 47904
rect 12604 46816 12924 47840
rect 12604 46752 12612 46816
rect 12676 46752 12692 46816
rect 12756 46752 12772 46816
rect 12836 46752 12852 46816
rect 12916 46752 12924 46816
rect 12604 45728 12924 46752
rect 12604 45664 12612 45728
rect 12676 45664 12692 45728
rect 12756 45664 12772 45728
rect 12836 45664 12852 45728
rect 12916 45664 12924 45728
rect 12604 44640 12924 45664
rect 12604 44576 12612 44640
rect 12676 44576 12692 44640
rect 12756 44576 12772 44640
rect 12836 44576 12852 44640
rect 12916 44576 12924 44640
rect 12604 43954 12924 44576
rect 12604 43718 12646 43954
rect 12882 43718 12924 43954
rect 12604 43552 12924 43718
rect 12604 43488 12612 43552
rect 12676 43488 12692 43552
rect 12756 43488 12772 43552
rect 12836 43488 12852 43552
rect 12916 43488 12924 43552
rect 12604 42464 12924 43488
rect 12604 42400 12612 42464
rect 12676 42400 12692 42464
rect 12756 42400 12772 42464
rect 12836 42400 12852 42464
rect 12916 42400 12924 42464
rect 12604 41376 12924 42400
rect 12604 41312 12612 41376
rect 12676 41312 12692 41376
rect 12756 41312 12772 41376
rect 12836 41312 12852 41376
rect 12916 41312 12924 41376
rect 12604 40288 12924 41312
rect 12604 40224 12612 40288
rect 12676 40224 12692 40288
rect 12756 40224 12772 40288
rect 12836 40224 12852 40288
rect 12916 40224 12924 40288
rect 12604 39200 12924 40224
rect 12604 39136 12612 39200
rect 12676 39136 12692 39200
rect 12756 39136 12772 39200
rect 12836 39136 12852 39200
rect 12916 39136 12924 39200
rect 12604 38954 12924 39136
rect 12604 38718 12646 38954
rect 12882 38718 12924 38954
rect 12604 38112 12924 38718
rect 12604 38048 12612 38112
rect 12676 38048 12692 38112
rect 12756 38048 12772 38112
rect 12836 38048 12852 38112
rect 12916 38048 12924 38112
rect 12604 37024 12924 38048
rect 12604 36960 12612 37024
rect 12676 36960 12692 37024
rect 12756 36960 12772 37024
rect 12836 36960 12852 37024
rect 12916 36960 12924 37024
rect 12604 35936 12924 36960
rect 12604 35872 12612 35936
rect 12676 35872 12692 35936
rect 12756 35872 12772 35936
rect 12836 35872 12852 35936
rect 12916 35872 12924 35936
rect 12604 34848 12924 35872
rect 12604 34784 12612 34848
rect 12676 34784 12692 34848
rect 12756 34784 12772 34848
rect 12836 34784 12852 34848
rect 12916 34784 12924 34848
rect 12604 33954 12924 34784
rect 12604 33760 12646 33954
rect 12882 33760 12924 33954
rect 12604 33696 12612 33760
rect 12676 33696 12692 33718
rect 12756 33696 12772 33718
rect 12836 33696 12852 33718
rect 12916 33696 12924 33760
rect 12604 32672 12924 33696
rect 12604 32608 12612 32672
rect 12676 32608 12692 32672
rect 12756 32608 12772 32672
rect 12836 32608 12852 32672
rect 12916 32608 12924 32672
rect 12604 31584 12924 32608
rect 12604 31520 12612 31584
rect 12676 31520 12692 31584
rect 12756 31520 12772 31584
rect 12836 31520 12852 31584
rect 12916 31520 12924 31584
rect 12604 30496 12924 31520
rect 12604 30432 12612 30496
rect 12676 30432 12692 30496
rect 12756 30432 12772 30496
rect 12836 30432 12852 30496
rect 12916 30432 12924 30496
rect 12604 29408 12924 30432
rect 12604 29344 12612 29408
rect 12676 29344 12692 29408
rect 12756 29344 12772 29408
rect 12836 29344 12852 29408
rect 12916 29344 12924 29408
rect 12604 28954 12924 29344
rect 12604 28718 12646 28954
rect 12882 28718 12924 28954
rect 12604 28320 12924 28718
rect 12604 28256 12612 28320
rect 12676 28256 12692 28320
rect 12756 28256 12772 28320
rect 12836 28256 12852 28320
rect 12916 28256 12924 28320
rect 12604 27232 12924 28256
rect 12604 27168 12612 27232
rect 12676 27168 12692 27232
rect 12756 27168 12772 27232
rect 12836 27168 12852 27232
rect 12916 27168 12924 27232
rect 12604 26144 12924 27168
rect 12604 26080 12612 26144
rect 12676 26080 12692 26144
rect 12756 26080 12772 26144
rect 12836 26080 12852 26144
rect 12916 26080 12924 26144
rect 12604 25056 12924 26080
rect 12604 24992 12612 25056
rect 12676 24992 12692 25056
rect 12756 24992 12772 25056
rect 12836 24992 12852 25056
rect 12916 24992 12924 25056
rect 12604 23968 12924 24992
rect 12604 23904 12612 23968
rect 12676 23954 12692 23968
rect 12756 23954 12772 23968
rect 12836 23954 12852 23968
rect 12916 23904 12924 23968
rect 12604 23718 12646 23904
rect 12882 23718 12924 23904
rect 12604 22880 12924 23718
rect 12604 22816 12612 22880
rect 12676 22816 12692 22880
rect 12756 22816 12772 22880
rect 12836 22816 12852 22880
rect 12916 22816 12924 22880
rect 12604 21792 12924 22816
rect 12604 21728 12612 21792
rect 12676 21728 12692 21792
rect 12756 21728 12772 21792
rect 12836 21728 12852 21792
rect 12916 21728 12924 21792
rect 12604 20704 12924 21728
rect 12604 20640 12612 20704
rect 12676 20640 12692 20704
rect 12756 20640 12772 20704
rect 12836 20640 12852 20704
rect 12916 20640 12924 20704
rect 12604 19616 12924 20640
rect 12604 19552 12612 19616
rect 12676 19552 12692 19616
rect 12756 19552 12772 19616
rect 12836 19552 12852 19616
rect 12916 19552 12924 19616
rect 12604 18954 12924 19552
rect 12604 18718 12646 18954
rect 12882 18718 12924 18954
rect 12604 18528 12924 18718
rect 12604 18464 12612 18528
rect 12676 18464 12692 18528
rect 12756 18464 12772 18528
rect 12836 18464 12852 18528
rect 12916 18464 12924 18528
rect 12604 17440 12924 18464
rect 12604 17376 12612 17440
rect 12676 17376 12692 17440
rect 12756 17376 12772 17440
rect 12836 17376 12852 17440
rect 12916 17376 12924 17440
rect 12604 16352 12924 17376
rect 12604 16288 12612 16352
rect 12676 16288 12692 16352
rect 12756 16288 12772 16352
rect 12836 16288 12852 16352
rect 12916 16288 12924 16352
rect 12604 15264 12924 16288
rect 12604 15200 12612 15264
rect 12676 15200 12692 15264
rect 12756 15200 12772 15264
rect 12836 15200 12852 15264
rect 12916 15200 12924 15264
rect 12604 14176 12924 15200
rect 12604 14112 12612 14176
rect 12676 14112 12692 14176
rect 12756 14112 12772 14176
rect 12836 14112 12852 14176
rect 12916 14112 12924 14176
rect 12604 13954 12924 14112
rect 12604 13718 12646 13954
rect 12882 13718 12924 13954
rect 12604 13088 12924 13718
rect 12604 13024 12612 13088
rect 12676 13024 12692 13088
rect 12756 13024 12772 13088
rect 12836 13024 12852 13088
rect 12916 13024 12924 13088
rect 12604 12000 12924 13024
rect 12604 11936 12612 12000
rect 12676 11936 12692 12000
rect 12756 11936 12772 12000
rect 12836 11936 12852 12000
rect 12916 11936 12924 12000
rect 12604 10912 12924 11936
rect 12604 10848 12612 10912
rect 12676 10848 12692 10912
rect 12756 10848 12772 10912
rect 12836 10848 12852 10912
rect 12916 10848 12924 10912
rect 12604 9824 12924 10848
rect 12604 9760 12612 9824
rect 12676 9760 12692 9824
rect 12756 9760 12772 9824
rect 12836 9760 12852 9824
rect 12916 9760 12924 9824
rect 12604 8954 12924 9760
rect 12604 8736 12646 8954
rect 12882 8736 12924 8954
rect 12604 8672 12612 8736
rect 12676 8672 12692 8718
rect 12756 8672 12772 8718
rect 12836 8672 12852 8718
rect 12916 8672 12924 8736
rect 12604 7648 12924 8672
rect 12604 7584 12612 7648
rect 12676 7584 12692 7648
rect 12756 7584 12772 7648
rect 12836 7584 12852 7648
rect 12916 7584 12924 7648
rect 12604 6560 12924 7584
rect 12604 6496 12612 6560
rect 12676 6496 12692 6560
rect 12756 6496 12772 6560
rect 12836 6496 12852 6560
rect 12916 6496 12924 6560
rect 12604 5472 12924 6496
rect 12604 5408 12612 5472
rect 12676 5408 12692 5472
rect 12756 5408 12772 5472
rect 12836 5408 12852 5472
rect 12916 5408 12924 5472
rect 12604 4384 12924 5408
rect 12604 4320 12612 4384
rect 12676 4320 12692 4384
rect 12756 4320 12772 4384
rect 12836 4320 12852 4384
rect 12916 4320 12924 4384
rect 12604 3954 12924 4320
rect 12604 3718 12646 3954
rect 12882 3718 12924 3954
rect 12604 3296 12924 3718
rect 12604 3232 12612 3296
rect 12676 3232 12692 3296
rect 12756 3232 12772 3296
rect 12836 3232 12852 3296
rect 12916 3232 12924 3296
rect 12604 2208 12924 3232
rect 12604 2144 12612 2208
rect 12676 2144 12692 2208
rect 12756 2144 12772 2208
rect 12836 2144 12852 2208
rect 12916 2144 12924 2208
rect 12604 2128 12924 2144
rect 16944 69120 17264 69680
rect 16944 69056 16952 69120
rect 17016 69056 17032 69120
rect 17096 69056 17112 69120
rect 17176 69056 17192 69120
rect 17256 69056 17264 69120
rect 16944 68294 17264 69056
rect 16944 68058 16986 68294
rect 17222 68058 17264 68294
rect 16944 68032 17264 68058
rect 16944 67968 16952 68032
rect 17016 67968 17032 68032
rect 17096 67968 17112 68032
rect 17176 67968 17192 68032
rect 17256 67968 17264 68032
rect 16944 66944 17264 67968
rect 16944 66880 16952 66944
rect 17016 66880 17032 66944
rect 17096 66880 17112 66944
rect 17176 66880 17192 66944
rect 17256 66880 17264 66944
rect 16944 65856 17264 66880
rect 16944 65792 16952 65856
rect 17016 65792 17032 65856
rect 17096 65792 17112 65856
rect 17176 65792 17192 65856
rect 17256 65792 17264 65856
rect 16944 64768 17264 65792
rect 16944 64704 16952 64768
rect 17016 64704 17032 64768
rect 17096 64704 17112 64768
rect 17176 64704 17192 64768
rect 17256 64704 17264 64768
rect 16944 63680 17264 64704
rect 16944 63616 16952 63680
rect 17016 63616 17032 63680
rect 17096 63616 17112 63680
rect 17176 63616 17192 63680
rect 17256 63616 17264 63680
rect 16944 63294 17264 63616
rect 16944 63058 16986 63294
rect 17222 63058 17264 63294
rect 16944 62592 17264 63058
rect 16944 62528 16952 62592
rect 17016 62528 17032 62592
rect 17096 62528 17112 62592
rect 17176 62528 17192 62592
rect 17256 62528 17264 62592
rect 16944 61504 17264 62528
rect 16944 61440 16952 61504
rect 17016 61440 17032 61504
rect 17096 61440 17112 61504
rect 17176 61440 17192 61504
rect 17256 61440 17264 61504
rect 16944 60416 17264 61440
rect 16944 60352 16952 60416
rect 17016 60352 17032 60416
rect 17096 60352 17112 60416
rect 17176 60352 17192 60416
rect 17256 60352 17264 60416
rect 16944 59328 17264 60352
rect 16944 59264 16952 59328
rect 17016 59264 17032 59328
rect 17096 59264 17112 59328
rect 17176 59264 17192 59328
rect 17256 59264 17264 59328
rect 16944 58294 17264 59264
rect 16944 58240 16986 58294
rect 17222 58240 17264 58294
rect 16944 58176 16952 58240
rect 17256 58176 17264 58240
rect 16944 58058 16986 58176
rect 17222 58058 17264 58176
rect 16944 57152 17264 58058
rect 16944 57088 16952 57152
rect 17016 57088 17032 57152
rect 17096 57088 17112 57152
rect 17176 57088 17192 57152
rect 17256 57088 17264 57152
rect 16944 56064 17264 57088
rect 16944 56000 16952 56064
rect 17016 56000 17032 56064
rect 17096 56000 17112 56064
rect 17176 56000 17192 56064
rect 17256 56000 17264 56064
rect 16944 54976 17264 56000
rect 16944 54912 16952 54976
rect 17016 54912 17032 54976
rect 17096 54912 17112 54976
rect 17176 54912 17192 54976
rect 17256 54912 17264 54976
rect 16944 53888 17264 54912
rect 16944 53824 16952 53888
rect 17016 53824 17032 53888
rect 17096 53824 17112 53888
rect 17176 53824 17192 53888
rect 17256 53824 17264 53888
rect 16944 53294 17264 53824
rect 16944 53058 16986 53294
rect 17222 53058 17264 53294
rect 16944 52800 17264 53058
rect 16944 52736 16952 52800
rect 17016 52736 17032 52800
rect 17096 52736 17112 52800
rect 17176 52736 17192 52800
rect 17256 52736 17264 52800
rect 16944 51712 17264 52736
rect 16944 51648 16952 51712
rect 17016 51648 17032 51712
rect 17096 51648 17112 51712
rect 17176 51648 17192 51712
rect 17256 51648 17264 51712
rect 16944 50624 17264 51648
rect 16944 50560 16952 50624
rect 17016 50560 17032 50624
rect 17096 50560 17112 50624
rect 17176 50560 17192 50624
rect 17256 50560 17264 50624
rect 16944 49536 17264 50560
rect 16944 49472 16952 49536
rect 17016 49472 17032 49536
rect 17096 49472 17112 49536
rect 17176 49472 17192 49536
rect 17256 49472 17264 49536
rect 16944 48448 17264 49472
rect 16944 48384 16952 48448
rect 17016 48384 17032 48448
rect 17096 48384 17112 48448
rect 17176 48384 17192 48448
rect 17256 48384 17264 48448
rect 16944 48294 17264 48384
rect 16944 48058 16986 48294
rect 17222 48058 17264 48294
rect 16944 47360 17264 48058
rect 16944 47296 16952 47360
rect 17016 47296 17032 47360
rect 17096 47296 17112 47360
rect 17176 47296 17192 47360
rect 17256 47296 17264 47360
rect 16944 46272 17264 47296
rect 16944 46208 16952 46272
rect 17016 46208 17032 46272
rect 17096 46208 17112 46272
rect 17176 46208 17192 46272
rect 17256 46208 17264 46272
rect 16944 45184 17264 46208
rect 16944 45120 16952 45184
rect 17016 45120 17032 45184
rect 17096 45120 17112 45184
rect 17176 45120 17192 45184
rect 17256 45120 17264 45184
rect 16944 44096 17264 45120
rect 16944 44032 16952 44096
rect 17016 44032 17032 44096
rect 17096 44032 17112 44096
rect 17176 44032 17192 44096
rect 17256 44032 17264 44096
rect 16944 43294 17264 44032
rect 16944 43058 16986 43294
rect 17222 43058 17264 43294
rect 16944 43008 17264 43058
rect 16944 42944 16952 43008
rect 17016 42944 17032 43008
rect 17096 42944 17112 43008
rect 17176 42944 17192 43008
rect 17256 42944 17264 43008
rect 16944 41920 17264 42944
rect 16944 41856 16952 41920
rect 17016 41856 17032 41920
rect 17096 41856 17112 41920
rect 17176 41856 17192 41920
rect 17256 41856 17264 41920
rect 16944 40832 17264 41856
rect 16944 40768 16952 40832
rect 17016 40768 17032 40832
rect 17096 40768 17112 40832
rect 17176 40768 17192 40832
rect 17256 40768 17264 40832
rect 16944 39744 17264 40768
rect 16944 39680 16952 39744
rect 17016 39680 17032 39744
rect 17096 39680 17112 39744
rect 17176 39680 17192 39744
rect 17256 39680 17264 39744
rect 16944 38656 17264 39680
rect 16944 38592 16952 38656
rect 17016 38592 17032 38656
rect 17096 38592 17112 38656
rect 17176 38592 17192 38656
rect 17256 38592 17264 38656
rect 16944 38294 17264 38592
rect 16944 38058 16986 38294
rect 17222 38058 17264 38294
rect 16944 37568 17264 38058
rect 16944 37504 16952 37568
rect 17016 37504 17032 37568
rect 17096 37504 17112 37568
rect 17176 37504 17192 37568
rect 17256 37504 17264 37568
rect 16944 36480 17264 37504
rect 16944 36416 16952 36480
rect 17016 36416 17032 36480
rect 17096 36416 17112 36480
rect 17176 36416 17192 36480
rect 17256 36416 17264 36480
rect 16944 35392 17264 36416
rect 16944 35328 16952 35392
rect 17016 35328 17032 35392
rect 17096 35328 17112 35392
rect 17176 35328 17192 35392
rect 17256 35328 17264 35392
rect 16944 34304 17264 35328
rect 16944 34240 16952 34304
rect 17016 34240 17032 34304
rect 17096 34240 17112 34304
rect 17176 34240 17192 34304
rect 17256 34240 17264 34304
rect 16944 33294 17264 34240
rect 16944 33216 16986 33294
rect 17222 33216 17264 33294
rect 16944 33152 16952 33216
rect 17256 33152 17264 33216
rect 16944 33058 16986 33152
rect 17222 33058 17264 33152
rect 16944 32128 17264 33058
rect 16944 32064 16952 32128
rect 17016 32064 17032 32128
rect 17096 32064 17112 32128
rect 17176 32064 17192 32128
rect 17256 32064 17264 32128
rect 16944 31040 17264 32064
rect 16944 30976 16952 31040
rect 17016 30976 17032 31040
rect 17096 30976 17112 31040
rect 17176 30976 17192 31040
rect 17256 30976 17264 31040
rect 16944 29952 17264 30976
rect 16944 29888 16952 29952
rect 17016 29888 17032 29952
rect 17096 29888 17112 29952
rect 17176 29888 17192 29952
rect 17256 29888 17264 29952
rect 16944 28864 17264 29888
rect 16944 28800 16952 28864
rect 17016 28800 17032 28864
rect 17096 28800 17112 28864
rect 17176 28800 17192 28864
rect 17256 28800 17264 28864
rect 16944 28294 17264 28800
rect 16944 28058 16986 28294
rect 17222 28058 17264 28294
rect 16944 27776 17264 28058
rect 16944 27712 16952 27776
rect 17016 27712 17032 27776
rect 17096 27712 17112 27776
rect 17176 27712 17192 27776
rect 17256 27712 17264 27776
rect 16944 26688 17264 27712
rect 16944 26624 16952 26688
rect 17016 26624 17032 26688
rect 17096 26624 17112 26688
rect 17176 26624 17192 26688
rect 17256 26624 17264 26688
rect 16944 25600 17264 26624
rect 16944 25536 16952 25600
rect 17016 25536 17032 25600
rect 17096 25536 17112 25600
rect 17176 25536 17192 25600
rect 17256 25536 17264 25600
rect 16944 24512 17264 25536
rect 16944 24448 16952 24512
rect 17016 24448 17032 24512
rect 17096 24448 17112 24512
rect 17176 24448 17192 24512
rect 17256 24448 17264 24512
rect 16944 23424 17264 24448
rect 16944 23360 16952 23424
rect 17016 23360 17032 23424
rect 17096 23360 17112 23424
rect 17176 23360 17192 23424
rect 17256 23360 17264 23424
rect 16944 23294 17264 23360
rect 16944 23058 16986 23294
rect 17222 23058 17264 23294
rect 16944 22336 17264 23058
rect 16944 22272 16952 22336
rect 17016 22272 17032 22336
rect 17096 22272 17112 22336
rect 17176 22272 17192 22336
rect 17256 22272 17264 22336
rect 16944 21248 17264 22272
rect 16944 21184 16952 21248
rect 17016 21184 17032 21248
rect 17096 21184 17112 21248
rect 17176 21184 17192 21248
rect 17256 21184 17264 21248
rect 16944 20160 17264 21184
rect 16944 20096 16952 20160
rect 17016 20096 17032 20160
rect 17096 20096 17112 20160
rect 17176 20096 17192 20160
rect 17256 20096 17264 20160
rect 16944 19072 17264 20096
rect 16944 19008 16952 19072
rect 17016 19008 17032 19072
rect 17096 19008 17112 19072
rect 17176 19008 17192 19072
rect 17256 19008 17264 19072
rect 16944 18294 17264 19008
rect 16944 18058 16986 18294
rect 17222 18058 17264 18294
rect 16944 17984 17264 18058
rect 16944 17920 16952 17984
rect 17016 17920 17032 17984
rect 17096 17920 17112 17984
rect 17176 17920 17192 17984
rect 17256 17920 17264 17984
rect 16944 16896 17264 17920
rect 16944 16832 16952 16896
rect 17016 16832 17032 16896
rect 17096 16832 17112 16896
rect 17176 16832 17192 16896
rect 17256 16832 17264 16896
rect 16944 15808 17264 16832
rect 16944 15744 16952 15808
rect 17016 15744 17032 15808
rect 17096 15744 17112 15808
rect 17176 15744 17192 15808
rect 17256 15744 17264 15808
rect 16944 14720 17264 15744
rect 16944 14656 16952 14720
rect 17016 14656 17032 14720
rect 17096 14656 17112 14720
rect 17176 14656 17192 14720
rect 17256 14656 17264 14720
rect 16944 13632 17264 14656
rect 16944 13568 16952 13632
rect 17016 13568 17032 13632
rect 17096 13568 17112 13632
rect 17176 13568 17192 13632
rect 17256 13568 17264 13632
rect 16944 13294 17264 13568
rect 16944 13058 16986 13294
rect 17222 13058 17264 13294
rect 16944 12544 17264 13058
rect 16944 12480 16952 12544
rect 17016 12480 17032 12544
rect 17096 12480 17112 12544
rect 17176 12480 17192 12544
rect 17256 12480 17264 12544
rect 16944 11456 17264 12480
rect 16944 11392 16952 11456
rect 17016 11392 17032 11456
rect 17096 11392 17112 11456
rect 17176 11392 17192 11456
rect 17256 11392 17264 11456
rect 16944 10368 17264 11392
rect 16944 10304 16952 10368
rect 17016 10304 17032 10368
rect 17096 10304 17112 10368
rect 17176 10304 17192 10368
rect 17256 10304 17264 10368
rect 16944 9280 17264 10304
rect 16944 9216 16952 9280
rect 17016 9216 17032 9280
rect 17096 9216 17112 9280
rect 17176 9216 17192 9280
rect 17256 9216 17264 9280
rect 16944 8294 17264 9216
rect 16944 8192 16986 8294
rect 17222 8192 17264 8294
rect 16944 8128 16952 8192
rect 17256 8128 17264 8192
rect 16944 8058 16986 8128
rect 17222 8058 17264 8128
rect 16944 7104 17264 8058
rect 16944 7040 16952 7104
rect 17016 7040 17032 7104
rect 17096 7040 17112 7104
rect 17176 7040 17192 7104
rect 17256 7040 17264 7104
rect 16944 6016 17264 7040
rect 16944 5952 16952 6016
rect 17016 5952 17032 6016
rect 17096 5952 17112 6016
rect 17176 5952 17192 6016
rect 17256 5952 17264 6016
rect 16944 4928 17264 5952
rect 16944 4864 16952 4928
rect 17016 4864 17032 4928
rect 17096 4864 17112 4928
rect 17176 4864 17192 4928
rect 17256 4864 17264 4928
rect 16944 3840 17264 4864
rect 16944 3776 16952 3840
rect 17016 3776 17032 3840
rect 17096 3776 17112 3840
rect 17176 3776 17192 3840
rect 17256 3776 17264 3840
rect 16944 3294 17264 3776
rect 16944 3058 16986 3294
rect 17222 3058 17264 3294
rect 16944 2752 17264 3058
rect 16944 2688 16952 2752
rect 17016 2688 17032 2752
rect 17096 2688 17112 2752
rect 17176 2688 17192 2752
rect 17256 2688 17264 2752
rect 16944 2128 17264 2688
rect 17604 69664 17924 69680
rect 17604 69600 17612 69664
rect 17676 69600 17692 69664
rect 17756 69600 17772 69664
rect 17836 69600 17852 69664
rect 17916 69600 17924 69664
rect 17604 68954 17924 69600
rect 17604 68718 17646 68954
rect 17882 68718 17924 68954
rect 17604 68576 17924 68718
rect 17604 68512 17612 68576
rect 17676 68512 17692 68576
rect 17756 68512 17772 68576
rect 17836 68512 17852 68576
rect 17916 68512 17924 68576
rect 17604 67488 17924 68512
rect 17604 67424 17612 67488
rect 17676 67424 17692 67488
rect 17756 67424 17772 67488
rect 17836 67424 17852 67488
rect 17916 67424 17924 67488
rect 17604 66400 17924 67424
rect 17604 66336 17612 66400
rect 17676 66336 17692 66400
rect 17756 66336 17772 66400
rect 17836 66336 17852 66400
rect 17916 66336 17924 66400
rect 17604 65312 17924 66336
rect 17604 65248 17612 65312
rect 17676 65248 17692 65312
rect 17756 65248 17772 65312
rect 17836 65248 17852 65312
rect 17916 65248 17924 65312
rect 17604 64224 17924 65248
rect 17604 64160 17612 64224
rect 17676 64160 17692 64224
rect 17756 64160 17772 64224
rect 17836 64160 17852 64224
rect 17916 64160 17924 64224
rect 17604 63954 17924 64160
rect 17604 63718 17646 63954
rect 17882 63718 17924 63954
rect 17604 63136 17924 63718
rect 17604 63072 17612 63136
rect 17676 63072 17692 63136
rect 17756 63072 17772 63136
rect 17836 63072 17852 63136
rect 17916 63072 17924 63136
rect 17604 62048 17924 63072
rect 17604 61984 17612 62048
rect 17676 61984 17692 62048
rect 17756 61984 17772 62048
rect 17836 61984 17852 62048
rect 17916 61984 17924 62048
rect 17604 60960 17924 61984
rect 17604 60896 17612 60960
rect 17676 60896 17692 60960
rect 17756 60896 17772 60960
rect 17836 60896 17852 60960
rect 17916 60896 17924 60960
rect 17604 59872 17924 60896
rect 17604 59808 17612 59872
rect 17676 59808 17692 59872
rect 17756 59808 17772 59872
rect 17836 59808 17852 59872
rect 17916 59808 17924 59872
rect 17604 58954 17924 59808
rect 17604 58784 17646 58954
rect 17882 58784 17924 58954
rect 17604 58720 17612 58784
rect 17916 58720 17924 58784
rect 17604 58718 17646 58720
rect 17882 58718 17924 58720
rect 17604 57696 17924 58718
rect 17604 57632 17612 57696
rect 17676 57632 17692 57696
rect 17756 57632 17772 57696
rect 17836 57632 17852 57696
rect 17916 57632 17924 57696
rect 17604 56608 17924 57632
rect 17604 56544 17612 56608
rect 17676 56544 17692 56608
rect 17756 56544 17772 56608
rect 17836 56544 17852 56608
rect 17916 56544 17924 56608
rect 17604 55520 17924 56544
rect 17604 55456 17612 55520
rect 17676 55456 17692 55520
rect 17756 55456 17772 55520
rect 17836 55456 17852 55520
rect 17916 55456 17924 55520
rect 17604 54432 17924 55456
rect 17604 54368 17612 54432
rect 17676 54368 17692 54432
rect 17756 54368 17772 54432
rect 17836 54368 17852 54432
rect 17916 54368 17924 54432
rect 17604 53954 17924 54368
rect 17604 53718 17646 53954
rect 17882 53718 17924 53954
rect 17604 53344 17924 53718
rect 17604 53280 17612 53344
rect 17676 53280 17692 53344
rect 17756 53280 17772 53344
rect 17836 53280 17852 53344
rect 17916 53280 17924 53344
rect 17604 52256 17924 53280
rect 17604 52192 17612 52256
rect 17676 52192 17692 52256
rect 17756 52192 17772 52256
rect 17836 52192 17852 52256
rect 17916 52192 17924 52256
rect 17604 51168 17924 52192
rect 17604 51104 17612 51168
rect 17676 51104 17692 51168
rect 17756 51104 17772 51168
rect 17836 51104 17852 51168
rect 17916 51104 17924 51168
rect 17604 50080 17924 51104
rect 17604 50016 17612 50080
rect 17676 50016 17692 50080
rect 17756 50016 17772 50080
rect 17836 50016 17852 50080
rect 17916 50016 17924 50080
rect 17604 48992 17924 50016
rect 17604 48928 17612 48992
rect 17676 48954 17692 48992
rect 17756 48954 17772 48992
rect 17836 48954 17852 48992
rect 17916 48928 17924 48992
rect 17604 48718 17646 48928
rect 17882 48718 17924 48928
rect 17604 47904 17924 48718
rect 17604 47840 17612 47904
rect 17676 47840 17692 47904
rect 17756 47840 17772 47904
rect 17836 47840 17852 47904
rect 17916 47840 17924 47904
rect 17604 46816 17924 47840
rect 17604 46752 17612 46816
rect 17676 46752 17692 46816
rect 17756 46752 17772 46816
rect 17836 46752 17852 46816
rect 17916 46752 17924 46816
rect 17604 45728 17924 46752
rect 21944 69120 22264 69680
rect 21944 69056 21952 69120
rect 22016 69056 22032 69120
rect 22096 69056 22112 69120
rect 22176 69056 22192 69120
rect 22256 69056 22264 69120
rect 21944 68294 22264 69056
rect 21944 68058 21986 68294
rect 22222 68058 22264 68294
rect 21944 68032 22264 68058
rect 21944 67968 21952 68032
rect 22016 67968 22032 68032
rect 22096 67968 22112 68032
rect 22176 67968 22192 68032
rect 22256 67968 22264 68032
rect 21944 66944 22264 67968
rect 21944 66880 21952 66944
rect 22016 66880 22032 66944
rect 22096 66880 22112 66944
rect 22176 66880 22192 66944
rect 22256 66880 22264 66944
rect 21944 65856 22264 66880
rect 21944 65792 21952 65856
rect 22016 65792 22032 65856
rect 22096 65792 22112 65856
rect 22176 65792 22192 65856
rect 22256 65792 22264 65856
rect 21944 64768 22264 65792
rect 21944 64704 21952 64768
rect 22016 64704 22032 64768
rect 22096 64704 22112 64768
rect 22176 64704 22192 64768
rect 22256 64704 22264 64768
rect 21944 63680 22264 64704
rect 21944 63616 21952 63680
rect 22016 63616 22032 63680
rect 22096 63616 22112 63680
rect 22176 63616 22192 63680
rect 22256 63616 22264 63680
rect 21944 63294 22264 63616
rect 21944 63058 21986 63294
rect 22222 63058 22264 63294
rect 21944 62592 22264 63058
rect 21944 62528 21952 62592
rect 22016 62528 22032 62592
rect 22096 62528 22112 62592
rect 22176 62528 22192 62592
rect 22256 62528 22264 62592
rect 21944 61504 22264 62528
rect 21944 61440 21952 61504
rect 22016 61440 22032 61504
rect 22096 61440 22112 61504
rect 22176 61440 22192 61504
rect 22256 61440 22264 61504
rect 21944 60416 22264 61440
rect 21944 60352 21952 60416
rect 22016 60352 22032 60416
rect 22096 60352 22112 60416
rect 22176 60352 22192 60416
rect 22256 60352 22264 60416
rect 21944 59328 22264 60352
rect 21944 59264 21952 59328
rect 22016 59264 22032 59328
rect 22096 59264 22112 59328
rect 22176 59264 22192 59328
rect 22256 59264 22264 59328
rect 21944 58294 22264 59264
rect 21944 58240 21986 58294
rect 22222 58240 22264 58294
rect 21944 58176 21952 58240
rect 22256 58176 22264 58240
rect 21944 58058 21986 58176
rect 22222 58058 22264 58176
rect 21944 57152 22264 58058
rect 21944 57088 21952 57152
rect 22016 57088 22032 57152
rect 22096 57088 22112 57152
rect 22176 57088 22192 57152
rect 22256 57088 22264 57152
rect 21944 56064 22264 57088
rect 21944 56000 21952 56064
rect 22016 56000 22032 56064
rect 22096 56000 22112 56064
rect 22176 56000 22192 56064
rect 22256 56000 22264 56064
rect 21944 54976 22264 56000
rect 21944 54912 21952 54976
rect 22016 54912 22032 54976
rect 22096 54912 22112 54976
rect 22176 54912 22192 54976
rect 22256 54912 22264 54976
rect 21944 53888 22264 54912
rect 21944 53824 21952 53888
rect 22016 53824 22032 53888
rect 22096 53824 22112 53888
rect 22176 53824 22192 53888
rect 22256 53824 22264 53888
rect 21944 53294 22264 53824
rect 21944 53058 21986 53294
rect 22222 53058 22264 53294
rect 21944 52800 22264 53058
rect 21944 52736 21952 52800
rect 22016 52736 22032 52800
rect 22096 52736 22112 52800
rect 22176 52736 22192 52800
rect 22256 52736 22264 52800
rect 21944 51712 22264 52736
rect 21944 51648 21952 51712
rect 22016 51648 22032 51712
rect 22096 51648 22112 51712
rect 22176 51648 22192 51712
rect 22256 51648 22264 51712
rect 21944 50624 22264 51648
rect 21944 50560 21952 50624
rect 22016 50560 22032 50624
rect 22096 50560 22112 50624
rect 22176 50560 22192 50624
rect 22256 50560 22264 50624
rect 21944 49536 22264 50560
rect 21944 49472 21952 49536
rect 22016 49472 22032 49536
rect 22096 49472 22112 49536
rect 22176 49472 22192 49536
rect 22256 49472 22264 49536
rect 21944 48448 22264 49472
rect 21944 48384 21952 48448
rect 22016 48384 22032 48448
rect 22096 48384 22112 48448
rect 22176 48384 22192 48448
rect 22256 48384 22264 48448
rect 21944 48294 22264 48384
rect 21944 48058 21986 48294
rect 22222 48058 22264 48294
rect 21944 47360 22264 48058
rect 21944 47296 21952 47360
rect 22016 47296 22032 47360
rect 22096 47296 22112 47360
rect 22176 47296 22192 47360
rect 22256 47296 22264 47360
rect 21944 46272 22264 47296
rect 21944 46208 21952 46272
rect 22016 46208 22032 46272
rect 22096 46208 22112 46272
rect 22176 46208 22192 46272
rect 22256 46208 22264 46272
rect 21035 45932 21101 45933
rect 21035 45868 21036 45932
rect 21100 45868 21101 45932
rect 21035 45867 21101 45868
rect 17604 45664 17612 45728
rect 17676 45664 17692 45728
rect 17756 45664 17772 45728
rect 17836 45664 17852 45728
rect 17916 45664 17924 45728
rect 17604 44640 17924 45664
rect 17604 44576 17612 44640
rect 17676 44576 17692 44640
rect 17756 44576 17772 44640
rect 17836 44576 17852 44640
rect 17916 44576 17924 44640
rect 17604 43954 17924 44576
rect 17604 43718 17646 43954
rect 17882 43718 17924 43954
rect 17604 43552 17924 43718
rect 17604 43488 17612 43552
rect 17676 43488 17692 43552
rect 17756 43488 17772 43552
rect 17836 43488 17852 43552
rect 17916 43488 17924 43552
rect 17604 42464 17924 43488
rect 17604 42400 17612 42464
rect 17676 42400 17692 42464
rect 17756 42400 17772 42464
rect 17836 42400 17852 42464
rect 17916 42400 17924 42464
rect 17604 41376 17924 42400
rect 17604 41312 17612 41376
rect 17676 41312 17692 41376
rect 17756 41312 17772 41376
rect 17836 41312 17852 41376
rect 17916 41312 17924 41376
rect 17604 40288 17924 41312
rect 17604 40224 17612 40288
rect 17676 40224 17692 40288
rect 17756 40224 17772 40288
rect 17836 40224 17852 40288
rect 17916 40224 17924 40288
rect 17604 39200 17924 40224
rect 17604 39136 17612 39200
rect 17676 39136 17692 39200
rect 17756 39136 17772 39200
rect 17836 39136 17852 39200
rect 17916 39136 17924 39200
rect 17604 38954 17924 39136
rect 17604 38718 17646 38954
rect 17882 38718 17924 38954
rect 17604 38112 17924 38718
rect 17604 38048 17612 38112
rect 17676 38048 17692 38112
rect 17756 38048 17772 38112
rect 17836 38048 17852 38112
rect 17916 38048 17924 38112
rect 17604 37024 17924 38048
rect 17604 36960 17612 37024
rect 17676 36960 17692 37024
rect 17756 36960 17772 37024
rect 17836 36960 17852 37024
rect 17916 36960 17924 37024
rect 17604 35936 17924 36960
rect 18091 36140 18157 36141
rect 18091 36076 18092 36140
rect 18156 36076 18157 36140
rect 18091 36075 18157 36076
rect 17604 35872 17612 35936
rect 17676 35872 17692 35936
rect 17756 35872 17772 35936
rect 17836 35872 17852 35936
rect 17916 35872 17924 35936
rect 17604 34848 17924 35872
rect 17604 34784 17612 34848
rect 17676 34784 17692 34848
rect 17756 34784 17772 34848
rect 17836 34784 17852 34848
rect 17916 34784 17924 34848
rect 17604 33954 17924 34784
rect 18094 34509 18154 36075
rect 18091 34508 18157 34509
rect 18091 34444 18092 34508
rect 18156 34444 18157 34508
rect 18091 34443 18157 34444
rect 17604 33760 17646 33954
rect 17882 33760 17924 33954
rect 21038 33829 21098 45867
rect 21944 45184 22264 46208
rect 21944 45120 21952 45184
rect 22016 45120 22032 45184
rect 22096 45120 22112 45184
rect 22176 45120 22192 45184
rect 22256 45120 22264 45184
rect 21944 44096 22264 45120
rect 21944 44032 21952 44096
rect 22016 44032 22032 44096
rect 22096 44032 22112 44096
rect 22176 44032 22192 44096
rect 22256 44032 22264 44096
rect 21944 43294 22264 44032
rect 21944 43058 21986 43294
rect 22222 43058 22264 43294
rect 21944 43008 22264 43058
rect 21944 42944 21952 43008
rect 22016 42944 22032 43008
rect 22096 42944 22112 43008
rect 22176 42944 22192 43008
rect 22256 42944 22264 43008
rect 21944 41920 22264 42944
rect 21944 41856 21952 41920
rect 22016 41856 22032 41920
rect 22096 41856 22112 41920
rect 22176 41856 22192 41920
rect 22256 41856 22264 41920
rect 21944 40832 22264 41856
rect 21944 40768 21952 40832
rect 22016 40768 22032 40832
rect 22096 40768 22112 40832
rect 22176 40768 22192 40832
rect 22256 40768 22264 40832
rect 21944 39744 22264 40768
rect 21944 39680 21952 39744
rect 22016 39680 22032 39744
rect 22096 39680 22112 39744
rect 22176 39680 22192 39744
rect 22256 39680 22264 39744
rect 21944 38656 22264 39680
rect 21944 38592 21952 38656
rect 22016 38592 22032 38656
rect 22096 38592 22112 38656
rect 22176 38592 22192 38656
rect 22256 38592 22264 38656
rect 21944 38294 22264 38592
rect 21944 38058 21986 38294
rect 22222 38058 22264 38294
rect 21944 37568 22264 38058
rect 21944 37504 21952 37568
rect 22016 37504 22032 37568
rect 22096 37504 22112 37568
rect 22176 37504 22192 37568
rect 22256 37504 22264 37568
rect 21944 36480 22264 37504
rect 21944 36416 21952 36480
rect 22016 36416 22032 36480
rect 22096 36416 22112 36480
rect 22176 36416 22192 36480
rect 22256 36416 22264 36480
rect 21944 35392 22264 36416
rect 21944 35328 21952 35392
rect 22016 35328 22032 35392
rect 22096 35328 22112 35392
rect 22176 35328 22192 35392
rect 22256 35328 22264 35392
rect 21944 34304 22264 35328
rect 21944 34240 21952 34304
rect 22016 34240 22032 34304
rect 22096 34240 22112 34304
rect 22176 34240 22192 34304
rect 22256 34240 22264 34304
rect 21035 33828 21101 33829
rect 21035 33764 21036 33828
rect 21100 33764 21101 33828
rect 21035 33763 21101 33764
rect 17604 33696 17612 33760
rect 17676 33696 17692 33718
rect 17756 33696 17772 33718
rect 17836 33696 17852 33718
rect 17916 33696 17924 33760
rect 17604 32672 17924 33696
rect 17604 32608 17612 32672
rect 17676 32608 17692 32672
rect 17756 32608 17772 32672
rect 17836 32608 17852 32672
rect 17916 32608 17924 32672
rect 17604 31584 17924 32608
rect 17604 31520 17612 31584
rect 17676 31520 17692 31584
rect 17756 31520 17772 31584
rect 17836 31520 17852 31584
rect 17916 31520 17924 31584
rect 17604 30496 17924 31520
rect 17604 30432 17612 30496
rect 17676 30432 17692 30496
rect 17756 30432 17772 30496
rect 17836 30432 17852 30496
rect 17916 30432 17924 30496
rect 17604 29408 17924 30432
rect 17604 29344 17612 29408
rect 17676 29344 17692 29408
rect 17756 29344 17772 29408
rect 17836 29344 17852 29408
rect 17916 29344 17924 29408
rect 17604 28954 17924 29344
rect 17604 28718 17646 28954
rect 17882 28718 17924 28954
rect 17604 28320 17924 28718
rect 17604 28256 17612 28320
rect 17676 28256 17692 28320
rect 17756 28256 17772 28320
rect 17836 28256 17852 28320
rect 17916 28256 17924 28320
rect 17604 27232 17924 28256
rect 17604 27168 17612 27232
rect 17676 27168 17692 27232
rect 17756 27168 17772 27232
rect 17836 27168 17852 27232
rect 17916 27168 17924 27232
rect 17604 26144 17924 27168
rect 17604 26080 17612 26144
rect 17676 26080 17692 26144
rect 17756 26080 17772 26144
rect 17836 26080 17852 26144
rect 17916 26080 17924 26144
rect 17604 25056 17924 26080
rect 17604 24992 17612 25056
rect 17676 24992 17692 25056
rect 17756 24992 17772 25056
rect 17836 24992 17852 25056
rect 17916 24992 17924 25056
rect 17604 23968 17924 24992
rect 17604 23904 17612 23968
rect 17676 23954 17692 23968
rect 17756 23954 17772 23968
rect 17836 23954 17852 23968
rect 17916 23904 17924 23968
rect 17604 23718 17646 23904
rect 17882 23718 17924 23904
rect 17604 22880 17924 23718
rect 17604 22816 17612 22880
rect 17676 22816 17692 22880
rect 17756 22816 17772 22880
rect 17836 22816 17852 22880
rect 17916 22816 17924 22880
rect 17604 21792 17924 22816
rect 21038 22677 21098 33763
rect 21944 33294 22264 34240
rect 21944 33216 21986 33294
rect 22222 33216 22264 33294
rect 21944 33152 21952 33216
rect 22256 33152 22264 33216
rect 21944 33058 21986 33152
rect 22222 33058 22264 33152
rect 21944 32128 22264 33058
rect 21944 32064 21952 32128
rect 22016 32064 22032 32128
rect 22096 32064 22112 32128
rect 22176 32064 22192 32128
rect 22256 32064 22264 32128
rect 21944 31040 22264 32064
rect 21944 30976 21952 31040
rect 22016 30976 22032 31040
rect 22096 30976 22112 31040
rect 22176 30976 22192 31040
rect 22256 30976 22264 31040
rect 21944 29952 22264 30976
rect 21944 29888 21952 29952
rect 22016 29888 22032 29952
rect 22096 29888 22112 29952
rect 22176 29888 22192 29952
rect 22256 29888 22264 29952
rect 21944 28864 22264 29888
rect 21944 28800 21952 28864
rect 22016 28800 22032 28864
rect 22096 28800 22112 28864
rect 22176 28800 22192 28864
rect 22256 28800 22264 28864
rect 21944 28294 22264 28800
rect 21944 28058 21986 28294
rect 22222 28058 22264 28294
rect 21944 27776 22264 28058
rect 21944 27712 21952 27776
rect 22016 27712 22032 27776
rect 22096 27712 22112 27776
rect 22176 27712 22192 27776
rect 22256 27712 22264 27776
rect 21944 26688 22264 27712
rect 21944 26624 21952 26688
rect 22016 26624 22032 26688
rect 22096 26624 22112 26688
rect 22176 26624 22192 26688
rect 22256 26624 22264 26688
rect 21944 25600 22264 26624
rect 21944 25536 21952 25600
rect 22016 25536 22032 25600
rect 22096 25536 22112 25600
rect 22176 25536 22192 25600
rect 22256 25536 22264 25600
rect 21944 24512 22264 25536
rect 21944 24448 21952 24512
rect 22016 24448 22032 24512
rect 22096 24448 22112 24512
rect 22176 24448 22192 24512
rect 22256 24448 22264 24512
rect 21944 23424 22264 24448
rect 21944 23360 21952 23424
rect 22016 23360 22032 23424
rect 22096 23360 22112 23424
rect 22176 23360 22192 23424
rect 22256 23360 22264 23424
rect 21944 23294 22264 23360
rect 21944 23058 21986 23294
rect 22222 23058 22264 23294
rect 21035 22676 21101 22677
rect 21035 22612 21036 22676
rect 21100 22612 21101 22676
rect 21035 22611 21101 22612
rect 21038 21997 21098 22611
rect 21944 22336 22264 23058
rect 21944 22272 21952 22336
rect 22016 22272 22032 22336
rect 22096 22272 22112 22336
rect 22176 22272 22192 22336
rect 22256 22272 22264 22336
rect 21035 21996 21101 21997
rect 21035 21932 21036 21996
rect 21100 21932 21101 21996
rect 21035 21931 21101 21932
rect 17604 21728 17612 21792
rect 17676 21728 17692 21792
rect 17756 21728 17772 21792
rect 17836 21728 17852 21792
rect 17916 21728 17924 21792
rect 17604 20704 17924 21728
rect 17604 20640 17612 20704
rect 17676 20640 17692 20704
rect 17756 20640 17772 20704
rect 17836 20640 17852 20704
rect 17916 20640 17924 20704
rect 17604 19616 17924 20640
rect 17604 19552 17612 19616
rect 17676 19552 17692 19616
rect 17756 19552 17772 19616
rect 17836 19552 17852 19616
rect 17916 19552 17924 19616
rect 17604 18954 17924 19552
rect 17604 18718 17646 18954
rect 17882 18718 17924 18954
rect 17604 18528 17924 18718
rect 17604 18464 17612 18528
rect 17676 18464 17692 18528
rect 17756 18464 17772 18528
rect 17836 18464 17852 18528
rect 17916 18464 17924 18528
rect 17604 17440 17924 18464
rect 17604 17376 17612 17440
rect 17676 17376 17692 17440
rect 17756 17376 17772 17440
rect 17836 17376 17852 17440
rect 17916 17376 17924 17440
rect 17604 16352 17924 17376
rect 17604 16288 17612 16352
rect 17676 16288 17692 16352
rect 17756 16288 17772 16352
rect 17836 16288 17852 16352
rect 17916 16288 17924 16352
rect 17604 15264 17924 16288
rect 17604 15200 17612 15264
rect 17676 15200 17692 15264
rect 17756 15200 17772 15264
rect 17836 15200 17852 15264
rect 17916 15200 17924 15264
rect 17604 14176 17924 15200
rect 17604 14112 17612 14176
rect 17676 14112 17692 14176
rect 17756 14112 17772 14176
rect 17836 14112 17852 14176
rect 17916 14112 17924 14176
rect 17604 13954 17924 14112
rect 17604 13718 17646 13954
rect 17882 13718 17924 13954
rect 17604 13088 17924 13718
rect 17604 13024 17612 13088
rect 17676 13024 17692 13088
rect 17756 13024 17772 13088
rect 17836 13024 17852 13088
rect 17916 13024 17924 13088
rect 17604 12000 17924 13024
rect 17604 11936 17612 12000
rect 17676 11936 17692 12000
rect 17756 11936 17772 12000
rect 17836 11936 17852 12000
rect 17916 11936 17924 12000
rect 17604 10912 17924 11936
rect 17604 10848 17612 10912
rect 17676 10848 17692 10912
rect 17756 10848 17772 10912
rect 17836 10848 17852 10912
rect 17916 10848 17924 10912
rect 17604 9824 17924 10848
rect 17604 9760 17612 9824
rect 17676 9760 17692 9824
rect 17756 9760 17772 9824
rect 17836 9760 17852 9824
rect 17916 9760 17924 9824
rect 17604 8954 17924 9760
rect 17604 8736 17646 8954
rect 17882 8736 17924 8954
rect 17604 8672 17612 8736
rect 17676 8672 17692 8718
rect 17756 8672 17772 8718
rect 17836 8672 17852 8718
rect 17916 8672 17924 8736
rect 17604 7648 17924 8672
rect 17604 7584 17612 7648
rect 17676 7584 17692 7648
rect 17756 7584 17772 7648
rect 17836 7584 17852 7648
rect 17916 7584 17924 7648
rect 17604 6560 17924 7584
rect 17604 6496 17612 6560
rect 17676 6496 17692 6560
rect 17756 6496 17772 6560
rect 17836 6496 17852 6560
rect 17916 6496 17924 6560
rect 17604 5472 17924 6496
rect 17604 5408 17612 5472
rect 17676 5408 17692 5472
rect 17756 5408 17772 5472
rect 17836 5408 17852 5472
rect 17916 5408 17924 5472
rect 17604 4384 17924 5408
rect 17604 4320 17612 4384
rect 17676 4320 17692 4384
rect 17756 4320 17772 4384
rect 17836 4320 17852 4384
rect 17916 4320 17924 4384
rect 17604 3954 17924 4320
rect 17604 3718 17646 3954
rect 17882 3718 17924 3954
rect 17604 3296 17924 3718
rect 17604 3232 17612 3296
rect 17676 3232 17692 3296
rect 17756 3232 17772 3296
rect 17836 3232 17852 3296
rect 17916 3232 17924 3296
rect 17604 2208 17924 3232
rect 17604 2144 17612 2208
rect 17676 2144 17692 2208
rect 17756 2144 17772 2208
rect 17836 2144 17852 2208
rect 17916 2144 17924 2208
rect 17604 2128 17924 2144
rect 21944 21248 22264 22272
rect 21944 21184 21952 21248
rect 22016 21184 22032 21248
rect 22096 21184 22112 21248
rect 22176 21184 22192 21248
rect 22256 21184 22264 21248
rect 21944 20160 22264 21184
rect 21944 20096 21952 20160
rect 22016 20096 22032 20160
rect 22096 20096 22112 20160
rect 22176 20096 22192 20160
rect 22256 20096 22264 20160
rect 21944 19072 22264 20096
rect 21944 19008 21952 19072
rect 22016 19008 22032 19072
rect 22096 19008 22112 19072
rect 22176 19008 22192 19072
rect 22256 19008 22264 19072
rect 21944 18294 22264 19008
rect 21944 18058 21986 18294
rect 22222 18058 22264 18294
rect 21944 17984 22264 18058
rect 21944 17920 21952 17984
rect 22016 17920 22032 17984
rect 22096 17920 22112 17984
rect 22176 17920 22192 17984
rect 22256 17920 22264 17984
rect 21944 16896 22264 17920
rect 21944 16832 21952 16896
rect 22016 16832 22032 16896
rect 22096 16832 22112 16896
rect 22176 16832 22192 16896
rect 22256 16832 22264 16896
rect 21944 15808 22264 16832
rect 21944 15744 21952 15808
rect 22016 15744 22032 15808
rect 22096 15744 22112 15808
rect 22176 15744 22192 15808
rect 22256 15744 22264 15808
rect 21944 14720 22264 15744
rect 21944 14656 21952 14720
rect 22016 14656 22032 14720
rect 22096 14656 22112 14720
rect 22176 14656 22192 14720
rect 22256 14656 22264 14720
rect 21944 13632 22264 14656
rect 21944 13568 21952 13632
rect 22016 13568 22032 13632
rect 22096 13568 22112 13632
rect 22176 13568 22192 13632
rect 22256 13568 22264 13632
rect 21944 13294 22264 13568
rect 21944 13058 21986 13294
rect 22222 13058 22264 13294
rect 21944 12544 22264 13058
rect 21944 12480 21952 12544
rect 22016 12480 22032 12544
rect 22096 12480 22112 12544
rect 22176 12480 22192 12544
rect 22256 12480 22264 12544
rect 21944 11456 22264 12480
rect 21944 11392 21952 11456
rect 22016 11392 22032 11456
rect 22096 11392 22112 11456
rect 22176 11392 22192 11456
rect 22256 11392 22264 11456
rect 21944 10368 22264 11392
rect 21944 10304 21952 10368
rect 22016 10304 22032 10368
rect 22096 10304 22112 10368
rect 22176 10304 22192 10368
rect 22256 10304 22264 10368
rect 21944 9280 22264 10304
rect 21944 9216 21952 9280
rect 22016 9216 22032 9280
rect 22096 9216 22112 9280
rect 22176 9216 22192 9280
rect 22256 9216 22264 9280
rect 21944 8294 22264 9216
rect 21944 8192 21986 8294
rect 22222 8192 22264 8294
rect 21944 8128 21952 8192
rect 22256 8128 22264 8192
rect 21944 8058 21986 8128
rect 22222 8058 22264 8128
rect 21944 7104 22264 8058
rect 21944 7040 21952 7104
rect 22016 7040 22032 7104
rect 22096 7040 22112 7104
rect 22176 7040 22192 7104
rect 22256 7040 22264 7104
rect 21944 6016 22264 7040
rect 21944 5952 21952 6016
rect 22016 5952 22032 6016
rect 22096 5952 22112 6016
rect 22176 5952 22192 6016
rect 22256 5952 22264 6016
rect 21944 4928 22264 5952
rect 21944 4864 21952 4928
rect 22016 4864 22032 4928
rect 22096 4864 22112 4928
rect 22176 4864 22192 4928
rect 22256 4864 22264 4928
rect 21944 3840 22264 4864
rect 21944 3776 21952 3840
rect 22016 3776 22032 3840
rect 22096 3776 22112 3840
rect 22176 3776 22192 3840
rect 22256 3776 22264 3840
rect 21944 3294 22264 3776
rect 21944 3058 21986 3294
rect 22222 3058 22264 3294
rect 21944 2752 22264 3058
rect 21944 2688 21952 2752
rect 22016 2688 22032 2752
rect 22096 2688 22112 2752
rect 22176 2688 22192 2752
rect 22256 2688 22264 2752
rect 21944 2128 22264 2688
rect 22604 69664 22924 69680
rect 22604 69600 22612 69664
rect 22676 69600 22692 69664
rect 22756 69600 22772 69664
rect 22836 69600 22852 69664
rect 22916 69600 22924 69664
rect 22604 68954 22924 69600
rect 22604 68718 22646 68954
rect 22882 68718 22924 68954
rect 22604 68576 22924 68718
rect 22604 68512 22612 68576
rect 22676 68512 22692 68576
rect 22756 68512 22772 68576
rect 22836 68512 22852 68576
rect 22916 68512 22924 68576
rect 22604 67488 22924 68512
rect 22604 67424 22612 67488
rect 22676 67424 22692 67488
rect 22756 67424 22772 67488
rect 22836 67424 22852 67488
rect 22916 67424 22924 67488
rect 22604 66400 22924 67424
rect 22604 66336 22612 66400
rect 22676 66336 22692 66400
rect 22756 66336 22772 66400
rect 22836 66336 22852 66400
rect 22916 66336 22924 66400
rect 22604 65312 22924 66336
rect 22604 65248 22612 65312
rect 22676 65248 22692 65312
rect 22756 65248 22772 65312
rect 22836 65248 22852 65312
rect 22916 65248 22924 65312
rect 22604 64224 22924 65248
rect 22604 64160 22612 64224
rect 22676 64160 22692 64224
rect 22756 64160 22772 64224
rect 22836 64160 22852 64224
rect 22916 64160 22924 64224
rect 22604 63954 22924 64160
rect 22604 63718 22646 63954
rect 22882 63718 22924 63954
rect 22604 63136 22924 63718
rect 22604 63072 22612 63136
rect 22676 63072 22692 63136
rect 22756 63072 22772 63136
rect 22836 63072 22852 63136
rect 22916 63072 22924 63136
rect 22604 62048 22924 63072
rect 22604 61984 22612 62048
rect 22676 61984 22692 62048
rect 22756 61984 22772 62048
rect 22836 61984 22852 62048
rect 22916 61984 22924 62048
rect 22604 60960 22924 61984
rect 22604 60896 22612 60960
rect 22676 60896 22692 60960
rect 22756 60896 22772 60960
rect 22836 60896 22852 60960
rect 22916 60896 22924 60960
rect 22604 59872 22924 60896
rect 22604 59808 22612 59872
rect 22676 59808 22692 59872
rect 22756 59808 22772 59872
rect 22836 59808 22852 59872
rect 22916 59808 22924 59872
rect 22604 58954 22924 59808
rect 22604 58784 22646 58954
rect 22882 58784 22924 58954
rect 22604 58720 22612 58784
rect 22916 58720 22924 58784
rect 22604 58718 22646 58720
rect 22882 58718 22924 58720
rect 22604 57696 22924 58718
rect 22604 57632 22612 57696
rect 22676 57632 22692 57696
rect 22756 57632 22772 57696
rect 22836 57632 22852 57696
rect 22916 57632 22924 57696
rect 22604 56608 22924 57632
rect 22604 56544 22612 56608
rect 22676 56544 22692 56608
rect 22756 56544 22772 56608
rect 22836 56544 22852 56608
rect 22916 56544 22924 56608
rect 22604 55520 22924 56544
rect 22604 55456 22612 55520
rect 22676 55456 22692 55520
rect 22756 55456 22772 55520
rect 22836 55456 22852 55520
rect 22916 55456 22924 55520
rect 22604 54432 22924 55456
rect 22604 54368 22612 54432
rect 22676 54368 22692 54432
rect 22756 54368 22772 54432
rect 22836 54368 22852 54432
rect 22916 54368 22924 54432
rect 22604 53954 22924 54368
rect 22604 53718 22646 53954
rect 22882 53718 22924 53954
rect 22604 53344 22924 53718
rect 22604 53280 22612 53344
rect 22676 53280 22692 53344
rect 22756 53280 22772 53344
rect 22836 53280 22852 53344
rect 22916 53280 22924 53344
rect 22604 52256 22924 53280
rect 22604 52192 22612 52256
rect 22676 52192 22692 52256
rect 22756 52192 22772 52256
rect 22836 52192 22852 52256
rect 22916 52192 22924 52256
rect 22604 51168 22924 52192
rect 22604 51104 22612 51168
rect 22676 51104 22692 51168
rect 22756 51104 22772 51168
rect 22836 51104 22852 51168
rect 22916 51104 22924 51168
rect 22604 50080 22924 51104
rect 22604 50016 22612 50080
rect 22676 50016 22692 50080
rect 22756 50016 22772 50080
rect 22836 50016 22852 50080
rect 22916 50016 22924 50080
rect 22604 48992 22924 50016
rect 22604 48928 22612 48992
rect 22676 48954 22692 48992
rect 22756 48954 22772 48992
rect 22836 48954 22852 48992
rect 22916 48928 22924 48992
rect 22604 48718 22646 48928
rect 22882 48718 22924 48928
rect 22604 47904 22924 48718
rect 22604 47840 22612 47904
rect 22676 47840 22692 47904
rect 22756 47840 22772 47904
rect 22836 47840 22852 47904
rect 22916 47840 22924 47904
rect 22604 46816 22924 47840
rect 22604 46752 22612 46816
rect 22676 46752 22692 46816
rect 22756 46752 22772 46816
rect 22836 46752 22852 46816
rect 22916 46752 22924 46816
rect 22604 45728 22924 46752
rect 22604 45664 22612 45728
rect 22676 45664 22692 45728
rect 22756 45664 22772 45728
rect 22836 45664 22852 45728
rect 22916 45664 22924 45728
rect 22604 44640 22924 45664
rect 22604 44576 22612 44640
rect 22676 44576 22692 44640
rect 22756 44576 22772 44640
rect 22836 44576 22852 44640
rect 22916 44576 22924 44640
rect 22604 43954 22924 44576
rect 22604 43718 22646 43954
rect 22882 43718 22924 43954
rect 22604 43552 22924 43718
rect 22604 43488 22612 43552
rect 22676 43488 22692 43552
rect 22756 43488 22772 43552
rect 22836 43488 22852 43552
rect 22916 43488 22924 43552
rect 22604 42464 22924 43488
rect 22604 42400 22612 42464
rect 22676 42400 22692 42464
rect 22756 42400 22772 42464
rect 22836 42400 22852 42464
rect 22916 42400 22924 42464
rect 22604 41376 22924 42400
rect 22604 41312 22612 41376
rect 22676 41312 22692 41376
rect 22756 41312 22772 41376
rect 22836 41312 22852 41376
rect 22916 41312 22924 41376
rect 22604 40288 22924 41312
rect 22604 40224 22612 40288
rect 22676 40224 22692 40288
rect 22756 40224 22772 40288
rect 22836 40224 22852 40288
rect 22916 40224 22924 40288
rect 22604 39200 22924 40224
rect 22604 39136 22612 39200
rect 22676 39136 22692 39200
rect 22756 39136 22772 39200
rect 22836 39136 22852 39200
rect 22916 39136 22924 39200
rect 22604 38954 22924 39136
rect 22604 38718 22646 38954
rect 22882 38718 22924 38954
rect 22604 38112 22924 38718
rect 22604 38048 22612 38112
rect 22676 38048 22692 38112
rect 22756 38048 22772 38112
rect 22836 38048 22852 38112
rect 22916 38048 22924 38112
rect 22604 37024 22924 38048
rect 22604 36960 22612 37024
rect 22676 36960 22692 37024
rect 22756 36960 22772 37024
rect 22836 36960 22852 37024
rect 22916 36960 22924 37024
rect 22604 35936 22924 36960
rect 22604 35872 22612 35936
rect 22676 35872 22692 35936
rect 22756 35872 22772 35936
rect 22836 35872 22852 35936
rect 22916 35872 22924 35936
rect 22604 34848 22924 35872
rect 22604 34784 22612 34848
rect 22676 34784 22692 34848
rect 22756 34784 22772 34848
rect 22836 34784 22852 34848
rect 22916 34784 22924 34848
rect 22604 33954 22924 34784
rect 22604 33760 22646 33954
rect 22882 33760 22924 33954
rect 22604 33696 22612 33760
rect 22676 33696 22692 33718
rect 22756 33696 22772 33718
rect 22836 33696 22852 33718
rect 22916 33696 22924 33760
rect 22604 32672 22924 33696
rect 22604 32608 22612 32672
rect 22676 32608 22692 32672
rect 22756 32608 22772 32672
rect 22836 32608 22852 32672
rect 22916 32608 22924 32672
rect 22604 31584 22924 32608
rect 22604 31520 22612 31584
rect 22676 31520 22692 31584
rect 22756 31520 22772 31584
rect 22836 31520 22852 31584
rect 22916 31520 22924 31584
rect 22604 30496 22924 31520
rect 22604 30432 22612 30496
rect 22676 30432 22692 30496
rect 22756 30432 22772 30496
rect 22836 30432 22852 30496
rect 22916 30432 22924 30496
rect 22604 29408 22924 30432
rect 22604 29344 22612 29408
rect 22676 29344 22692 29408
rect 22756 29344 22772 29408
rect 22836 29344 22852 29408
rect 22916 29344 22924 29408
rect 22604 28954 22924 29344
rect 22604 28718 22646 28954
rect 22882 28718 22924 28954
rect 22604 28320 22924 28718
rect 22604 28256 22612 28320
rect 22676 28256 22692 28320
rect 22756 28256 22772 28320
rect 22836 28256 22852 28320
rect 22916 28256 22924 28320
rect 22604 27232 22924 28256
rect 22604 27168 22612 27232
rect 22676 27168 22692 27232
rect 22756 27168 22772 27232
rect 22836 27168 22852 27232
rect 22916 27168 22924 27232
rect 22604 26144 22924 27168
rect 22604 26080 22612 26144
rect 22676 26080 22692 26144
rect 22756 26080 22772 26144
rect 22836 26080 22852 26144
rect 22916 26080 22924 26144
rect 22604 25056 22924 26080
rect 22604 24992 22612 25056
rect 22676 24992 22692 25056
rect 22756 24992 22772 25056
rect 22836 24992 22852 25056
rect 22916 24992 22924 25056
rect 22604 23968 22924 24992
rect 22604 23904 22612 23968
rect 22676 23954 22692 23968
rect 22756 23954 22772 23968
rect 22836 23954 22852 23968
rect 22916 23904 22924 23968
rect 22604 23718 22646 23904
rect 22882 23718 22924 23904
rect 22604 22880 22924 23718
rect 22604 22816 22612 22880
rect 22676 22816 22692 22880
rect 22756 22816 22772 22880
rect 22836 22816 22852 22880
rect 22916 22816 22924 22880
rect 22604 21792 22924 22816
rect 22604 21728 22612 21792
rect 22676 21728 22692 21792
rect 22756 21728 22772 21792
rect 22836 21728 22852 21792
rect 22916 21728 22924 21792
rect 22604 20704 22924 21728
rect 22604 20640 22612 20704
rect 22676 20640 22692 20704
rect 22756 20640 22772 20704
rect 22836 20640 22852 20704
rect 22916 20640 22924 20704
rect 22604 19616 22924 20640
rect 22604 19552 22612 19616
rect 22676 19552 22692 19616
rect 22756 19552 22772 19616
rect 22836 19552 22852 19616
rect 22916 19552 22924 19616
rect 22604 18954 22924 19552
rect 22604 18718 22646 18954
rect 22882 18718 22924 18954
rect 22604 18528 22924 18718
rect 22604 18464 22612 18528
rect 22676 18464 22692 18528
rect 22756 18464 22772 18528
rect 22836 18464 22852 18528
rect 22916 18464 22924 18528
rect 22604 17440 22924 18464
rect 22604 17376 22612 17440
rect 22676 17376 22692 17440
rect 22756 17376 22772 17440
rect 22836 17376 22852 17440
rect 22916 17376 22924 17440
rect 22604 16352 22924 17376
rect 22604 16288 22612 16352
rect 22676 16288 22692 16352
rect 22756 16288 22772 16352
rect 22836 16288 22852 16352
rect 22916 16288 22924 16352
rect 22604 15264 22924 16288
rect 22604 15200 22612 15264
rect 22676 15200 22692 15264
rect 22756 15200 22772 15264
rect 22836 15200 22852 15264
rect 22916 15200 22924 15264
rect 22604 14176 22924 15200
rect 22604 14112 22612 14176
rect 22676 14112 22692 14176
rect 22756 14112 22772 14176
rect 22836 14112 22852 14176
rect 22916 14112 22924 14176
rect 22604 13954 22924 14112
rect 22604 13718 22646 13954
rect 22882 13718 22924 13954
rect 22604 13088 22924 13718
rect 22604 13024 22612 13088
rect 22676 13024 22692 13088
rect 22756 13024 22772 13088
rect 22836 13024 22852 13088
rect 22916 13024 22924 13088
rect 22604 12000 22924 13024
rect 22604 11936 22612 12000
rect 22676 11936 22692 12000
rect 22756 11936 22772 12000
rect 22836 11936 22852 12000
rect 22916 11936 22924 12000
rect 22604 10912 22924 11936
rect 22604 10848 22612 10912
rect 22676 10848 22692 10912
rect 22756 10848 22772 10912
rect 22836 10848 22852 10912
rect 22916 10848 22924 10912
rect 22604 9824 22924 10848
rect 22604 9760 22612 9824
rect 22676 9760 22692 9824
rect 22756 9760 22772 9824
rect 22836 9760 22852 9824
rect 22916 9760 22924 9824
rect 22604 8954 22924 9760
rect 22604 8736 22646 8954
rect 22882 8736 22924 8954
rect 22604 8672 22612 8736
rect 22676 8672 22692 8718
rect 22756 8672 22772 8718
rect 22836 8672 22852 8718
rect 22916 8672 22924 8736
rect 22604 7648 22924 8672
rect 22604 7584 22612 7648
rect 22676 7584 22692 7648
rect 22756 7584 22772 7648
rect 22836 7584 22852 7648
rect 22916 7584 22924 7648
rect 22604 6560 22924 7584
rect 22604 6496 22612 6560
rect 22676 6496 22692 6560
rect 22756 6496 22772 6560
rect 22836 6496 22852 6560
rect 22916 6496 22924 6560
rect 22604 5472 22924 6496
rect 22604 5408 22612 5472
rect 22676 5408 22692 5472
rect 22756 5408 22772 5472
rect 22836 5408 22852 5472
rect 22916 5408 22924 5472
rect 22604 4384 22924 5408
rect 22604 4320 22612 4384
rect 22676 4320 22692 4384
rect 22756 4320 22772 4384
rect 22836 4320 22852 4384
rect 22916 4320 22924 4384
rect 22604 3954 22924 4320
rect 22604 3718 22646 3954
rect 22882 3718 22924 3954
rect 22604 3296 22924 3718
rect 22604 3232 22612 3296
rect 22676 3232 22692 3296
rect 22756 3232 22772 3296
rect 22836 3232 22852 3296
rect 22916 3232 22924 3296
rect 22604 2208 22924 3232
rect 22604 2144 22612 2208
rect 22676 2144 22692 2208
rect 22756 2144 22772 2208
rect 22836 2144 22852 2208
rect 22916 2144 22924 2208
rect 22604 2128 22924 2144
rect 26944 69120 27264 69680
rect 26944 69056 26952 69120
rect 27016 69056 27032 69120
rect 27096 69056 27112 69120
rect 27176 69056 27192 69120
rect 27256 69056 27264 69120
rect 26944 68294 27264 69056
rect 26944 68058 26986 68294
rect 27222 68058 27264 68294
rect 26944 68032 27264 68058
rect 26944 67968 26952 68032
rect 27016 67968 27032 68032
rect 27096 67968 27112 68032
rect 27176 67968 27192 68032
rect 27256 67968 27264 68032
rect 26944 66944 27264 67968
rect 26944 66880 26952 66944
rect 27016 66880 27032 66944
rect 27096 66880 27112 66944
rect 27176 66880 27192 66944
rect 27256 66880 27264 66944
rect 26944 65856 27264 66880
rect 26944 65792 26952 65856
rect 27016 65792 27032 65856
rect 27096 65792 27112 65856
rect 27176 65792 27192 65856
rect 27256 65792 27264 65856
rect 26944 64768 27264 65792
rect 26944 64704 26952 64768
rect 27016 64704 27032 64768
rect 27096 64704 27112 64768
rect 27176 64704 27192 64768
rect 27256 64704 27264 64768
rect 26944 63680 27264 64704
rect 26944 63616 26952 63680
rect 27016 63616 27032 63680
rect 27096 63616 27112 63680
rect 27176 63616 27192 63680
rect 27256 63616 27264 63680
rect 26944 63294 27264 63616
rect 26944 63058 26986 63294
rect 27222 63058 27264 63294
rect 26944 62592 27264 63058
rect 26944 62528 26952 62592
rect 27016 62528 27032 62592
rect 27096 62528 27112 62592
rect 27176 62528 27192 62592
rect 27256 62528 27264 62592
rect 26944 61504 27264 62528
rect 26944 61440 26952 61504
rect 27016 61440 27032 61504
rect 27096 61440 27112 61504
rect 27176 61440 27192 61504
rect 27256 61440 27264 61504
rect 26944 60416 27264 61440
rect 26944 60352 26952 60416
rect 27016 60352 27032 60416
rect 27096 60352 27112 60416
rect 27176 60352 27192 60416
rect 27256 60352 27264 60416
rect 26944 59328 27264 60352
rect 26944 59264 26952 59328
rect 27016 59264 27032 59328
rect 27096 59264 27112 59328
rect 27176 59264 27192 59328
rect 27256 59264 27264 59328
rect 26944 58294 27264 59264
rect 26944 58240 26986 58294
rect 27222 58240 27264 58294
rect 26944 58176 26952 58240
rect 27256 58176 27264 58240
rect 26944 58058 26986 58176
rect 27222 58058 27264 58176
rect 26944 57152 27264 58058
rect 26944 57088 26952 57152
rect 27016 57088 27032 57152
rect 27096 57088 27112 57152
rect 27176 57088 27192 57152
rect 27256 57088 27264 57152
rect 26944 56064 27264 57088
rect 26944 56000 26952 56064
rect 27016 56000 27032 56064
rect 27096 56000 27112 56064
rect 27176 56000 27192 56064
rect 27256 56000 27264 56064
rect 26944 54976 27264 56000
rect 26944 54912 26952 54976
rect 27016 54912 27032 54976
rect 27096 54912 27112 54976
rect 27176 54912 27192 54976
rect 27256 54912 27264 54976
rect 26944 53888 27264 54912
rect 26944 53824 26952 53888
rect 27016 53824 27032 53888
rect 27096 53824 27112 53888
rect 27176 53824 27192 53888
rect 27256 53824 27264 53888
rect 26944 53294 27264 53824
rect 26944 53058 26986 53294
rect 27222 53058 27264 53294
rect 26944 52800 27264 53058
rect 26944 52736 26952 52800
rect 27016 52736 27032 52800
rect 27096 52736 27112 52800
rect 27176 52736 27192 52800
rect 27256 52736 27264 52800
rect 26944 51712 27264 52736
rect 26944 51648 26952 51712
rect 27016 51648 27032 51712
rect 27096 51648 27112 51712
rect 27176 51648 27192 51712
rect 27256 51648 27264 51712
rect 26944 50624 27264 51648
rect 26944 50560 26952 50624
rect 27016 50560 27032 50624
rect 27096 50560 27112 50624
rect 27176 50560 27192 50624
rect 27256 50560 27264 50624
rect 26944 49536 27264 50560
rect 26944 49472 26952 49536
rect 27016 49472 27032 49536
rect 27096 49472 27112 49536
rect 27176 49472 27192 49536
rect 27256 49472 27264 49536
rect 26944 48448 27264 49472
rect 26944 48384 26952 48448
rect 27016 48384 27032 48448
rect 27096 48384 27112 48448
rect 27176 48384 27192 48448
rect 27256 48384 27264 48448
rect 26944 48294 27264 48384
rect 26944 48058 26986 48294
rect 27222 48058 27264 48294
rect 26944 47360 27264 48058
rect 26944 47296 26952 47360
rect 27016 47296 27032 47360
rect 27096 47296 27112 47360
rect 27176 47296 27192 47360
rect 27256 47296 27264 47360
rect 26944 46272 27264 47296
rect 26944 46208 26952 46272
rect 27016 46208 27032 46272
rect 27096 46208 27112 46272
rect 27176 46208 27192 46272
rect 27256 46208 27264 46272
rect 26944 45184 27264 46208
rect 26944 45120 26952 45184
rect 27016 45120 27032 45184
rect 27096 45120 27112 45184
rect 27176 45120 27192 45184
rect 27256 45120 27264 45184
rect 26944 44096 27264 45120
rect 26944 44032 26952 44096
rect 27016 44032 27032 44096
rect 27096 44032 27112 44096
rect 27176 44032 27192 44096
rect 27256 44032 27264 44096
rect 26944 43294 27264 44032
rect 26944 43058 26986 43294
rect 27222 43058 27264 43294
rect 26944 43008 27264 43058
rect 26944 42944 26952 43008
rect 27016 42944 27032 43008
rect 27096 42944 27112 43008
rect 27176 42944 27192 43008
rect 27256 42944 27264 43008
rect 26944 41920 27264 42944
rect 26944 41856 26952 41920
rect 27016 41856 27032 41920
rect 27096 41856 27112 41920
rect 27176 41856 27192 41920
rect 27256 41856 27264 41920
rect 26944 40832 27264 41856
rect 26944 40768 26952 40832
rect 27016 40768 27032 40832
rect 27096 40768 27112 40832
rect 27176 40768 27192 40832
rect 27256 40768 27264 40832
rect 26944 39744 27264 40768
rect 26944 39680 26952 39744
rect 27016 39680 27032 39744
rect 27096 39680 27112 39744
rect 27176 39680 27192 39744
rect 27256 39680 27264 39744
rect 26944 38656 27264 39680
rect 26944 38592 26952 38656
rect 27016 38592 27032 38656
rect 27096 38592 27112 38656
rect 27176 38592 27192 38656
rect 27256 38592 27264 38656
rect 26944 38294 27264 38592
rect 26944 38058 26986 38294
rect 27222 38058 27264 38294
rect 26944 37568 27264 38058
rect 26944 37504 26952 37568
rect 27016 37504 27032 37568
rect 27096 37504 27112 37568
rect 27176 37504 27192 37568
rect 27256 37504 27264 37568
rect 26944 36480 27264 37504
rect 26944 36416 26952 36480
rect 27016 36416 27032 36480
rect 27096 36416 27112 36480
rect 27176 36416 27192 36480
rect 27256 36416 27264 36480
rect 26944 35392 27264 36416
rect 26944 35328 26952 35392
rect 27016 35328 27032 35392
rect 27096 35328 27112 35392
rect 27176 35328 27192 35392
rect 27256 35328 27264 35392
rect 26944 34304 27264 35328
rect 26944 34240 26952 34304
rect 27016 34240 27032 34304
rect 27096 34240 27112 34304
rect 27176 34240 27192 34304
rect 27256 34240 27264 34304
rect 26944 33294 27264 34240
rect 26944 33216 26986 33294
rect 27222 33216 27264 33294
rect 26944 33152 26952 33216
rect 27256 33152 27264 33216
rect 26944 33058 26986 33152
rect 27222 33058 27264 33152
rect 26944 32128 27264 33058
rect 26944 32064 26952 32128
rect 27016 32064 27032 32128
rect 27096 32064 27112 32128
rect 27176 32064 27192 32128
rect 27256 32064 27264 32128
rect 26944 31040 27264 32064
rect 26944 30976 26952 31040
rect 27016 30976 27032 31040
rect 27096 30976 27112 31040
rect 27176 30976 27192 31040
rect 27256 30976 27264 31040
rect 26944 29952 27264 30976
rect 26944 29888 26952 29952
rect 27016 29888 27032 29952
rect 27096 29888 27112 29952
rect 27176 29888 27192 29952
rect 27256 29888 27264 29952
rect 26944 28864 27264 29888
rect 26944 28800 26952 28864
rect 27016 28800 27032 28864
rect 27096 28800 27112 28864
rect 27176 28800 27192 28864
rect 27256 28800 27264 28864
rect 26944 28294 27264 28800
rect 26944 28058 26986 28294
rect 27222 28058 27264 28294
rect 26944 27776 27264 28058
rect 26944 27712 26952 27776
rect 27016 27712 27032 27776
rect 27096 27712 27112 27776
rect 27176 27712 27192 27776
rect 27256 27712 27264 27776
rect 26944 26688 27264 27712
rect 26944 26624 26952 26688
rect 27016 26624 27032 26688
rect 27096 26624 27112 26688
rect 27176 26624 27192 26688
rect 27256 26624 27264 26688
rect 26944 25600 27264 26624
rect 26944 25536 26952 25600
rect 27016 25536 27032 25600
rect 27096 25536 27112 25600
rect 27176 25536 27192 25600
rect 27256 25536 27264 25600
rect 26944 24512 27264 25536
rect 26944 24448 26952 24512
rect 27016 24448 27032 24512
rect 27096 24448 27112 24512
rect 27176 24448 27192 24512
rect 27256 24448 27264 24512
rect 26944 23424 27264 24448
rect 26944 23360 26952 23424
rect 27016 23360 27032 23424
rect 27096 23360 27112 23424
rect 27176 23360 27192 23424
rect 27256 23360 27264 23424
rect 26944 23294 27264 23360
rect 26944 23058 26986 23294
rect 27222 23058 27264 23294
rect 26944 22336 27264 23058
rect 26944 22272 26952 22336
rect 27016 22272 27032 22336
rect 27096 22272 27112 22336
rect 27176 22272 27192 22336
rect 27256 22272 27264 22336
rect 26944 21248 27264 22272
rect 26944 21184 26952 21248
rect 27016 21184 27032 21248
rect 27096 21184 27112 21248
rect 27176 21184 27192 21248
rect 27256 21184 27264 21248
rect 26944 20160 27264 21184
rect 26944 20096 26952 20160
rect 27016 20096 27032 20160
rect 27096 20096 27112 20160
rect 27176 20096 27192 20160
rect 27256 20096 27264 20160
rect 26944 19072 27264 20096
rect 26944 19008 26952 19072
rect 27016 19008 27032 19072
rect 27096 19008 27112 19072
rect 27176 19008 27192 19072
rect 27256 19008 27264 19072
rect 26944 18294 27264 19008
rect 26944 18058 26986 18294
rect 27222 18058 27264 18294
rect 26944 17984 27264 18058
rect 26944 17920 26952 17984
rect 27016 17920 27032 17984
rect 27096 17920 27112 17984
rect 27176 17920 27192 17984
rect 27256 17920 27264 17984
rect 26944 16896 27264 17920
rect 26944 16832 26952 16896
rect 27016 16832 27032 16896
rect 27096 16832 27112 16896
rect 27176 16832 27192 16896
rect 27256 16832 27264 16896
rect 26944 15808 27264 16832
rect 26944 15744 26952 15808
rect 27016 15744 27032 15808
rect 27096 15744 27112 15808
rect 27176 15744 27192 15808
rect 27256 15744 27264 15808
rect 26944 14720 27264 15744
rect 26944 14656 26952 14720
rect 27016 14656 27032 14720
rect 27096 14656 27112 14720
rect 27176 14656 27192 14720
rect 27256 14656 27264 14720
rect 26944 13632 27264 14656
rect 26944 13568 26952 13632
rect 27016 13568 27032 13632
rect 27096 13568 27112 13632
rect 27176 13568 27192 13632
rect 27256 13568 27264 13632
rect 26944 13294 27264 13568
rect 26944 13058 26986 13294
rect 27222 13058 27264 13294
rect 26944 12544 27264 13058
rect 26944 12480 26952 12544
rect 27016 12480 27032 12544
rect 27096 12480 27112 12544
rect 27176 12480 27192 12544
rect 27256 12480 27264 12544
rect 26944 11456 27264 12480
rect 26944 11392 26952 11456
rect 27016 11392 27032 11456
rect 27096 11392 27112 11456
rect 27176 11392 27192 11456
rect 27256 11392 27264 11456
rect 26944 10368 27264 11392
rect 26944 10304 26952 10368
rect 27016 10304 27032 10368
rect 27096 10304 27112 10368
rect 27176 10304 27192 10368
rect 27256 10304 27264 10368
rect 26944 9280 27264 10304
rect 26944 9216 26952 9280
rect 27016 9216 27032 9280
rect 27096 9216 27112 9280
rect 27176 9216 27192 9280
rect 27256 9216 27264 9280
rect 26944 8294 27264 9216
rect 26944 8192 26986 8294
rect 27222 8192 27264 8294
rect 26944 8128 26952 8192
rect 27256 8128 27264 8192
rect 26944 8058 26986 8128
rect 27222 8058 27264 8128
rect 26944 7104 27264 8058
rect 26944 7040 26952 7104
rect 27016 7040 27032 7104
rect 27096 7040 27112 7104
rect 27176 7040 27192 7104
rect 27256 7040 27264 7104
rect 26944 6016 27264 7040
rect 26944 5952 26952 6016
rect 27016 5952 27032 6016
rect 27096 5952 27112 6016
rect 27176 5952 27192 6016
rect 27256 5952 27264 6016
rect 26944 4928 27264 5952
rect 26944 4864 26952 4928
rect 27016 4864 27032 4928
rect 27096 4864 27112 4928
rect 27176 4864 27192 4928
rect 27256 4864 27264 4928
rect 26944 3840 27264 4864
rect 26944 3776 26952 3840
rect 27016 3776 27032 3840
rect 27096 3776 27112 3840
rect 27176 3776 27192 3840
rect 27256 3776 27264 3840
rect 26944 3294 27264 3776
rect 26944 3058 26986 3294
rect 27222 3058 27264 3294
rect 26944 2752 27264 3058
rect 26944 2688 26952 2752
rect 27016 2688 27032 2752
rect 27096 2688 27112 2752
rect 27176 2688 27192 2752
rect 27256 2688 27264 2752
rect 26944 2128 27264 2688
rect 27604 69664 27924 69680
rect 27604 69600 27612 69664
rect 27676 69600 27692 69664
rect 27756 69600 27772 69664
rect 27836 69600 27852 69664
rect 27916 69600 27924 69664
rect 27604 68954 27924 69600
rect 27604 68718 27646 68954
rect 27882 68718 27924 68954
rect 27604 68576 27924 68718
rect 27604 68512 27612 68576
rect 27676 68512 27692 68576
rect 27756 68512 27772 68576
rect 27836 68512 27852 68576
rect 27916 68512 27924 68576
rect 27604 67488 27924 68512
rect 31944 69120 32264 69680
rect 31944 69056 31952 69120
rect 32016 69056 32032 69120
rect 32096 69056 32112 69120
rect 32176 69056 32192 69120
rect 32256 69056 32264 69120
rect 31944 68294 32264 69056
rect 31944 68058 31986 68294
rect 32222 68058 32264 68294
rect 31944 68032 32264 68058
rect 31944 67968 31952 68032
rect 32016 67968 32032 68032
rect 32096 67968 32112 68032
rect 32176 67968 32192 68032
rect 32256 67968 32264 68032
rect 31707 67692 31773 67693
rect 31707 67628 31708 67692
rect 31772 67628 31773 67692
rect 31707 67627 31773 67628
rect 27604 67424 27612 67488
rect 27676 67424 27692 67488
rect 27756 67424 27772 67488
rect 27836 67424 27852 67488
rect 27916 67424 27924 67488
rect 27604 66400 27924 67424
rect 27604 66336 27612 66400
rect 27676 66336 27692 66400
rect 27756 66336 27772 66400
rect 27836 66336 27852 66400
rect 27916 66336 27924 66400
rect 27604 65312 27924 66336
rect 27604 65248 27612 65312
rect 27676 65248 27692 65312
rect 27756 65248 27772 65312
rect 27836 65248 27852 65312
rect 27916 65248 27924 65312
rect 27604 64224 27924 65248
rect 27604 64160 27612 64224
rect 27676 64160 27692 64224
rect 27756 64160 27772 64224
rect 27836 64160 27852 64224
rect 27916 64160 27924 64224
rect 27604 63954 27924 64160
rect 27604 63718 27646 63954
rect 27882 63718 27924 63954
rect 27604 63136 27924 63718
rect 27604 63072 27612 63136
rect 27676 63072 27692 63136
rect 27756 63072 27772 63136
rect 27836 63072 27852 63136
rect 27916 63072 27924 63136
rect 27604 62048 27924 63072
rect 27604 61984 27612 62048
rect 27676 61984 27692 62048
rect 27756 61984 27772 62048
rect 27836 61984 27852 62048
rect 27916 61984 27924 62048
rect 27604 60960 27924 61984
rect 27604 60896 27612 60960
rect 27676 60896 27692 60960
rect 27756 60896 27772 60960
rect 27836 60896 27852 60960
rect 27916 60896 27924 60960
rect 27604 59872 27924 60896
rect 27604 59808 27612 59872
rect 27676 59808 27692 59872
rect 27756 59808 27772 59872
rect 27836 59808 27852 59872
rect 27916 59808 27924 59872
rect 27604 58954 27924 59808
rect 27604 58784 27646 58954
rect 27882 58784 27924 58954
rect 27604 58720 27612 58784
rect 27916 58720 27924 58784
rect 27604 58718 27646 58720
rect 27882 58718 27924 58720
rect 27604 57696 27924 58718
rect 27604 57632 27612 57696
rect 27676 57632 27692 57696
rect 27756 57632 27772 57696
rect 27836 57632 27852 57696
rect 27916 57632 27924 57696
rect 27604 56608 27924 57632
rect 27604 56544 27612 56608
rect 27676 56544 27692 56608
rect 27756 56544 27772 56608
rect 27836 56544 27852 56608
rect 27916 56544 27924 56608
rect 27604 55520 27924 56544
rect 27604 55456 27612 55520
rect 27676 55456 27692 55520
rect 27756 55456 27772 55520
rect 27836 55456 27852 55520
rect 27916 55456 27924 55520
rect 27604 54432 27924 55456
rect 27604 54368 27612 54432
rect 27676 54368 27692 54432
rect 27756 54368 27772 54432
rect 27836 54368 27852 54432
rect 27916 54368 27924 54432
rect 27604 53954 27924 54368
rect 27604 53718 27646 53954
rect 27882 53718 27924 53954
rect 27604 53344 27924 53718
rect 27604 53280 27612 53344
rect 27676 53280 27692 53344
rect 27756 53280 27772 53344
rect 27836 53280 27852 53344
rect 27916 53280 27924 53344
rect 27604 52256 27924 53280
rect 27604 52192 27612 52256
rect 27676 52192 27692 52256
rect 27756 52192 27772 52256
rect 27836 52192 27852 52256
rect 27916 52192 27924 52256
rect 27604 51168 27924 52192
rect 27604 51104 27612 51168
rect 27676 51104 27692 51168
rect 27756 51104 27772 51168
rect 27836 51104 27852 51168
rect 27916 51104 27924 51168
rect 27604 50080 27924 51104
rect 31710 50965 31770 67627
rect 31944 66944 32264 67968
rect 31944 66880 31952 66944
rect 32016 66880 32032 66944
rect 32096 66880 32112 66944
rect 32176 66880 32192 66944
rect 32256 66880 32264 66944
rect 31944 65856 32264 66880
rect 31944 65792 31952 65856
rect 32016 65792 32032 65856
rect 32096 65792 32112 65856
rect 32176 65792 32192 65856
rect 32256 65792 32264 65856
rect 31944 64768 32264 65792
rect 31944 64704 31952 64768
rect 32016 64704 32032 64768
rect 32096 64704 32112 64768
rect 32176 64704 32192 64768
rect 32256 64704 32264 64768
rect 31944 63680 32264 64704
rect 31944 63616 31952 63680
rect 32016 63616 32032 63680
rect 32096 63616 32112 63680
rect 32176 63616 32192 63680
rect 32256 63616 32264 63680
rect 31944 63294 32264 63616
rect 31944 63058 31986 63294
rect 32222 63058 32264 63294
rect 31944 62592 32264 63058
rect 31944 62528 31952 62592
rect 32016 62528 32032 62592
rect 32096 62528 32112 62592
rect 32176 62528 32192 62592
rect 32256 62528 32264 62592
rect 31944 61504 32264 62528
rect 31944 61440 31952 61504
rect 32016 61440 32032 61504
rect 32096 61440 32112 61504
rect 32176 61440 32192 61504
rect 32256 61440 32264 61504
rect 31944 60416 32264 61440
rect 31944 60352 31952 60416
rect 32016 60352 32032 60416
rect 32096 60352 32112 60416
rect 32176 60352 32192 60416
rect 32256 60352 32264 60416
rect 31944 59328 32264 60352
rect 31944 59264 31952 59328
rect 32016 59264 32032 59328
rect 32096 59264 32112 59328
rect 32176 59264 32192 59328
rect 32256 59264 32264 59328
rect 31944 58294 32264 59264
rect 31944 58240 31986 58294
rect 32222 58240 32264 58294
rect 31944 58176 31952 58240
rect 32256 58176 32264 58240
rect 31944 58058 31986 58176
rect 32222 58058 32264 58176
rect 31944 57152 32264 58058
rect 31944 57088 31952 57152
rect 32016 57088 32032 57152
rect 32096 57088 32112 57152
rect 32176 57088 32192 57152
rect 32256 57088 32264 57152
rect 31944 56064 32264 57088
rect 31944 56000 31952 56064
rect 32016 56000 32032 56064
rect 32096 56000 32112 56064
rect 32176 56000 32192 56064
rect 32256 56000 32264 56064
rect 31944 54976 32264 56000
rect 31944 54912 31952 54976
rect 32016 54912 32032 54976
rect 32096 54912 32112 54976
rect 32176 54912 32192 54976
rect 32256 54912 32264 54976
rect 31944 53888 32264 54912
rect 31944 53824 31952 53888
rect 32016 53824 32032 53888
rect 32096 53824 32112 53888
rect 32176 53824 32192 53888
rect 32256 53824 32264 53888
rect 31944 53294 32264 53824
rect 31944 53058 31986 53294
rect 32222 53058 32264 53294
rect 31944 52800 32264 53058
rect 31944 52736 31952 52800
rect 32016 52736 32032 52800
rect 32096 52736 32112 52800
rect 32176 52736 32192 52800
rect 32256 52736 32264 52800
rect 31944 51712 32264 52736
rect 31944 51648 31952 51712
rect 32016 51648 32032 51712
rect 32096 51648 32112 51712
rect 32176 51648 32192 51712
rect 32256 51648 32264 51712
rect 31707 50964 31773 50965
rect 31707 50900 31708 50964
rect 31772 50900 31773 50964
rect 31707 50899 31773 50900
rect 27604 50016 27612 50080
rect 27676 50016 27692 50080
rect 27756 50016 27772 50080
rect 27836 50016 27852 50080
rect 27916 50016 27924 50080
rect 27604 48992 27924 50016
rect 27604 48928 27612 48992
rect 27676 48954 27692 48992
rect 27756 48954 27772 48992
rect 27836 48954 27852 48992
rect 27916 48928 27924 48992
rect 27604 48718 27646 48928
rect 27882 48718 27924 48928
rect 27604 47904 27924 48718
rect 27604 47840 27612 47904
rect 27676 47840 27692 47904
rect 27756 47840 27772 47904
rect 27836 47840 27852 47904
rect 27916 47840 27924 47904
rect 27604 46816 27924 47840
rect 27604 46752 27612 46816
rect 27676 46752 27692 46816
rect 27756 46752 27772 46816
rect 27836 46752 27852 46816
rect 27916 46752 27924 46816
rect 27604 45728 27924 46752
rect 27604 45664 27612 45728
rect 27676 45664 27692 45728
rect 27756 45664 27772 45728
rect 27836 45664 27852 45728
rect 27916 45664 27924 45728
rect 27604 44640 27924 45664
rect 27604 44576 27612 44640
rect 27676 44576 27692 44640
rect 27756 44576 27772 44640
rect 27836 44576 27852 44640
rect 27916 44576 27924 44640
rect 27604 43954 27924 44576
rect 27604 43718 27646 43954
rect 27882 43718 27924 43954
rect 27604 43552 27924 43718
rect 27604 43488 27612 43552
rect 27676 43488 27692 43552
rect 27756 43488 27772 43552
rect 27836 43488 27852 43552
rect 27916 43488 27924 43552
rect 27604 42464 27924 43488
rect 27604 42400 27612 42464
rect 27676 42400 27692 42464
rect 27756 42400 27772 42464
rect 27836 42400 27852 42464
rect 27916 42400 27924 42464
rect 27604 41376 27924 42400
rect 31944 50624 32264 51648
rect 32604 69664 32924 69680
rect 32604 69600 32612 69664
rect 32676 69600 32692 69664
rect 32756 69600 32772 69664
rect 32836 69600 32852 69664
rect 32916 69600 32924 69664
rect 32604 68954 32924 69600
rect 32604 68718 32646 68954
rect 32882 68718 32924 68954
rect 32604 68576 32924 68718
rect 32604 68512 32612 68576
rect 32676 68512 32692 68576
rect 32756 68512 32772 68576
rect 32836 68512 32852 68576
rect 32916 68512 32924 68576
rect 32604 67488 32924 68512
rect 32604 67424 32612 67488
rect 32676 67424 32692 67488
rect 32756 67424 32772 67488
rect 32836 67424 32852 67488
rect 32916 67424 32924 67488
rect 32604 66400 32924 67424
rect 32604 66336 32612 66400
rect 32676 66336 32692 66400
rect 32756 66336 32772 66400
rect 32836 66336 32852 66400
rect 32916 66336 32924 66400
rect 32604 65312 32924 66336
rect 32604 65248 32612 65312
rect 32676 65248 32692 65312
rect 32756 65248 32772 65312
rect 32836 65248 32852 65312
rect 32916 65248 32924 65312
rect 32604 64224 32924 65248
rect 32604 64160 32612 64224
rect 32676 64160 32692 64224
rect 32756 64160 32772 64224
rect 32836 64160 32852 64224
rect 32916 64160 32924 64224
rect 32604 63954 32924 64160
rect 32604 63718 32646 63954
rect 32882 63718 32924 63954
rect 32604 63136 32924 63718
rect 32604 63072 32612 63136
rect 32676 63072 32692 63136
rect 32756 63072 32772 63136
rect 32836 63072 32852 63136
rect 32916 63072 32924 63136
rect 32604 62048 32924 63072
rect 32604 61984 32612 62048
rect 32676 61984 32692 62048
rect 32756 61984 32772 62048
rect 32836 61984 32852 62048
rect 32916 61984 32924 62048
rect 32604 60960 32924 61984
rect 32604 60896 32612 60960
rect 32676 60896 32692 60960
rect 32756 60896 32772 60960
rect 32836 60896 32852 60960
rect 32916 60896 32924 60960
rect 32604 59872 32924 60896
rect 32604 59808 32612 59872
rect 32676 59808 32692 59872
rect 32756 59808 32772 59872
rect 32836 59808 32852 59872
rect 32916 59808 32924 59872
rect 32604 58954 32924 59808
rect 32604 58784 32646 58954
rect 32882 58784 32924 58954
rect 32604 58720 32612 58784
rect 32916 58720 32924 58784
rect 32604 58718 32646 58720
rect 32882 58718 32924 58720
rect 32604 57696 32924 58718
rect 36944 69120 37264 69680
rect 36944 69056 36952 69120
rect 37016 69056 37032 69120
rect 37096 69056 37112 69120
rect 37176 69056 37192 69120
rect 37256 69056 37264 69120
rect 36944 68294 37264 69056
rect 36944 68058 36986 68294
rect 37222 68058 37264 68294
rect 36944 68032 37264 68058
rect 36944 67968 36952 68032
rect 37016 67968 37032 68032
rect 37096 67968 37112 68032
rect 37176 67968 37192 68032
rect 37256 67968 37264 68032
rect 36944 66944 37264 67968
rect 36944 66880 36952 66944
rect 37016 66880 37032 66944
rect 37096 66880 37112 66944
rect 37176 66880 37192 66944
rect 37256 66880 37264 66944
rect 36944 65856 37264 66880
rect 36944 65792 36952 65856
rect 37016 65792 37032 65856
rect 37096 65792 37112 65856
rect 37176 65792 37192 65856
rect 37256 65792 37264 65856
rect 36944 64768 37264 65792
rect 36944 64704 36952 64768
rect 37016 64704 37032 64768
rect 37096 64704 37112 64768
rect 37176 64704 37192 64768
rect 37256 64704 37264 64768
rect 36944 63680 37264 64704
rect 36944 63616 36952 63680
rect 37016 63616 37032 63680
rect 37096 63616 37112 63680
rect 37176 63616 37192 63680
rect 37256 63616 37264 63680
rect 36944 63294 37264 63616
rect 36944 63058 36986 63294
rect 37222 63058 37264 63294
rect 36944 62592 37264 63058
rect 36944 62528 36952 62592
rect 37016 62528 37032 62592
rect 37096 62528 37112 62592
rect 37176 62528 37192 62592
rect 37256 62528 37264 62592
rect 36944 61504 37264 62528
rect 36944 61440 36952 61504
rect 37016 61440 37032 61504
rect 37096 61440 37112 61504
rect 37176 61440 37192 61504
rect 37256 61440 37264 61504
rect 36944 60416 37264 61440
rect 36944 60352 36952 60416
rect 37016 60352 37032 60416
rect 37096 60352 37112 60416
rect 37176 60352 37192 60416
rect 37256 60352 37264 60416
rect 36944 59328 37264 60352
rect 36944 59264 36952 59328
rect 37016 59264 37032 59328
rect 37096 59264 37112 59328
rect 37176 59264 37192 59328
rect 37256 59264 37264 59328
rect 33179 58308 33245 58309
rect 33179 58244 33180 58308
rect 33244 58244 33245 58308
rect 33179 58243 33245 58244
rect 36944 58294 37264 59264
rect 32604 57632 32612 57696
rect 32676 57632 32692 57696
rect 32756 57632 32772 57696
rect 32836 57632 32852 57696
rect 32916 57632 32924 57696
rect 32604 56608 32924 57632
rect 32604 56544 32612 56608
rect 32676 56544 32692 56608
rect 32756 56544 32772 56608
rect 32836 56544 32852 56608
rect 32916 56544 32924 56608
rect 32604 55520 32924 56544
rect 32604 55456 32612 55520
rect 32676 55456 32692 55520
rect 32756 55456 32772 55520
rect 32836 55456 32852 55520
rect 32916 55456 32924 55520
rect 32604 54432 32924 55456
rect 32604 54368 32612 54432
rect 32676 54368 32692 54432
rect 32756 54368 32772 54432
rect 32836 54368 32852 54432
rect 32916 54368 32924 54432
rect 32604 53954 32924 54368
rect 32604 53718 32646 53954
rect 32882 53718 32924 53954
rect 32604 53344 32924 53718
rect 32604 53280 32612 53344
rect 32676 53280 32692 53344
rect 32756 53280 32772 53344
rect 32836 53280 32852 53344
rect 32916 53280 32924 53344
rect 32604 52256 32924 53280
rect 32604 52192 32612 52256
rect 32676 52192 32692 52256
rect 32756 52192 32772 52256
rect 32836 52192 32852 52256
rect 32916 52192 32924 52256
rect 32604 51168 32924 52192
rect 32604 51104 32612 51168
rect 32676 51104 32692 51168
rect 32756 51104 32772 51168
rect 32836 51104 32852 51168
rect 32916 51104 32924 51168
rect 32443 50964 32509 50965
rect 32443 50900 32444 50964
rect 32508 50900 32509 50964
rect 32443 50899 32509 50900
rect 31944 50560 31952 50624
rect 32016 50560 32032 50624
rect 32096 50560 32112 50624
rect 32176 50560 32192 50624
rect 32256 50560 32264 50624
rect 31944 49536 32264 50560
rect 31944 49472 31952 49536
rect 32016 49472 32032 49536
rect 32096 49472 32112 49536
rect 32176 49472 32192 49536
rect 32256 49472 32264 49536
rect 31944 48448 32264 49472
rect 31944 48384 31952 48448
rect 32016 48384 32032 48448
rect 32096 48384 32112 48448
rect 32176 48384 32192 48448
rect 32256 48384 32264 48448
rect 31944 48294 32264 48384
rect 31944 48058 31986 48294
rect 32222 48058 32264 48294
rect 31944 47360 32264 48058
rect 31944 47296 31952 47360
rect 32016 47296 32032 47360
rect 32096 47296 32112 47360
rect 32176 47296 32192 47360
rect 32256 47296 32264 47360
rect 31944 46272 32264 47296
rect 31944 46208 31952 46272
rect 32016 46208 32032 46272
rect 32096 46208 32112 46272
rect 32176 46208 32192 46272
rect 32256 46208 32264 46272
rect 31944 45184 32264 46208
rect 31944 45120 31952 45184
rect 32016 45120 32032 45184
rect 32096 45120 32112 45184
rect 32176 45120 32192 45184
rect 32256 45120 32264 45184
rect 31944 44096 32264 45120
rect 31944 44032 31952 44096
rect 32016 44032 32032 44096
rect 32096 44032 32112 44096
rect 32176 44032 32192 44096
rect 32256 44032 32264 44096
rect 31944 43294 32264 44032
rect 31944 43058 31986 43294
rect 32222 43058 32264 43294
rect 31944 43008 32264 43058
rect 31944 42944 31952 43008
rect 32016 42944 32032 43008
rect 32096 42944 32112 43008
rect 32176 42944 32192 43008
rect 32256 42944 32264 43008
rect 31944 41920 32264 42944
rect 31944 41856 31952 41920
rect 32016 41856 32032 41920
rect 32096 41856 32112 41920
rect 32176 41856 32192 41920
rect 32256 41856 32264 41920
rect 31707 41444 31773 41445
rect 31707 41430 31708 41444
rect 27604 41312 27612 41376
rect 27676 41312 27692 41376
rect 27756 41312 27772 41376
rect 27836 41312 27852 41376
rect 27916 41312 27924 41376
rect 27604 40288 27924 41312
rect 27604 40224 27612 40288
rect 27676 40224 27692 40288
rect 27756 40224 27772 40288
rect 27836 40224 27852 40288
rect 27916 40224 27924 40288
rect 27604 39200 27924 40224
rect 27604 39136 27612 39200
rect 27676 39136 27692 39200
rect 27756 39136 27772 39200
rect 27836 39136 27852 39200
rect 27916 39136 27924 39200
rect 27604 38954 27924 39136
rect 27604 38718 27646 38954
rect 27882 38718 27924 38954
rect 27604 38112 27924 38718
rect 27604 38048 27612 38112
rect 27676 38048 27692 38112
rect 27756 38048 27772 38112
rect 27836 38048 27852 38112
rect 27916 38048 27924 38112
rect 27604 37024 27924 38048
rect 27604 36960 27612 37024
rect 27676 36960 27692 37024
rect 27756 36960 27772 37024
rect 27836 36960 27852 37024
rect 27916 36960 27924 37024
rect 27604 35936 27924 36960
rect 27604 35872 27612 35936
rect 27676 35872 27692 35936
rect 27756 35872 27772 35936
rect 27836 35872 27852 35936
rect 27916 35872 27924 35936
rect 27604 34848 27924 35872
rect 27604 34784 27612 34848
rect 27676 34784 27692 34848
rect 27756 34784 27772 34848
rect 27836 34784 27852 34848
rect 27916 34784 27924 34848
rect 27604 33954 27924 34784
rect 27604 33760 27646 33954
rect 27882 33760 27924 33954
rect 27604 33696 27612 33760
rect 27676 33696 27692 33718
rect 27756 33696 27772 33718
rect 27836 33696 27852 33718
rect 27916 33696 27924 33760
rect 27604 32672 27924 33696
rect 27604 32608 27612 32672
rect 27676 32608 27692 32672
rect 27756 32608 27772 32672
rect 27836 32608 27852 32672
rect 27916 32608 27924 32672
rect 27604 31584 27924 32608
rect 31526 41380 31708 41430
rect 31772 41380 31773 41444
rect 31526 41379 31773 41380
rect 31526 41370 31770 41379
rect 31526 31770 31586 41370
rect 31944 40832 32264 41856
rect 32446 41445 32506 50899
rect 32604 50080 32924 51104
rect 32604 50016 32612 50080
rect 32676 50016 32692 50080
rect 32756 50016 32772 50080
rect 32836 50016 32852 50080
rect 32916 50016 32924 50080
rect 32604 48992 32924 50016
rect 32604 48928 32612 48992
rect 32676 48954 32692 48992
rect 32756 48954 32772 48992
rect 32836 48954 32852 48992
rect 32916 48928 32924 48992
rect 32604 48718 32646 48928
rect 32882 48718 32924 48928
rect 32604 47904 32924 48718
rect 32604 47840 32612 47904
rect 32676 47840 32692 47904
rect 32756 47840 32772 47904
rect 32836 47840 32852 47904
rect 32916 47840 32924 47904
rect 32604 46816 32924 47840
rect 32604 46752 32612 46816
rect 32676 46752 32692 46816
rect 32756 46752 32772 46816
rect 32836 46752 32852 46816
rect 32916 46752 32924 46816
rect 32604 45728 32924 46752
rect 32604 45664 32612 45728
rect 32676 45664 32692 45728
rect 32756 45664 32772 45728
rect 32836 45664 32852 45728
rect 32916 45664 32924 45728
rect 32604 44640 32924 45664
rect 32604 44576 32612 44640
rect 32676 44576 32692 44640
rect 32756 44576 32772 44640
rect 32836 44576 32852 44640
rect 32916 44576 32924 44640
rect 32604 43954 32924 44576
rect 32604 43718 32646 43954
rect 32882 43718 32924 43954
rect 32604 43552 32924 43718
rect 32604 43488 32612 43552
rect 32676 43488 32692 43552
rect 32756 43488 32772 43552
rect 32836 43488 32852 43552
rect 32916 43488 32924 43552
rect 32604 42464 32924 43488
rect 32604 42400 32612 42464
rect 32676 42400 32692 42464
rect 32756 42400 32772 42464
rect 32836 42400 32852 42464
rect 32916 42400 32924 42464
rect 32443 41444 32509 41445
rect 32443 41380 32444 41444
rect 32508 41380 32509 41444
rect 32443 41379 32509 41380
rect 31944 40768 31952 40832
rect 32016 40768 32032 40832
rect 32096 40768 32112 40832
rect 32176 40768 32192 40832
rect 32256 40768 32264 40832
rect 31944 39744 32264 40768
rect 31944 39680 31952 39744
rect 32016 39680 32032 39744
rect 32096 39680 32112 39744
rect 32176 39680 32192 39744
rect 32256 39680 32264 39744
rect 31944 38656 32264 39680
rect 31944 38592 31952 38656
rect 32016 38592 32032 38656
rect 32096 38592 32112 38656
rect 32176 38592 32192 38656
rect 32256 38592 32264 38656
rect 31944 38294 32264 38592
rect 31944 38058 31986 38294
rect 32222 38058 32264 38294
rect 31944 37568 32264 38058
rect 31944 37504 31952 37568
rect 32016 37504 32032 37568
rect 32096 37504 32112 37568
rect 32176 37504 32192 37568
rect 32256 37504 32264 37568
rect 31944 36480 32264 37504
rect 31944 36416 31952 36480
rect 32016 36416 32032 36480
rect 32096 36416 32112 36480
rect 32176 36416 32192 36480
rect 32256 36416 32264 36480
rect 31944 35392 32264 36416
rect 31944 35328 31952 35392
rect 32016 35328 32032 35392
rect 32096 35328 32112 35392
rect 32176 35328 32192 35392
rect 32256 35328 32264 35392
rect 31944 34304 32264 35328
rect 31944 34240 31952 34304
rect 32016 34240 32032 34304
rect 32096 34240 32112 34304
rect 32176 34240 32192 34304
rect 32256 34240 32264 34304
rect 31944 33294 32264 34240
rect 31944 33216 31986 33294
rect 32222 33216 32264 33294
rect 31944 33152 31952 33216
rect 32256 33152 32264 33216
rect 31944 33058 31986 33152
rect 32222 33058 32264 33152
rect 31944 32128 32264 33058
rect 31944 32064 31952 32128
rect 32016 32064 32032 32128
rect 32096 32064 32112 32128
rect 32176 32064 32192 32128
rect 32256 32064 32264 32128
rect 31526 31710 31770 31770
rect 27604 31520 27612 31584
rect 27676 31520 27692 31584
rect 27756 31520 27772 31584
rect 27836 31520 27852 31584
rect 27916 31520 27924 31584
rect 27604 30496 27924 31520
rect 27604 30432 27612 30496
rect 27676 30432 27692 30496
rect 27756 30432 27772 30496
rect 27836 30432 27852 30496
rect 27916 30432 27924 30496
rect 27604 29408 27924 30432
rect 27604 29344 27612 29408
rect 27676 29344 27692 29408
rect 27756 29344 27772 29408
rect 27836 29344 27852 29408
rect 27916 29344 27924 29408
rect 27604 28954 27924 29344
rect 27604 28718 27646 28954
rect 27882 28718 27924 28954
rect 31710 28797 31770 31710
rect 31944 31040 32264 32064
rect 31944 30976 31952 31040
rect 32016 30976 32032 31040
rect 32096 30976 32112 31040
rect 32176 30976 32192 31040
rect 32256 30976 32264 31040
rect 31944 29952 32264 30976
rect 31944 29888 31952 29952
rect 32016 29888 32032 29952
rect 32096 29888 32112 29952
rect 32176 29888 32192 29952
rect 32256 29888 32264 29952
rect 31944 28864 32264 29888
rect 31944 28800 31952 28864
rect 32016 28800 32032 28864
rect 32096 28800 32112 28864
rect 32176 28800 32192 28864
rect 32256 28800 32264 28864
rect 31707 28796 31773 28797
rect 31707 28732 31708 28796
rect 31772 28732 31773 28796
rect 31707 28731 31773 28732
rect 27604 28320 27924 28718
rect 27604 28256 27612 28320
rect 27676 28256 27692 28320
rect 27756 28256 27772 28320
rect 27836 28256 27852 28320
rect 27916 28256 27924 28320
rect 27604 27232 27924 28256
rect 27604 27168 27612 27232
rect 27676 27168 27692 27232
rect 27756 27168 27772 27232
rect 27836 27168 27852 27232
rect 27916 27168 27924 27232
rect 27604 26144 27924 27168
rect 27604 26080 27612 26144
rect 27676 26080 27692 26144
rect 27756 26080 27772 26144
rect 27836 26080 27852 26144
rect 27916 26080 27924 26144
rect 27604 25056 27924 26080
rect 27604 24992 27612 25056
rect 27676 24992 27692 25056
rect 27756 24992 27772 25056
rect 27836 24992 27852 25056
rect 27916 24992 27924 25056
rect 27604 23968 27924 24992
rect 27604 23904 27612 23968
rect 27676 23954 27692 23968
rect 27756 23954 27772 23968
rect 27836 23954 27852 23968
rect 27916 23904 27924 23968
rect 27604 23718 27646 23904
rect 27882 23718 27924 23904
rect 27604 22880 27924 23718
rect 27604 22816 27612 22880
rect 27676 22816 27692 22880
rect 27756 22816 27772 22880
rect 27836 22816 27852 22880
rect 27916 22816 27924 22880
rect 27604 21792 27924 22816
rect 27604 21728 27612 21792
rect 27676 21728 27692 21792
rect 27756 21728 27772 21792
rect 27836 21728 27852 21792
rect 27916 21728 27924 21792
rect 27604 20704 27924 21728
rect 27604 20640 27612 20704
rect 27676 20640 27692 20704
rect 27756 20640 27772 20704
rect 27836 20640 27852 20704
rect 27916 20640 27924 20704
rect 27604 19616 27924 20640
rect 27604 19552 27612 19616
rect 27676 19552 27692 19616
rect 27756 19552 27772 19616
rect 27836 19552 27852 19616
rect 27916 19552 27924 19616
rect 27604 18954 27924 19552
rect 27604 18718 27646 18954
rect 27882 18718 27924 18954
rect 27604 18528 27924 18718
rect 27604 18464 27612 18528
rect 27676 18464 27692 18528
rect 27756 18464 27772 18528
rect 27836 18464 27852 18528
rect 27916 18464 27924 18528
rect 27604 17440 27924 18464
rect 27604 17376 27612 17440
rect 27676 17376 27692 17440
rect 27756 17376 27772 17440
rect 27836 17376 27852 17440
rect 27916 17376 27924 17440
rect 27604 16352 27924 17376
rect 27604 16288 27612 16352
rect 27676 16288 27692 16352
rect 27756 16288 27772 16352
rect 27836 16288 27852 16352
rect 27916 16288 27924 16352
rect 27604 15264 27924 16288
rect 27604 15200 27612 15264
rect 27676 15200 27692 15264
rect 27756 15200 27772 15264
rect 27836 15200 27852 15264
rect 27916 15200 27924 15264
rect 27604 14176 27924 15200
rect 27604 14112 27612 14176
rect 27676 14112 27692 14176
rect 27756 14112 27772 14176
rect 27836 14112 27852 14176
rect 27916 14112 27924 14176
rect 27604 13954 27924 14112
rect 27604 13718 27646 13954
rect 27882 13718 27924 13954
rect 27604 13088 27924 13718
rect 27604 13024 27612 13088
rect 27676 13024 27692 13088
rect 27756 13024 27772 13088
rect 27836 13024 27852 13088
rect 27916 13024 27924 13088
rect 27604 12000 27924 13024
rect 27604 11936 27612 12000
rect 27676 11936 27692 12000
rect 27756 11936 27772 12000
rect 27836 11936 27852 12000
rect 27916 11936 27924 12000
rect 27604 10912 27924 11936
rect 27604 10848 27612 10912
rect 27676 10848 27692 10912
rect 27756 10848 27772 10912
rect 27836 10848 27852 10912
rect 27916 10848 27924 10912
rect 27604 9824 27924 10848
rect 27604 9760 27612 9824
rect 27676 9760 27692 9824
rect 27756 9760 27772 9824
rect 27836 9760 27852 9824
rect 27916 9760 27924 9824
rect 27604 8954 27924 9760
rect 27604 8736 27646 8954
rect 27882 8736 27924 8954
rect 27604 8672 27612 8736
rect 27676 8672 27692 8718
rect 27756 8672 27772 8718
rect 27836 8672 27852 8718
rect 27916 8672 27924 8736
rect 27604 7648 27924 8672
rect 27604 7584 27612 7648
rect 27676 7584 27692 7648
rect 27756 7584 27772 7648
rect 27836 7584 27852 7648
rect 27916 7584 27924 7648
rect 27604 6560 27924 7584
rect 27604 6496 27612 6560
rect 27676 6496 27692 6560
rect 27756 6496 27772 6560
rect 27836 6496 27852 6560
rect 27916 6496 27924 6560
rect 27604 5472 27924 6496
rect 27604 5408 27612 5472
rect 27676 5408 27692 5472
rect 27756 5408 27772 5472
rect 27836 5408 27852 5472
rect 27916 5408 27924 5472
rect 27604 4384 27924 5408
rect 27604 4320 27612 4384
rect 27676 4320 27692 4384
rect 27756 4320 27772 4384
rect 27836 4320 27852 4384
rect 27916 4320 27924 4384
rect 27604 3954 27924 4320
rect 27604 3718 27646 3954
rect 27882 3718 27924 3954
rect 27604 3296 27924 3718
rect 27604 3232 27612 3296
rect 27676 3232 27692 3296
rect 27756 3232 27772 3296
rect 27836 3232 27852 3296
rect 27916 3232 27924 3296
rect 27604 2208 27924 3232
rect 27604 2144 27612 2208
rect 27676 2144 27692 2208
rect 27756 2144 27772 2208
rect 27836 2144 27852 2208
rect 27916 2144 27924 2208
rect 27604 2128 27924 2144
rect 31944 28294 32264 28800
rect 31944 28058 31986 28294
rect 32222 28058 32264 28294
rect 31944 27776 32264 28058
rect 31944 27712 31952 27776
rect 32016 27712 32032 27776
rect 32096 27712 32112 27776
rect 32176 27712 32192 27776
rect 32256 27712 32264 27776
rect 31944 26688 32264 27712
rect 31944 26624 31952 26688
rect 32016 26624 32032 26688
rect 32096 26624 32112 26688
rect 32176 26624 32192 26688
rect 32256 26624 32264 26688
rect 31944 25600 32264 26624
rect 31944 25536 31952 25600
rect 32016 25536 32032 25600
rect 32096 25536 32112 25600
rect 32176 25536 32192 25600
rect 32256 25536 32264 25600
rect 31944 24512 32264 25536
rect 31944 24448 31952 24512
rect 32016 24448 32032 24512
rect 32096 24448 32112 24512
rect 32176 24448 32192 24512
rect 32256 24448 32264 24512
rect 31944 23424 32264 24448
rect 31944 23360 31952 23424
rect 32016 23360 32032 23424
rect 32096 23360 32112 23424
rect 32176 23360 32192 23424
rect 32256 23360 32264 23424
rect 31944 23294 32264 23360
rect 31944 23058 31986 23294
rect 32222 23058 32264 23294
rect 31944 22336 32264 23058
rect 31944 22272 31952 22336
rect 32016 22272 32032 22336
rect 32096 22272 32112 22336
rect 32176 22272 32192 22336
rect 32256 22272 32264 22336
rect 31944 21248 32264 22272
rect 31944 21184 31952 21248
rect 32016 21184 32032 21248
rect 32096 21184 32112 21248
rect 32176 21184 32192 21248
rect 32256 21184 32264 21248
rect 31944 20160 32264 21184
rect 31944 20096 31952 20160
rect 32016 20096 32032 20160
rect 32096 20096 32112 20160
rect 32176 20096 32192 20160
rect 32256 20096 32264 20160
rect 31944 19072 32264 20096
rect 31944 19008 31952 19072
rect 32016 19008 32032 19072
rect 32096 19008 32112 19072
rect 32176 19008 32192 19072
rect 32256 19008 32264 19072
rect 31944 18294 32264 19008
rect 31944 18058 31986 18294
rect 32222 18058 32264 18294
rect 31944 17984 32264 18058
rect 31944 17920 31952 17984
rect 32016 17920 32032 17984
rect 32096 17920 32112 17984
rect 32176 17920 32192 17984
rect 32256 17920 32264 17984
rect 31944 16896 32264 17920
rect 31944 16832 31952 16896
rect 32016 16832 32032 16896
rect 32096 16832 32112 16896
rect 32176 16832 32192 16896
rect 32256 16832 32264 16896
rect 31944 15808 32264 16832
rect 31944 15744 31952 15808
rect 32016 15744 32032 15808
rect 32096 15744 32112 15808
rect 32176 15744 32192 15808
rect 32256 15744 32264 15808
rect 31944 14720 32264 15744
rect 31944 14656 31952 14720
rect 32016 14656 32032 14720
rect 32096 14656 32112 14720
rect 32176 14656 32192 14720
rect 32256 14656 32264 14720
rect 31944 13632 32264 14656
rect 31944 13568 31952 13632
rect 32016 13568 32032 13632
rect 32096 13568 32112 13632
rect 32176 13568 32192 13632
rect 32256 13568 32264 13632
rect 31944 13294 32264 13568
rect 31944 13058 31986 13294
rect 32222 13058 32264 13294
rect 31944 12544 32264 13058
rect 31944 12480 31952 12544
rect 32016 12480 32032 12544
rect 32096 12480 32112 12544
rect 32176 12480 32192 12544
rect 32256 12480 32264 12544
rect 31944 11456 32264 12480
rect 31944 11392 31952 11456
rect 32016 11392 32032 11456
rect 32096 11392 32112 11456
rect 32176 11392 32192 11456
rect 32256 11392 32264 11456
rect 31944 10368 32264 11392
rect 31944 10304 31952 10368
rect 32016 10304 32032 10368
rect 32096 10304 32112 10368
rect 32176 10304 32192 10368
rect 32256 10304 32264 10368
rect 31944 9280 32264 10304
rect 31944 9216 31952 9280
rect 32016 9216 32032 9280
rect 32096 9216 32112 9280
rect 32176 9216 32192 9280
rect 32256 9216 32264 9280
rect 31944 8294 32264 9216
rect 31944 8192 31986 8294
rect 32222 8192 32264 8294
rect 31944 8128 31952 8192
rect 32256 8128 32264 8192
rect 31944 8058 31986 8128
rect 32222 8058 32264 8128
rect 31944 7104 32264 8058
rect 31944 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32264 7104
rect 31944 6016 32264 7040
rect 31944 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32264 6016
rect 31944 4928 32264 5952
rect 31944 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32264 4928
rect 31944 3840 32264 4864
rect 31944 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32264 3840
rect 31944 3294 32264 3776
rect 31944 3058 31986 3294
rect 32222 3058 32264 3294
rect 31944 2752 32264 3058
rect 31944 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32264 2752
rect 31944 2128 32264 2688
rect 32604 41376 32924 42400
rect 32604 41312 32612 41376
rect 32676 41312 32692 41376
rect 32756 41312 32772 41376
rect 32836 41312 32852 41376
rect 32916 41312 32924 41376
rect 32604 40288 32924 41312
rect 32604 40224 32612 40288
rect 32676 40224 32692 40288
rect 32756 40224 32772 40288
rect 32836 40224 32852 40288
rect 32916 40224 32924 40288
rect 32604 39200 32924 40224
rect 32604 39136 32612 39200
rect 32676 39136 32692 39200
rect 32756 39136 32772 39200
rect 32836 39136 32852 39200
rect 32916 39136 32924 39200
rect 32604 38954 32924 39136
rect 32604 38718 32646 38954
rect 32882 38718 32924 38954
rect 32604 38112 32924 38718
rect 32604 38048 32612 38112
rect 32676 38048 32692 38112
rect 32756 38048 32772 38112
rect 32836 38048 32852 38112
rect 32916 38048 32924 38112
rect 32604 37024 32924 38048
rect 32604 36960 32612 37024
rect 32676 36960 32692 37024
rect 32756 36960 32772 37024
rect 32836 36960 32852 37024
rect 32916 36960 32924 37024
rect 32604 35936 32924 36960
rect 32604 35872 32612 35936
rect 32676 35872 32692 35936
rect 32756 35872 32772 35936
rect 32836 35872 32852 35936
rect 32916 35872 32924 35936
rect 32604 34848 32924 35872
rect 32604 34784 32612 34848
rect 32676 34784 32692 34848
rect 32756 34784 32772 34848
rect 32836 34784 32852 34848
rect 32916 34784 32924 34848
rect 32604 33954 32924 34784
rect 32604 33760 32646 33954
rect 32882 33760 32924 33954
rect 32604 33696 32612 33760
rect 32676 33696 32692 33718
rect 32756 33696 32772 33718
rect 32836 33696 32852 33718
rect 32916 33696 32924 33760
rect 32604 32672 32924 33696
rect 32604 32608 32612 32672
rect 32676 32608 32692 32672
rect 32756 32608 32772 32672
rect 32836 32608 32852 32672
rect 32916 32608 32924 32672
rect 32604 31584 32924 32608
rect 32604 31520 32612 31584
rect 32676 31520 32692 31584
rect 32756 31520 32772 31584
rect 32836 31520 32852 31584
rect 32916 31520 32924 31584
rect 32604 30496 32924 31520
rect 32604 30432 32612 30496
rect 32676 30432 32692 30496
rect 32756 30432 32772 30496
rect 32836 30432 32852 30496
rect 32916 30432 32924 30496
rect 32604 29408 32924 30432
rect 32604 29344 32612 29408
rect 32676 29344 32692 29408
rect 32756 29344 32772 29408
rect 32836 29344 32852 29408
rect 32916 29344 32924 29408
rect 32604 28954 32924 29344
rect 32604 28718 32646 28954
rect 32882 28718 32924 28954
rect 32604 28320 32924 28718
rect 32604 28256 32612 28320
rect 32676 28256 32692 28320
rect 32756 28256 32772 28320
rect 32836 28256 32852 28320
rect 32916 28256 32924 28320
rect 32604 27232 32924 28256
rect 32604 27168 32612 27232
rect 32676 27168 32692 27232
rect 32756 27168 32772 27232
rect 32836 27168 32852 27232
rect 32916 27168 32924 27232
rect 32604 26144 32924 27168
rect 32604 26080 32612 26144
rect 32676 26080 32692 26144
rect 32756 26080 32772 26144
rect 32836 26080 32852 26144
rect 32916 26080 32924 26144
rect 32604 25056 32924 26080
rect 32604 24992 32612 25056
rect 32676 24992 32692 25056
rect 32756 24992 32772 25056
rect 32836 24992 32852 25056
rect 32916 24992 32924 25056
rect 32604 23968 32924 24992
rect 32604 23904 32612 23968
rect 32676 23954 32692 23968
rect 32756 23954 32772 23968
rect 32836 23954 32852 23968
rect 32916 23904 32924 23968
rect 32604 23718 32646 23904
rect 32882 23718 32924 23904
rect 32604 22880 32924 23718
rect 32604 22816 32612 22880
rect 32676 22816 32692 22880
rect 32756 22816 32772 22880
rect 32836 22816 32852 22880
rect 32916 22816 32924 22880
rect 32604 21792 32924 22816
rect 32604 21728 32612 21792
rect 32676 21728 32692 21792
rect 32756 21728 32772 21792
rect 32836 21728 32852 21792
rect 32916 21728 32924 21792
rect 32604 20704 32924 21728
rect 32604 20640 32612 20704
rect 32676 20640 32692 20704
rect 32756 20640 32772 20704
rect 32836 20640 32852 20704
rect 32916 20640 32924 20704
rect 32604 19616 32924 20640
rect 32604 19552 32612 19616
rect 32676 19552 32692 19616
rect 32756 19552 32772 19616
rect 32836 19552 32852 19616
rect 32916 19552 32924 19616
rect 32604 18954 32924 19552
rect 32604 18718 32646 18954
rect 32882 18718 32924 18954
rect 32604 18528 32924 18718
rect 32604 18464 32612 18528
rect 32676 18464 32692 18528
rect 32756 18464 32772 18528
rect 32836 18464 32852 18528
rect 32916 18464 32924 18528
rect 32604 17440 32924 18464
rect 32604 17376 32612 17440
rect 32676 17376 32692 17440
rect 32756 17376 32772 17440
rect 32836 17376 32852 17440
rect 32916 17376 32924 17440
rect 32604 16352 32924 17376
rect 32604 16288 32612 16352
rect 32676 16288 32692 16352
rect 32756 16288 32772 16352
rect 32836 16288 32852 16352
rect 32916 16288 32924 16352
rect 32604 15264 32924 16288
rect 32604 15200 32612 15264
rect 32676 15200 32692 15264
rect 32756 15200 32772 15264
rect 32836 15200 32852 15264
rect 32916 15200 32924 15264
rect 32604 14176 32924 15200
rect 32604 14112 32612 14176
rect 32676 14112 32692 14176
rect 32756 14112 32772 14176
rect 32836 14112 32852 14176
rect 32916 14112 32924 14176
rect 32604 13954 32924 14112
rect 32604 13718 32646 13954
rect 32882 13718 32924 13954
rect 32604 13088 32924 13718
rect 32604 13024 32612 13088
rect 32676 13024 32692 13088
rect 32756 13024 32772 13088
rect 32836 13024 32852 13088
rect 32916 13024 32924 13088
rect 32604 12000 32924 13024
rect 32604 11936 32612 12000
rect 32676 11936 32692 12000
rect 32756 11936 32772 12000
rect 32836 11936 32852 12000
rect 32916 11936 32924 12000
rect 32604 10912 32924 11936
rect 33182 10981 33242 58243
rect 36944 58240 36986 58294
rect 37222 58240 37264 58294
rect 36944 58176 36952 58240
rect 37256 58176 37264 58240
rect 36944 58058 36986 58176
rect 37222 58058 37264 58176
rect 36944 57152 37264 58058
rect 36944 57088 36952 57152
rect 37016 57088 37032 57152
rect 37096 57088 37112 57152
rect 37176 57088 37192 57152
rect 37256 57088 37264 57152
rect 36944 56064 37264 57088
rect 36944 56000 36952 56064
rect 37016 56000 37032 56064
rect 37096 56000 37112 56064
rect 37176 56000 37192 56064
rect 37256 56000 37264 56064
rect 33915 55860 33981 55861
rect 33915 55796 33916 55860
rect 33980 55796 33981 55860
rect 33915 55795 33981 55796
rect 33547 55724 33613 55725
rect 33547 55660 33548 55724
rect 33612 55660 33613 55724
rect 33547 55659 33613 55660
rect 33363 51236 33429 51237
rect 33363 51172 33364 51236
rect 33428 51172 33429 51236
rect 33363 51171 33429 51172
rect 33179 10980 33245 10981
rect 33179 10916 33180 10980
rect 33244 10916 33245 10980
rect 33179 10915 33245 10916
rect 32604 10848 32612 10912
rect 32676 10848 32692 10912
rect 32756 10848 32772 10912
rect 32836 10848 32852 10912
rect 32916 10848 32924 10912
rect 32604 9824 32924 10848
rect 32604 9760 32612 9824
rect 32676 9760 32692 9824
rect 32756 9760 32772 9824
rect 32836 9760 32852 9824
rect 32916 9760 32924 9824
rect 32604 8954 32924 9760
rect 33366 9621 33426 51171
rect 33363 9620 33429 9621
rect 33363 9556 33364 9620
rect 33428 9556 33429 9620
rect 33363 9555 33429 9556
rect 32604 8736 32646 8954
rect 32882 8736 32924 8954
rect 32604 8672 32612 8736
rect 32676 8672 32692 8718
rect 32756 8672 32772 8718
rect 32836 8672 32852 8718
rect 32916 8672 32924 8736
rect 32604 7648 32924 8672
rect 33550 7853 33610 55659
rect 33918 14381 33978 55795
rect 36944 54976 37264 56000
rect 36944 54912 36952 54976
rect 37016 54912 37032 54976
rect 37096 54912 37112 54976
rect 37176 54912 37192 54976
rect 37256 54912 37264 54976
rect 36944 53888 37264 54912
rect 36944 53824 36952 53888
rect 37016 53824 37032 53888
rect 37096 53824 37112 53888
rect 37176 53824 37192 53888
rect 37256 53824 37264 53888
rect 36944 53294 37264 53824
rect 36944 53058 36986 53294
rect 37222 53058 37264 53294
rect 36944 52800 37264 53058
rect 36944 52736 36952 52800
rect 37016 52736 37032 52800
rect 37096 52736 37112 52800
rect 37176 52736 37192 52800
rect 37256 52736 37264 52800
rect 36944 51712 37264 52736
rect 36944 51648 36952 51712
rect 37016 51648 37032 51712
rect 37096 51648 37112 51712
rect 37176 51648 37192 51712
rect 37256 51648 37264 51712
rect 36944 50624 37264 51648
rect 36944 50560 36952 50624
rect 37016 50560 37032 50624
rect 37096 50560 37112 50624
rect 37176 50560 37192 50624
rect 37256 50560 37264 50624
rect 36944 49536 37264 50560
rect 36944 49472 36952 49536
rect 37016 49472 37032 49536
rect 37096 49472 37112 49536
rect 37176 49472 37192 49536
rect 37256 49472 37264 49536
rect 36944 48448 37264 49472
rect 36944 48384 36952 48448
rect 37016 48384 37032 48448
rect 37096 48384 37112 48448
rect 37176 48384 37192 48448
rect 37256 48384 37264 48448
rect 36944 48294 37264 48384
rect 36944 48058 36986 48294
rect 37222 48058 37264 48294
rect 36944 47360 37264 48058
rect 36944 47296 36952 47360
rect 37016 47296 37032 47360
rect 37096 47296 37112 47360
rect 37176 47296 37192 47360
rect 37256 47296 37264 47360
rect 36944 46272 37264 47296
rect 36944 46208 36952 46272
rect 37016 46208 37032 46272
rect 37096 46208 37112 46272
rect 37176 46208 37192 46272
rect 37256 46208 37264 46272
rect 36944 45184 37264 46208
rect 36944 45120 36952 45184
rect 37016 45120 37032 45184
rect 37096 45120 37112 45184
rect 37176 45120 37192 45184
rect 37256 45120 37264 45184
rect 36944 44096 37264 45120
rect 36944 44032 36952 44096
rect 37016 44032 37032 44096
rect 37096 44032 37112 44096
rect 37176 44032 37192 44096
rect 37256 44032 37264 44096
rect 36944 43294 37264 44032
rect 36944 43058 36986 43294
rect 37222 43058 37264 43294
rect 36944 43008 37264 43058
rect 36944 42944 36952 43008
rect 37016 42944 37032 43008
rect 37096 42944 37112 43008
rect 37176 42944 37192 43008
rect 37256 42944 37264 43008
rect 36944 41920 37264 42944
rect 36944 41856 36952 41920
rect 37016 41856 37032 41920
rect 37096 41856 37112 41920
rect 37176 41856 37192 41920
rect 37256 41856 37264 41920
rect 36944 40832 37264 41856
rect 36944 40768 36952 40832
rect 37016 40768 37032 40832
rect 37096 40768 37112 40832
rect 37176 40768 37192 40832
rect 37256 40768 37264 40832
rect 36944 39744 37264 40768
rect 36944 39680 36952 39744
rect 37016 39680 37032 39744
rect 37096 39680 37112 39744
rect 37176 39680 37192 39744
rect 37256 39680 37264 39744
rect 36944 38656 37264 39680
rect 36944 38592 36952 38656
rect 37016 38592 37032 38656
rect 37096 38592 37112 38656
rect 37176 38592 37192 38656
rect 37256 38592 37264 38656
rect 36944 38294 37264 38592
rect 36944 38058 36986 38294
rect 37222 38058 37264 38294
rect 36944 37568 37264 38058
rect 36944 37504 36952 37568
rect 37016 37504 37032 37568
rect 37096 37504 37112 37568
rect 37176 37504 37192 37568
rect 37256 37504 37264 37568
rect 36944 36480 37264 37504
rect 36944 36416 36952 36480
rect 37016 36416 37032 36480
rect 37096 36416 37112 36480
rect 37176 36416 37192 36480
rect 37256 36416 37264 36480
rect 36944 35392 37264 36416
rect 36944 35328 36952 35392
rect 37016 35328 37032 35392
rect 37096 35328 37112 35392
rect 37176 35328 37192 35392
rect 37256 35328 37264 35392
rect 36944 34304 37264 35328
rect 36944 34240 36952 34304
rect 37016 34240 37032 34304
rect 37096 34240 37112 34304
rect 37176 34240 37192 34304
rect 37256 34240 37264 34304
rect 36944 33294 37264 34240
rect 36944 33216 36986 33294
rect 37222 33216 37264 33294
rect 36944 33152 36952 33216
rect 37256 33152 37264 33216
rect 36944 33058 36986 33152
rect 37222 33058 37264 33152
rect 36944 32128 37264 33058
rect 36944 32064 36952 32128
rect 37016 32064 37032 32128
rect 37096 32064 37112 32128
rect 37176 32064 37192 32128
rect 37256 32064 37264 32128
rect 36944 31040 37264 32064
rect 36944 30976 36952 31040
rect 37016 30976 37032 31040
rect 37096 30976 37112 31040
rect 37176 30976 37192 31040
rect 37256 30976 37264 31040
rect 36944 29952 37264 30976
rect 36944 29888 36952 29952
rect 37016 29888 37032 29952
rect 37096 29888 37112 29952
rect 37176 29888 37192 29952
rect 37256 29888 37264 29952
rect 36944 28864 37264 29888
rect 36944 28800 36952 28864
rect 37016 28800 37032 28864
rect 37096 28800 37112 28864
rect 37176 28800 37192 28864
rect 37256 28800 37264 28864
rect 36944 28294 37264 28800
rect 36944 28058 36986 28294
rect 37222 28058 37264 28294
rect 36944 27776 37264 28058
rect 36944 27712 36952 27776
rect 37016 27712 37032 27776
rect 37096 27712 37112 27776
rect 37176 27712 37192 27776
rect 37256 27712 37264 27776
rect 36944 26688 37264 27712
rect 36944 26624 36952 26688
rect 37016 26624 37032 26688
rect 37096 26624 37112 26688
rect 37176 26624 37192 26688
rect 37256 26624 37264 26688
rect 36944 25600 37264 26624
rect 36944 25536 36952 25600
rect 37016 25536 37032 25600
rect 37096 25536 37112 25600
rect 37176 25536 37192 25600
rect 37256 25536 37264 25600
rect 36944 24512 37264 25536
rect 36944 24448 36952 24512
rect 37016 24448 37032 24512
rect 37096 24448 37112 24512
rect 37176 24448 37192 24512
rect 37256 24448 37264 24512
rect 36944 23424 37264 24448
rect 36944 23360 36952 23424
rect 37016 23360 37032 23424
rect 37096 23360 37112 23424
rect 37176 23360 37192 23424
rect 37256 23360 37264 23424
rect 36944 23294 37264 23360
rect 36944 23058 36986 23294
rect 37222 23058 37264 23294
rect 36944 22336 37264 23058
rect 36944 22272 36952 22336
rect 37016 22272 37032 22336
rect 37096 22272 37112 22336
rect 37176 22272 37192 22336
rect 37256 22272 37264 22336
rect 36944 21248 37264 22272
rect 36944 21184 36952 21248
rect 37016 21184 37032 21248
rect 37096 21184 37112 21248
rect 37176 21184 37192 21248
rect 37256 21184 37264 21248
rect 36944 20160 37264 21184
rect 36944 20096 36952 20160
rect 37016 20096 37032 20160
rect 37096 20096 37112 20160
rect 37176 20096 37192 20160
rect 37256 20096 37264 20160
rect 36944 19072 37264 20096
rect 36944 19008 36952 19072
rect 37016 19008 37032 19072
rect 37096 19008 37112 19072
rect 37176 19008 37192 19072
rect 37256 19008 37264 19072
rect 36944 18294 37264 19008
rect 36944 18058 36986 18294
rect 37222 18058 37264 18294
rect 36944 17984 37264 18058
rect 36944 17920 36952 17984
rect 37016 17920 37032 17984
rect 37096 17920 37112 17984
rect 37176 17920 37192 17984
rect 37256 17920 37264 17984
rect 36944 16896 37264 17920
rect 36944 16832 36952 16896
rect 37016 16832 37032 16896
rect 37096 16832 37112 16896
rect 37176 16832 37192 16896
rect 37256 16832 37264 16896
rect 36944 15808 37264 16832
rect 36944 15744 36952 15808
rect 37016 15744 37032 15808
rect 37096 15744 37112 15808
rect 37176 15744 37192 15808
rect 37256 15744 37264 15808
rect 36944 14720 37264 15744
rect 36944 14656 36952 14720
rect 37016 14656 37032 14720
rect 37096 14656 37112 14720
rect 37176 14656 37192 14720
rect 37256 14656 37264 14720
rect 33915 14380 33981 14381
rect 33915 14316 33916 14380
rect 33980 14316 33981 14380
rect 33915 14315 33981 14316
rect 36944 13632 37264 14656
rect 36944 13568 36952 13632
rect 37016 13568 37032 13632
rect 37096 13568 37112 13632
rect 37176 13568 37192 13632
rect 37256 13568 37264 13632
rect 36944 13294 37264 13568
rect 36944 13058 36986 13294
rect 37222 13058 37264 13294
rect 36944 12544 37264 13058
rect 36944 12480 36952 12544
rect 37016 12480 37032 12544
rect 37096 12480 37112 12544
rect 37176 12480 37192 12544
rect 37256 12480 37264 12544
rect 36944 11456 37264 12480
rect 36944 11392 36952 11456
rect 37016 11392 37032 11456
rect 37096 11392 37112 11456
rect 37176 11392 37192 11456
rect 37256 11392 37264 11456
rect 36944 10368 37264 11392
rect 36944 10304 36952 10368
rect 37016 10304 37032 10368
rect 37096 10304 37112 10368
rect 37176 10304 37192 10368
rect 37256 10304 37264 10368
rect 36944 9280 37264 10304
rect 36944 9216 36952 9280
rect 37016 9216 37032 9280
rect 37096 9216 37112 9280
rect 37176 9216 37192 9280
rect 37256 9216 37264 9280
rect 36944 8294 37264 9216
rect 36944 8192 36986 8294
rect 37222 8192 37264 8294
rect 36944 8128 36952 8192
rect 37256 8128 37264 8192
rect 36944 8058 36986 8128
rect 37222 8058 37264 8128
rect 33547 7852 33613 7853
rect 33547 7788 33548 7852
rect 33612 7788 33613 7852
rect 33547 7787 33613 7788
rect 32604 7584 32612 7648
rect 32676 7584 32692 7648
rect 32756 7584 32772 7648
rect 32836 7584 32852 7648
rect 32916 7584 32924 7648
rect 32604 6560 32924 7584
rect 32604 6496 32612 6560
rect 32676 6496 32692 6560
rect 32756 6496 32772 6560
rect 32836 6496 32852 6560
rect 32916 6496 32924 6560
rect 32604 5472 32924 6496
rect 32604 5408 32612 5472
rect 32676 5408 32692 5472
rect 32756 5408 32772 5472
rect 32836 5408 32852 5472
rect 32916 5408 32924 5472
rect 32604 4384 32924 5408
rect 32604 4320 32612 4384
rect 32676 4320 32692 4384
rect 32756 4320 32772 4384
rect 32836 4320 32852 4384
rect 32916 4320 32924 4384
rect 32604 3954 32924 4320
rect 32604 3718 32646 3954
rect 32882 3718 32924 3954
rect 32604 3296 32924 3718
rect 32604 3232 32612 3296
rect 32676 3232 32692 3296
rect 32756 3232 32772 3296
rect 32836 3232 32852 3296
rect 32916 3232 32924 3296
rect 32604 2208 32924 3232
rect 32604 2144 32612 2208
rect 32676 2144 32692 2208
rect 32756 2144 32772 2208
rect 32836 2144 32852 2208
rect 32916 2144 32924 2208
rect 32604 2128 32924 2144
rect 36944 7104 37264 8058
rect 36944 7040 36952 7104
rect 37016 7040 37032 7104
rect 37096 7040 37112 7104
rect 37176 7040 37192 7104
rect 37256 7040 37264 7104
rect 36944 6016 37264 7040
rect 36944 5952 36952 6016
rect 37016 5952 37032 6016
rect 37096 5952 37112 6016
rect 37176 5952 37192 6016
rect 37256 5952 37264 6016
rect 36944 4928 37264 5952
rect 36944 4864 36952 4928
rect 37016 4864 37032 4928
rect 37096 4864 37112 4928
rect 37176 4864 37192 4928
rect 37256 4864 37264 4928
rect 36944 3840 37264 4864
rect 36944 3776 36952 3840
rect 37016 3776 37032 3840
rect 37096 3776 37112 3840
rect 37176 3776 37192 3840
rect 37256 3776 37264 3840
rect 36944 3294 37264 3776
rect 36944 3058 36986 3294
rect 37222 3058 37264 3294
rect 36944 2752 37264 3058
rect 36944 2688 36952 2752
rect 37016 2688 37032 2752
rect 37096 2688 37112 2752
rect 37176 2688 37192 2752
rect 37256 2688 37264 2752
rect 36944 2128 37264 2688
rect 37604 69664 37924 69680
rect 37604 69600 37612 69664
rect 37676 69600 37692 69664
rect 37756 69600 37772 69664
rect 37836 69600 37852 69664
rect 37916 69600 37924 69664
rect 37604 68954 37924 69600
rect 37604 68718 37646 68954
rect 37882 68718 37924 68954
rect 37604 68576 37924 68718
rect 37604 68512 37612 68576
rect 37676 68512 37692 68576
rect 37756 68512 37772 68576
rect 37836 68512 37852 68576
rect 37916 68512 37924 68576
rect 37604 67488 37924 68512
rect 37604 67424 37612 67488
rect 37676 67424 37692 67488
rect 37756 67424 37772 67488
rect 37836 67424 37852 67488
rect 37916 67424 37924 67488
rect 37604 66400 37924 67424
rect 37604 66336 37612 66400
rect 37676 66336 37692 66400
rect 37756 66336 37772 66400
rect 37836 66336 37852 66400
rect 37916 66336 37924 66400
rect 37604 65312 37924 66336
rect 37604 65248 37612 65312
rect 37676 65248 37692 65312
rect 37756 65248 37772 65312
rect 37836 65248 37852 65312
rect 37916 65248 37924 65312
rect 37604 64224 37924 65248
rect 37604 64160 37612 64224
rect 37676 64160 37692 64224
rect 37756 64160 37772 64224
rect 37836 64160 37852 64224
rect 37916 64160 37924 64224
rect 37604 63954 37924 64160
rect 37604 63718 37646 63954
rect 37882 63718 37924 63954
rect 37604 63136 37924 63718
rect 37604 63072 37612 63136
rect 37676 63072 37692 63136
rect 37756 63072 37772 63136
rect 37836 63072 37852 63136
rect 37916 63072 37924 63136
rect 37604 62048 37924 63072
rect 37604 61984 37612 62048
rect 37676 61984 37692 62048
rect 37756 61984 37772 62048
rect 37836 61984 37852 62048
rect 37916 61984 37924 62048
rect 37604 60960 37924 61984
rect 37604 60896 37612 60960
rect 37676 60896 37692 60960
rect 37756 60896 37772 60960
rect 37836 60896 37852 60960
rect 37916 60896 37924 60960
rect 37604 59872 37924 60896
rect 37604 59808 37612 59872
rect 37676 59808 37692 59872
rect 37756 59808 37772 59872
rect 37836 59808 37852 59872
rect 37916 59808 37924 59872
rect 37604 58954 37924 59808
rect 37604 58784 37646 58954
rect 37882 58784 37924 58954
rect 37604 58720 37612 58784
rect 37916 58720 37924 58784
rect 37604 58718 37646 58720
rect 37882 58718 37924 58720
rect 37604 57696 37924 58718
rect 37604 57632 37612 57696
rect 37676 57632 37692 57696
rect 37756 57632 37772 57696
rect 37836 57632 37852 57696
rect 37916 57632 37924 57696
rect 37604 56608 37924 57632
rect 37604 56544 37612 56608
rect 37676 56544 37692 56608
rect 37756 56544 37772 56608
rect 37836 56544 37852 56608
rect 37916 56544 37924 56608
rect 37604 55520 37924 56544
rect 37604 55456 37612 55520
rect 37676 55456 37692 55520
rect 37756 55456 37772 55520
rect 37836 55456 37852 55520
rect 37916 55456 37924 55520
rect 37604 54432 37924 55456
rect 37604 54368 37612 54432
rect 37676 54368 37692 54432
rect 37756 54368 37772 54432
rect 37836 54368 37852 54432
rect 37916 54368 37924 54432
rect 37604 53954 37924 54368
rect 37604 53718 37646 53954
rect 37882 53718 37924 53954
rect 37604 53344 37924 53718
rect 37604 53280 37612 53344
rect 37676 53280 37692 53344
rect 37756 53280 37772 53344
rect 37836 53280 37852 53344
rect 37916 53280 37924 53344
rect 37604 52256 37924 53280
rect 37604 52192 37612 52256
rect 37676 52192 37692 52256
rect 37756 52192 37772 52256
rect 37836 52192 37852 52256
rect 37916 52192 37924 52256
rect 37604 51168 37924 52192
rect 37604 51104 37612 51168
rect 37676 51104 37692 51168
rect 37756 51104 37772 51168
rect 37836 51104 37852 51168
rect 37916 51104 37924 51168
rect 37604 50080 37924 51104
rect 37604 50016 37612 50080
rect 37676 50016 37692 50080
rect 37756 50016 37772 50080
rect 37836 50016 37852 50080
rect 37916 50016 37924 50080
rect 37604 48992 37924 50016
rect 37604 48928 37612 48992
rect 37676 48954 37692 48992
rect 37756 48954 37772 48992
rect 37836 48954 37852 48992
rect 37916 48928 37924 48992
rect 37604 48718 37646 48928
rect 37882 48718 37924 48928
rect 37604 47904 37924 48718
rect 37604 47840 37612 47904
rect 37676 47840 37692 47904
rect 37756 47840 37772 47904
rect 37836 47840 37852 47904
rect 37916 47840 37924 47904
rect 37604 46816 37924 47840
rect 37604 46752 37612 46816
rect 37676 46752 37692 46816
rect 37756 46752 37772 46816
rect 37836 46752 37852 46816
rect 37916 46752 37924 46816
rect 37604 45728 37924 46752
rect 37604 45664 37612 45728
rect 37676 45664 37692 45728
rect 37756 45664 37772 45728
rect 37836 45664 37852 45728
rect 37916 45664 37924 45728
rect 37604 44640 37924 45664
rect 37604 44576 37612 44640
rect 37676 44576 37692 44640
rect 37756 44576 37772 44640
rect 37836 44576 37852 44640
rect 37916 44576 37924 44640
rect 37604 43954 37924 44576
rect 37604 43718 37646 43954
rect 37882 43718 37924 43954
rect 37604 43552 37924 43718
rect 37604 43488 37612 43552
rect 37676 43488 37692 43552
rect 37756 43488 37772 43552
rect 37836 43488 37852 43552
rect 37916 43488 37924 43552
rect 37604 42464 37924 43488
rect 37604 42400 37612 42464
rect 37676 42400 37692 42464
rect 37756 42400 37772 42464
rect 37836 42400 37852 42464
rect 37916 42400 37924 42464
rect 37604 41376 37924 42400
rect 37604 41312 37612 41376
rect 37676 41312 37692 41376
rect 37756 41312 37772 41376
rect 37836 41312 37852 41376
rect 37916 41312 37924 41376
rect 37604 40288 37924 41312
rect 37604 40224 37612 40288
rect 37676 40224 37692 40288
rect 37756 40224 37772 40288
rect 37836 40224 37852 40288
rect 37916 40224 37924 40288
rect 37604 39200 37924 40224
rect 37604 39136 37612 39200
rect 37676 39136 37692 39200
rect 37756 39136 37772 39200
rect 37836 39136 37852 39200
rect 37916 39136 37924 39200
rect 37604 38954 37924 39136
rect 37604 38718 37646 38954
rect 37882 38718 37924 38954
rect 37604 38112 37924 38718
rect 37604 38048 37612 38112
rect 37676 38048 37692 38112
rect 37756 38048 37772 38112
rect 37836 38048 37852 38112
rect 37916 38048 37924 38112
rect 37604 37024 37924 38048
rect 37604 36960 37612 37024
rect 37676 36960 37692 37024
rect 37756 36960 37772 37024
rect 37836 36960 37852 37024
rect 37916 36960 37924 37024
rect 37604 35936 37924 36960
rect 37604 35872 37612 35936
rect 37676 35872 37692 35936
rect 37756 35872 37772 35936
rect 37836 35872 37852 35936
rect 37916 35872 37924 35936
rect 37604 34848 37924 35872
rect 37604 34784 37612 34848
rect 37676 34784 37692 34848
rect 37756 34784 37772 34848
rect 37836 34784 37852 34848
rect 37916 34784 37924 34848
rect 37604 33954 37924 34784
rect 37604 33760 37646 33954
rect 37882 33760 37924 33954
rect 37604 33696 37612 33760
rect 37676 33696 37692 33718
rect 37756 33696 37772 33718
rect 37836 33696 37852 33718
rect 37916 33696 37924 33760
rect 37604 32672 37924 33696
rect 37604 32608 37612 32672
rect 37676 32608 37692 32672
rect 37756 32608 37772 32672
rect 37836 32608 37852 32672
rect 37916 32608 37924 32672
rect 37604 31584 37924 32608
rect 37604 31520 37612 31584
rect 37676 31520 37692 31584
rect 37756 31520 37772 31584
rect 37836 31520 37852 31584
rect 37916 31520 37924 31584
rect 37604 30496 37924 31520
rect 37604 30432 37612 30496
rect 37676 30432 37692 30496
rect 37756 30432 37772 30496
rect 37836 30432 37852 30496
rect 37916 30432 37924 30496
rect 37604 29408 37924 30432
rect 37604 29344 37612 29408
rect 37676 29344 37692 29408
rect 37756 29344 37772 29408
rect 37836 29344 37852 29408
rect 37916 29344 37924 29408
rect 37604 28954 37924 29344
rect 37604 28718 37646 28954
rect 37882 28718 37924 28954
rect 37604 28320 37924 28718
rect 37604 28256 37612 28320
rect 37676 28256 37692 28320
rect 37756 28256 37772 28320
rect 37836 28256 37852 28320
rect 37916 28256 37924 28320
rect 37604 27232 37924 28256
rect 37604 27168 37612 27232
rect 37676 27168 37692 27232
rect 37756 27168 37772 27232
rect 37836 27168 37852 27232
rect 37916 27168 37924 27232
rect 37604 26144 37924 27168
rect 37604 26080 37612 26144
rect 37676 26080 37692 26144
rect 37756 26080 37772 26144
rect 37836 26080 37852 26144
rect 37916 26080 37924 26144
rect 37604 25056 37924 26080
rect 37604 24992 37612 25056
rect 37676 24992 37692 25056
rect 37756 24992 37772 25056
rect 37836 24992 37852 25056
rect 37916 24992 37924 25056
rect 37604 23968 37924 24992
rect 37604 23904 37612 23968
rect 37676 23954 37692 23968
rect 37756 23954 37772 23968
rect 37836 23954 37852 23968
rect 37916 23904 37924 23968
rect 37604 23718 37646 23904
rect 37882 23718 37924 23904
rect 37604 22880 37924 23718
rect 37604 22816 37612 22880
rect 37676 22816 37692 22880
rect 37756 22816 37772 22880
rect 37836 22816 37852 22880
rect 37916 22816 37924 22880
rect 37604 21792 37924 22816
rect 37604 21728 37612 21792
rect 37676 21728 37692 21792
rect 37756 21728 37772 21792
rect 37836 21728 37852 21792
rect 37916 21728 37924 21792
rect 37604 20704 37924 21728
rect 37604 20640 37612 20704
rect 37676 20640 37692 20704
rect 37756 20640 37772 20704
rect 37836 20640 37852 20704
rect 37916 20640 37924 20704
rect 37604 19616 37924 20640
rect 37604 19552 37612 19616
rect 37676 19552 37692 19616
rect 37756 19552 37772 19616
rect 37836 19552 37852 19616
rect 37916 19552 37924 19616
rect 37604 18954 37924 19552
rect 37604 18718 37646 18954
rect 37882 18718 37924 18954
rect 37604 18528 37924 18718
rect 37604 18464 37612 18528
rect 37676 18464 37692 18528
rect 37756 18464 37772 18528
rect 37836 18464 37852 18528
rect 37916 18464 37924 18528
rect 37604 17440 37924 18464
rect 37604 17376 37612 17440
rect 37676 17376 37692 17440
rect 37756 17376 37772 17440
rect 37836 17376 37852 17440
rect 37916 17376 37924 17440
rect 37604 16352 37924 17376
rect 37604 16288 37612 16352
rect 37676 16288 37692 16352
rect 37756 16288 37772 16352
rect 37836 16288 37852 16352
rect 37916 16288 37924 16352
rect 37604 15264 37924 16288
rect 37604 15200 37612 15264
rect 37676 15200 37692 15264
rect 37756 15200 37772 15264
rect 37836 15200 37852 15264
rect 37916 15200 37924 15264
rect 37604 14176 37924 15200
rect 37604 14112 37612 14176
rect 37676 14112 37692 14176
rect 37756 14112 37772 14176
rect 37836 14112 37852 14176
rect 37916 14112 37924 14176
rect 37604 13954 37924 14112
rect 37604 13718 37646 13954
rect 37882 13718 37924 13954
rect 37604 13088 37924 13718
rect 37604 13024 37612 13088
rect 37676 13024 37692 13088
rect 37756 13024 37772 13088
rect 37836 13024 37852 13088
rect 37916 13024 37924 13088
rect 37604 12000 37924 13024
rect 37604 11936 37612 12000
rect 37676 11936 37692 12000
rect 37756 11936 37772 12000
rect 37836 11936 37852 12000
rect 37916 11936 37924 12000
rect 37604 10912 37924 11936
rect 37604 10848 37612 10912
rect 37676 10848 37692 10912
rect 37756 10848 37772 10912
rect 37836 10848 37852 10912
rect 37916 10848 37924 10912
rect 37604 9824 37924 10848
rect 37604 9760 37612 9824
rect 37676 9760 37692 9824
rect 37756 9760 37772 9824
rect 37836 9760 37852 9824
rect 37916 9760 37924 9824
rect 37604 8954 37924 9760
rect 37604 8736 37646 8954
rect 37882 8736 37924 8954
rect 37604 8672 37612 8736
rect 37676 8672 37692 8718
rect 37756 8672 37772 8718
rect 37836 8672 37852 8718
rect 37916 8672 37924 8736
rect 37604 7648 37924 8672
rect 37604 7584 37612 7648
rect 37676 7584 37692 7648
rect 37756 7584 37772 7648
rect 37836 7584 37852 7648
rect 37916 7584 37924 7648
rect 37604 6560 37924 7584
rect 37604 6496 37612 6560
rect 37676 6496 37692 6560
rect 37756 6496 37772 6560
rect 37836 6496 37852 6560
rect 37916 6496 37924 6560
rect 37604 5472 37924 6496
rect 37604 5408 37612 5472
rect 37676 5408 37692 5472
rect 37756 5408 37772 5472
rect 37836 5408 37852 5472
rect 37916 5408 37924 5472
rect 37604 4384 37924 5408
rect 37604 4320 37612 4384
rect 37676 4320 37692 4384
rect 37756 4320 37772 4384
rect 37836 4320 37852 4384
rect 37916 4320 37924 4384
rect 37604 3954 37924 4320
rect 37604 3718 37646 3954
rect 37882 3718 37924 3954
rect 37604 3296 37924 3718
rect 37604 3232 37612 3296
rect 37676 3232 37692 3296
rect 37756 3232 37772 3296
rect 37836 3232 37852 3296
rect 37916 3232 37924 3296
rect 37604 2208 37924 3232
rect 37604 2144 37612 2208
rect 37676 2144 37692 2208
rect 37756 2144 37772 2208
rect 37836 2144 37852 2208
rect 37916 2144 37924 2208
rect 37604 2128 37924 2144
<< via4 >>
rect 1986 68058 2222 68294
rect 1986 63058 2222 63294
rect 1986 58240 2222 58294
rect 1986 58176 2016 58240
rect 2016 58176 2032 58240
rect 2032 58176 2096 58240
rect 2096 58176 2112 58240
rect 2112 58176 2176 58240
rect 2176 58176 2192 58240
rect 2192 58176 2222 58240
rect 1986 58058 2222 58176
rect 1986 53058 2222 53294
rect 1986 48058 2222 48294
rect 1986 43058 2222 43294
rect 1986 38058 2222 38294
rect 1986 33216 2222 33294
rect 1986 33152 2016 33216
rect 2016 33152 2032 33216
rect 2032 33152 2096 33216
rect 2096 33152 2112 33216
rect 2112 33152 2176 33216
rect 2176 33152 2192 33216
rect 2192 33152 2222 33216
rect 1986 33058 2222 33152
rect 1986 28058 2222 28294
rect 1986 23058 2222 23294
rect 1986 18058 2222 18294
rect 1986 13058 2222 13294
rect 1986 8192 2222 8294
rect 1986 8128 2016 8192
rect 2016 8128 2032 8192
rect 2032 8128 2096 8192
rect 2096 8128 2112 8192
rect 2112 8128 2176 8192
rect 2176 8128 2192 8192
rect 2192 8128 2222 8192
rect 1986 8058 2222 8128
rect 1986 3058 2222 3294
rect 2646 68718 2882 68954
rect 2646 63718 2882 63954
rect 2646 58784 2882 58954
rect 2646 58720 2676 58784
rect 2676 58720 2692 58784
rect 2692 58720 2756 58784
rect 2756 58720 2772 58784
rect 2772 58720 2836 58784
rect 2836 58720 2852 58784
rect 2852 58720 2882 58784
rect 2646 58718 2882 58720
rect 2646 53718 2882 53954
rect 2646 48928 2676 48954
rect 2676 48928 2692 48954
rect 2692 48928 2756 48954
rect 2756 48928 2772 48954
rect 2772 48928 2836 48954
rect 2836 48928 2852 48954
rect 2852 48928 2882 48954
rect 2646 48718 2882 48928
rect 2646 43718 2882 43954
rect 2646 38718 2882 38954
rect 2646 33760 2882 33954
rect 2646 33718 2676 33760
rect 2676 33718 2692 33760
rect 2692 33718 2756 33760
rect 2756 33718 2772 33760
rect 2772 33718 2836 33760
rect 2836 33718 2852 33760
rect 2852 33718 2882 33760
rect 2646 28718 2882 28954
rect 2646 23904 2676 23954
rect 2676 23904 2692 23954
rect 2692 23904 2756 23954
rect 2756 23904 2772 23954
rect 2772 23904 2836 23954
rect 2836 23904 2852 23954
rect 2852 23904 2882 23954
rect 2646 23718 2882 23904
rect 2646 18718 2882 18954
rect 2646 13718 2882 13954
rect 2646 8736 2882 8954
rect 2646 8718 2676 8736
rect 2676 8718 2692 8736
rect 2692 8718 2756 8736
rect 2756 8718 2772 8736
rect 2772 8718 2836 8736
rect 2836 8718 2852 8736
rect 2852 8718 2882 8736
rect 2646 3718 2882 3954
rect 6986 68058 7222 68294
rect 6986 63058 7222 63294
rect 6986 58240 7222 58294
rect 6986 58176 7016 58240
rect 7016 58176 7032 58240
rect 7032 58176 7096 58240
rect 7096 58176 7112 58240
rect 7112 58176 7176 58240
rect 7176 58176 7192 58240
rect 7192 58176 7222 58240
rect 6986 58058 7222 58176
rect 6986 53058 7222 53294
rect 6986 48058 7222 48294
rect 6986 43058 7222 43294
rect 6986 38058 7222 38294
rect 6986 33216 7222 33294
rect 6986 33152 7016 33216
rect 7016 33152 7032 33216
rect 7032 33152 7096 33216
rect 7096 33152 7112 33216
rect 7112 33152 7176 33216
rect 7176 33152 7192 33216
rect 7192 33152 7222 33216
rect 6986 33058 7222 33152
rect 6986 28058 7222 28294
rect 6986 23058 7222 23294
rect 6986 18058 7222 18294
rect 6986 13058 7222 13294
rect 6986 8192 7222 8294
rect 6986 8128 7016 8192
rect 7016 8128 7032 8192
rect 7032 8128 7096 8192
rect 7096 8128 7112 8192
rect 7112 8128 7176 8192
rect 7176 8128 7192 8192
rect 7192 8128 7222 8192
rect 6986 8058 7222 8128
rect 6986 3058 7222 3294
rect 7646 68718 7882 68954
rect 7646 63718 7882 63954
rect 7646 58784 7882 58954
rect 7646 58720 7676 58784
rect 7676 58720 7692 58784
rect 7692 58720 7756 58784
rect 7756 58720 7772 58784
rect 7772 58720 7836 58784
rect 7836 58720 7852 58784
rect 7852 58720 7882 58784
rect 7646 58718 7882 58720
rect 7646 53718 7882 53954
rect 7646 48928 7676 48954
rect 7676 48928 7692 48954
rect 7692 48928 7756 48954
rect 7756 48928 7772 48954
rect 7772 48928 7836 48954
rect 7836 48928 7852 48954
rect 7852 48928 7882 48954
rect 7646 48718 7882 48928
rect 7646 43718 7882 43954
rect 7646 38718 7882 38954
rect 7646 33760 7882 33954
rect 7646 33718 7676 33760
rect 7676 33718 7692 33760
rect 7692 33718 7756 33760
rect 7756 33718 7772 33760
rect 7772 33718 7836 33760
rect 7836 33718 7852 33760
rect 7852 33718 7882 33760
rect 7646 28718 7882 28954
rect 7646 23904 7676 23954
rect 7676 23904 7692 23954
rect 7692 23904 7756 23954
rect 7756 23904 7772 23954
rect 7772 23904 7836 23954
rect 7836 23904 7852 23954
rect 7852 23904 7882 23954
rect 7646 23718 7882 23904
rect 7646 18718 7882 18954
rect 7646 13718 7882 13954
rect 7646 8736 7882 8954
rect 7646 8718 7676 8736
rect 7676 8718 7692 8736
rect 7692 8718 7756 8736
rect 7756 8718 7772 8736
rect 7772 8718 7836 8736
rect 7836 8718 7852 8736
rect 7852 8718 7882 8736
rect 7646 3718 7882 3954
rect 11986 68058 12222 68294
rect 11986 63058 12222 63294
rect 11986 58240 12222 58294
rect 11986 58176 12016 58240
rect 12016 58176 12032 58240
rect 12032 58176 12096 58240
rect 12096 58176 12112 58240
rect 12112 58176 12176 58240
rect 12176 58176 12192 58240
rect 12192 58176 12222 58240
rect 11986 58058 12222 58176
rect 11986 53058 12222 53294
rect 11986 48058 12222 48294
rect 11986 43058 12222 43294
rect 11986 38058 12222 38294
rect 11986 33216 12222 33294
rect 11986 33152 12016 33216
rect 12016 33152 12032 33216
rect 12032 33152 12096 33216
rect 12096 33152 12112 33216
rect 12112 33152 12176 33216
rect 12176 33152 12192 33216
rect 12192 33152 12222 33216
rect 11986 33058 12222 33152
rect 11986 28058 12222 28294
rect 11986 23058 12222 23294
rect 11986 18058 12222 18294
rect 11986 13058 12222 13294
rect 11986 8192 12222 8294
rect 11986 8128 12016 8192
rect 12016 8128 12032 8192
rect 12032 8128 12096 8192
rect 12096 8128 12112 8192
rect 12112 8128 12176 8192
rect 12176 8128 12192 8192
rect 12192 8128 12222 8192
rect 11986 8058 12222 8128
rect 11986 3058 12222 3294
rect 12646 68718 12882 68954
rect 12646 63718 12882 63954
rect 12646 58784 12882 58954
rect 12646 58720 12676 58784
rect 12676 58720 12692 58784
rect 12692 58720 12756 58784
rect 12756 58720 12772 58784
rect 12772 58720 12836 58784
rect 12836 58720 12852 58784
rect 12852 58720 12882 58784
rect 12646 58718 12882 58720
rect 12646 53718 12882 53954
rect 12646 48928 12676 48954
rect 12676 48928 12692 48954
rect 12692 48928 12756 48954
rect 12756 48928 12772 48954
rect 12772 48928 12836 48954
rect 12836 48928 12852 48954
rect 12852 48928 12882 48954
rect 12646 48718 12882 48928
rect 12646 43718 12882 43954
rect 12646 38718 12882 38954
rect 12646 33760 12882 33954
rect 12646 33718 12676 33760
rect 12676 33718 12692 33760
rect 12692 33718 12756 33760
rect 12756 33718 12772 33760
rect 12772 33718 12836 33760
rect 12836 33718 12852 33760
rect 12852 33718 12882 33760
rect 12646 28718 12882 28954
rect 12646 23904 12676 23954
rect 12676 23904 12692 23954
rect 12692 23904 12756 23954
rect 12756 23904 12772 23954
rect 12772 23904 12836 23954
rect 12836 23904 12852 23954
rect 12852 23904 12882 23954
rect 12646 23718 12882 23904
rect 12646 18718 12882 18954
rect 12646 13718 12882 13954
rect 12646 8736 12882 8954
rect 12646 8718 12676 8736
rect 12676 8718 12692 8736
rect 12692 8718 12756 8736
rect 12756 8718 12772 8736
rect 12772 8718 12836 8736
rect 12836 8718 12852 8736
rect 12852 8718 12882 8736
rect 12646 3718 12882 3954
rect 16986 68058 17222 68294
rect 16986 63058 17222 63294
rect 16986 58240 17222 58294
rect 16986 58176 17016 58240
rect 17016 58176 17032 58240
rect 17032 58176 17096 58240
rect 17096 58176 17112 58240
rect 17112 58176 17176 58240
rect 17176 58176 17192 58240
rect 17192 58176 17222 58240
rect 16986 58058 17222 58176
rect 16986 53058 17222 53294
rect 16986 48058 17222 48294
rect 16986 43058 17222 43294
rect 16986 38058 17222 38294
rect 16986 33216 17222 33294
rect 16986 33152 17016 33216
rect 17016 33152 17032 33216
rect 17032 33152 17096 33216
rect 17096 33152 17112 33216
rect 17112 33152 17176 33216
rect 17176 33152 17192 33216
rect 17192 33152 17222 33216
rect 16986 33058 17222 33152
rect 16986 28058 17222 28294
rect 16986 23058 17222 23294
rect 16986 18058 17222 18294
rect 16986 13058 17222 13294
rect 16986 8192 17222 8294
rect 16986 8128 17016 8192
rect 17016 8128 17032 8192
rect 17032 8128 17096 8192
rect 17096 8128 17112 8192
rect 17112 8128 17176 8192
rect 17176 8128 17192 8192
rect 17192 8128 17222 8192
rect 16986 8058 17222 8128
rect 16986 3058 17222 3294
rect 17646 68718 17882 68954
rect 17646 63718 17882 63954
rect 17646 58784 17882 58954
rect 17646 58720 17676 58784
rect 17676 58720 17692 58784
rect 17692 58720 17756 58784
rect 17756 58720 17772 58784
rect 17772 58720 17836 58784
rect 17836 58720 17852 58784
rect 17852 58720 17882 58784
rect 17646 58718 17882 58720
rect 17646 53718 17882 53954
rect 17646 48928 17676 48954
rect 17676 48928 17692 48954
rect 17692 48928 17756 48954
rect 17756 48928 17772 48954
rect 17772 48928 17836 48954
rect 17836 48928 17852 48954
rect 17852 48928 17882 48954
rect 17646 48718 17882 48928
rect 21986 68058 22222 68294
rect 21986 63058 22222 63294
rect 21986 58240 22222 58294
rect 21986 58176 22016 58240
rect 22016 58176 22032 58240
rect 22032 58176 22096 58240
rect 22096 58176 22112 58240
rect 22112 58176 22176 58240
rect 22176 58176 22192 58240
rect 22192 58176 22222 58240
rect 21986 58058 22222 58176
rect 21986 53058 22222 53294
rect 21986 48058 22222 48294
rect 17646 43718 17882 43954
rect 17646 38718 17882 38954
rect 17646 33760 17882 33954
rect 21986 43058 22222 43294
rect 21986 38058 22222 38294
rect 17646 33718 17676 33760
rect 17676 33718 17692 33760
rect 17692 33718 17756 33760
rect 17756 33718 17772 33760
rect 17772 33718 17836 33760
rect 17836 33718 17852 33760
rect 17852 33718 17882 33760
rect 17646 28718 17882 28954
rect 17646 23904 17676 23954
rect 17676 23904 17692 23954
rect 17692 23904 17756 23954
rect 17756 23904 17772 23954
rect 17772 23904 17836 23954
rect 17836 23904 17852 23954
rect 17852 23904 17882 23954
rect 17646 23718 17882 23904
rect 21986 33216 22222 33294
rect 21986 33152 22016 33216
rect 22016 33152 22032 33216
rect 22032 33152 22096 33216
rect 22096 33152 22112 33216
rect 22112 33152 22176 33216
rect 22176 33152 22192 33216
rect 22192 33152 22222 33216
rect 21986 33058 22222 33152
rect 21986 28058 22222 28294
rect 21986 23058 22222 23294
rect 17646 18718 17882 18954
rect 17646 13718 17882 13954
rect 17646 8736 17882 8954
rect 17646 8718 17676 8736
rect 17676 8718 17692 8736
rect 17692 8718 17756 8736
rect 17756 8718 17772 8736
rect 17772 8718 17836 8736
rect 17836 8718 17852 8736
rect 17852 8718 17882 8736
rect 17646 3718 17882 3954
rect 21986 18058 22222 18294
rect 21986 13058 22222 13294
rect 21986 8192 22222 8294
rect 21986 8128 22016 8192
rect 22016 8128 22032 8192
rect 22032 8128 22096 8192
rect 22096 8128 22112 8192
rect 22112 8128 22176 8192
rect 22176 8128 22192 8192
rect 22192 8128 22222 8192
rect 21986 8058 22222 8128
rect 21986 3058 22222 3294
rect 22646 68718 22882 68954
rect 22646 63718 22882 63954
rect 22646 58784 22882 58954
rect 22646 58720 22676 58784
rect 22676 58720 22692 58784
rect 22692 58720 22756 58784
rect 22756 58720 22772 58784
rect 22772 58720 22836 58784
rect 22836 58720 22852 58784
rect 22852 58720 22882 58784
rect 22646 58718 22882 58720
rect 22646 53718 22882 53954
rect 22646 48928 22676 48954
rect 22676 48928 22692 48954
rect 22692 48928 22756 48954
rect 22756 48928 22772 48954
rect 22772 48928 22836 48954
rect 22836 48928 22852 48954
rect 22852 48928 22882 48954
rect 22646 48718 22882 48928
rect 22646 43718 22882 43954
rect 22646 38718 22882 38954
rect 22646 33760 22882 33954
rect 22646 33718 22676 33760
rect 22676 33718 22692 33760
rect 22692 33718 22756 33760
rect 22756 33718 22772 33760
rect 22772 33718 22836 33760
rect 22836 33718 22852 33760
rect 22852 33718 22882 33760
rect 22646 28718 22882 28954
rect 22646 23904 22676 23954
rect 22676 23904 22692 23954
rect 22692 23904 22756 23954
rect 22756 23904 22772 23954
rect 22772 23904 22836 23954
rect 22836 23904 22852 23954
rect 22852 23904 22882 23954
rect 22646 23718 22882 23904
rect 22646 18718 22882 18954
rect 22646 13718 22882 13954
rect 22646 8736 22882 8954
rect 22646 8718 22676 8736
rect 22676 8718 22692 8736
rect 22692 8718 22756 8736
rect 22756 8718 22772 8736
rect 22772 8718 22836 8736
rect 22836 8718 22852 8736
rect 22852 8718 22882 8736
rect 22646 3718 22882 3954
rect 26986 68058 27222 68294
rect 26986 63058 27222 63294
rect 26986 58240 27222 58294
rect 26986 58176 27016 58240
rect 27016 58176 27032 58240
rect 27032 58176 27096 58240
rect 27096 58176 27112 58240
rect 27112 58176 27176 58240
rect 27176 58176 27192 58240
rect 27192 58176 27222 58240
rect 26986 58058 27222 58176
rect 26986 53058 27222 53294
rect 26986 48058 27222 48294
rect 26986 43058 27222 43294
rect 26986 38058 27222 38294
rect 26986 33216 27222 33294
rect 26986 33152 27016 33216
rect 27016 33152 27032 33216
rect 27032 33152 27096 33216
rect 27096 33152 27112 33216
rect 27112 33152 27176 33216
rect 27176 33152 27192 33216
rect 27192 33152 27222 33216
rect 26986 33058 27222 33152
rect 26986 28058 27222 28294
rect 26986 23058 27222 23294
rect 26986 18058 27222 18294
rect 26986 13058 27222 13294
rect 26986 8192 27222 8294
rect 26986 8128 27016 8192
rect 27016 8128 27032 8192
rect 27032 8128 27096 8192
rect 27096 8128 27112 8192
rect 27112 8128 27176 8192
rect 27176 8128 27192 8192
rect 27192 8128 27222 8192
rect 26986 8058 27222 8128
rect 26986 3058 27222 3294
rect 27646 68718 27882 68954
rect 31986 68058 32222 68294
rect 27646 63718 27882 63954
rect 27646 58784 27882 58954
rect 27646 58720 27676 58784
rect 27676 58720 27692 58784
rect 27692 58720 27756 58784
rect 27756 58720 27772 58784
rect 27772 58720 27836 58784
rect 27836 58720 27852 58784
rect 27852 58720 27882 58784
rect 27646 58718 27882 58720
rect 27646 53718 27882 53954
rect 31986 63058 32222 63294
rect 31986 58240 32222 58294
rect 31986 58176 32016 58240
rect 32016 58176 32032 58240
rect 32032 58176 32096 58240
rect 32096 58176 32112 58240
rect 32112 58176 32176 58240
rect 32176 58176 32192 58240
rect 32192 58176 32222 58240
rect 31986 58058 32222 58176
rect 31986 53058 32222 53294
rect 27646 48928 27676 48954
rect 27676 48928 27692 48954
rect 27692 48928 27756 48954
rect 27756 48928 27772 48954
rect 27772 48928 27836 48954
rect 27836 48928 27852 48954
rect 27852 48928 27882 48954
rect 27646 48718 27882 48928
rect 27646 43718 27882 43954
rect 32646 68718 32882 68954
rect 32646 63718 32882 63954
rect 32646 58784 32882 58954
rect 32646 58720 32676 58784
rect 32676 58720 32692 58784
rect 32692 58720 32756 58784
rect 32756 58720 32772 58784
rect 32772 58720 32836 58784
rect 32836 58720 32852 58784
rect 32852 58720 32882 58784
rect 32646 58718 32882 58720
rect 36986 68058 37222 68294
rect 36986 63058 37222 63294
rect 32646 53718 32882 53954
rect 31986 48058 32222 48294
rect 31986 43058 32222 43294
rect 27646 38718 27882 38954
rect 27646 33760 27882 33954
rect 27646 33718 27676 33760
rect 27676 33718 27692 33760
rect 27692 33718 27756 33760
rect 27756 33718 27772 33760
rect 27772 33718 27836 33760
rect 27836 33718 27852 33760
rect 27852 33718 27882 33760
rect 32646 48928 32676 48954
rect 32676 48928 32692 48954
rect 32692 48928 32756 48954
rect 32756 48928 32772 48954
rect 32772 48928 32836 48954
rect 32836 48928 32852 48954
rect 32852 48928 32882 48954
rect 32646 48718 32882 48928
rect 32646 43718 32882 43954
rect 31986 38058 32222 38294
rect 31986 33216 32222 33294
rect 31986 33152 32016 33216
rect 32016 33152 32032 33216
rect 32032 33152 32096 33216
rect 32096 33152 32112 33216
rect 32112 33152 32176 33216
rect 32176 33152 32192 33216
rect 32192 33152 32222 33216
rect 31986 33058 32222 33152
rect 27646 28718 27882 28954
rect 27646 23904 27676 23954
rect 27676 23904 27692 23954
rect 27692 23904 27756 23954
rect 27756 23904 27772 23954
rect 27772 23904 27836 23954
rect 27836 23904 27852 23954
rect 27852 23904 27882 23954
rect 27646 23718 27882 23904
rect 27646 18718 27882 18954
rect 27646 13718 27882 13954
rect 27646 8736 27882 8954
rect 27646 8718 27676 8736
rect 27676 8718 27692 8736
rect 27692 8718 27756 8736
rect 27756 8718 27772 8736
rect 27772 8718 27836 8736
rect 27836 8718 27852 8736
rect 27852 8718 27882 8736
rect 27646 3718 27882 3954
rect 31986 28058 32222 28294
rect 31986 23058 32222 23294
rect 31986 18058 32222 18294
rect 31986 13058 32222 13294
rect 31986 8192 32222 8294
rect 31986 8128 32016 8192
rect 32016 8128 32032 8192
rect 32032 8128 32096 8192
rect 32096 8128 32112 8192
rect 32112 8128 32176 8192
rect 32176 8128 32192 8192
rect 32192 8128 32222 8192
rect 31986 8058 32222 8128
rect 31986 3058 32222 3294
rect 32646 38718 32882 38954
rect 32646 33760 32882 33954
rect 32646 33718 32676 33760
rect 32676 33718 32692 33760
rect 32692 33718 32756 33760
rect 32756 33718 32772 33760
rect 32772 33718 32836 33760
rect 32836 33718 32852 33760
rect 32852 33718 32882 33760
rect 32646 28718 32882 28954
rect 32646 23904 32676 23954
rect 32676 23904 32692 23954
rect 32692 23904 32756 23954
rect 32756 23904 32772 23954
rect 32772 23904 32836 23954
rect 32836 23904 32852 23954
rect 32852 23904 32882 23954
rect 32646 23718 32882 23904
rect 32646 18718 32882 18954
rect 32646 13718 32882 13954
rect 36986 58240 37222 58294
rect 36986 58176 37016 58240
rect 37016 58176 37032 58240
rect 37032 58176 37096 58240
rect 37096 58176 37112 58240
rect 37112 58176 37176 58240
rect 37176 58176 37192 58240
rect 37192 58176 37222 58240
rect 36986 58058 37222 58176
rect 32646 8736 32882 8954
rect 32646 8718 32676 8736
rect 32676 8718 32692 8736
rect 32692 8718 32756 8736
rect 32756 8718 32772 8736
rect 32772 8718 32836 8736
rect 32836 8718 32852 8736
rect 32852 8718 32882 8736
rect 36986 53058 37222 53294
rect 36986 48058 37222 48294
rect 36986 43058 37222 43294
rect 36986 38058 37222 38294
rect 36986 33216 37222 33294
rect 36986 33152 37016 33216
rect 37016 33152 37032 33216
rect 37032 33152 37096 33216
rect 37096 33152 37112 33216
rect 37112 33152 37176 33216
rect 37176 33152 37192 33216
rect 37192 33152 37222 33216
rect 36986 33058 37222 33152
rect 36986 28058 37222 28294
rect 36986 23058 37222 23294
rect 36986 18058 37222 18294
rect 36986 13058 37222 13294
rect 36986 8192 37222 8294
rect 36986 8128 37016 8192
rect 37016 8128 37032 8192
rect 37032 8128 37096 8192
rect 37096 8128 37112 8192
rect 37112 8128 37176 8192
rect 37176 8128 37192 8192
rect 37192 8128 37222 8192
rect 36986 8058 37222 8128
rect 32646 3718 32882 3954
rect 36986 3058 37222 3294
rect 37646 68718 37882 68954
rect 37646 63718 37882 63954
rect 37646 58784 37882 58954
rect 37646 58720 37676 58784
rect 37676 58720 37692 58784
rect 37692 58720 37756 58784
rect 37756 58720 37772 58784
rect 37772 58720 37836 58784
rect 37836 58720 37852 58784
rect 37852 58720 37882 58784
rect 37646 58718 37882 58720
rect 37646 53718 37882 53954
rect 37646 48928 37676 48954
rect 37676 48928 37692 48954
rect 37692 48928 37756 48954
rect 37756 48928 37772 48954
rect 37772 48928 37836 48954
rect 37836 48928 37852 48954
rect 37852 48928 37882 48954
rect 37646 48718 37882 48928
rect 37646 43718 37882 43954
rect 37646 38718 37882 38954
rect 37646 33760 37882 33954
rect 37646 33718 37676 33760
rect 37676 33718 37692 33760
rect 37692 33718 37756 33760
rect 37756 33718 37772 33760
rect 37772 33718 37836 33760
rect 37836 33718 37852 33760
rect 37852 33718 37882 33760
rect 37646 28718 37882 28954
rect 37646 23904 37676 23954
rect 37676 23904 37692 23954
rect 37692 23904 37756 23954
rect 37756 23904 37772 23954
rect 37772 23904 37836 23954
rect 37836 23904 37852 23954
rect 37852 23904 37882 23954
rect 37646 23718 37882 23904
rect 37646 18718 37882 18954
rect 37646 13718 37882 13954
rect 37646 8736 37882 8954
rect 37646 8718 37676 8736
rect 37676 8718 37692 8736
rect 37692 8718 37756 8736
rect 37756 8718 37772 8736
rect 37772 8718 37836 8736
rect 37836 8718 37852 8736
rect 37852 8718 37882 8736
rect 37646 3718 37882 3954
<< metal5 >>
rect 1056 68954 40896 68996
rect 1056 68718 2646 68954
rect 2882 68718 7646 68954
rect 7882 68718 12646 68954
rect 12882 68718 17646 68954
rect 17882 68718 22646 68954
rect 22882 68718 27646 68954
rect 27882 68718 32646 68954
rect 32882 68718 37646 68954
rect 37882 68718 40896 68954
rect 1056 68676 40896 68718
rect 1056 68294 40896 68336
rect 1056 68058 1986 68294
rect 2222 68058 6986 68294
rect 7222 68058 11986 68294
rect 12222 68058 16986 68294
rect 17222 68058 21986 68294
rect 22222 68058 26986 68294
rect 27222 68058 31986 68294
rect 32222 68058 36986 68294
rect 37222 68058 40896 68294
rect 1056 68016 40896 68058
rect 1056 63954 40896 63996
rect 1056 63718 2646 63954
rect 2882 63718 7646 63954
rect 7882 63718 12646 63954
rect 12882 63718 17646 63954
rect 17882 63718 22646 63954
rect 22882 63718 27646 63954
rect 27882 63718 32646 63954
rect 32882 63718 37646 63954
rect 37882 63718 40896 63954
rect 1056 63676 40896 63718
rect 1056 63294 40896 63336
rect 1056 63058 1986 63294
rect 2222 63058 6986 63294
rect 7222 63058 11986 63294
rect 12222 63058 16986 63294
rect 17222 63058 21986 63294
rect 22222 63058 26986 63294
rect 27222 63058 31986 63294
rect 32222 63058 36986 63294
rect 37222 63058 40896 63294
rect 1056 63016 40896 63058
rect 1056 58954 40896 58996
rect 1056 58718 2646 58954
rect 2882 58718 7646 58954
rect 7882 58718 12646 58954
rect 12882 58718 17646 58954
rect 17882 58718 22646 58954
rect 22882 58718 27646 58954
rect 27882 58718 32646 58954
rect 32882 58718 37646 58954
rect 37882 58718 40896 58954
rect 1056 58676 40896 58718
rect 1056 58294 40896 58336
rect 1056 58058 1986 58294
rect 2222 58058 6986 58294
rect 7222 58058 11986 58294
rect 12222 58058 16986 58294
rect 17222 58058 21986 58294
rect 22222 58058 26986 58294
rect 27222 58058 31986 58294
rect 32222 58058 36986 58294
rect 37222 58058 40896 58294
rect 1056 58016 40896 58058
rect 1056 53954 40896 53996
rect 1056 53718 2646 53954
rect 2882 53718 7646 53954
rect 7882 53718 12646 53954
rect 12882 53718 17646 53954
rect 17882 53718 22646 53954
rect 22882 53718 27646 53954
rect 27882 53718 32646 53954
rect 32882 53718 37646 53954
rect 37882 53718 40896 53954
rect 1056 53676 40896 53718
rect 1056 53294 40896 53336
rect 1056 53058 1986 53294
rect 2222 53058 6986 53294
rect 7222 53058 11986 53294
rect 12222 53058 16986 53294
rect 17222 53058 21986 53294
rect 22222 53058 26986 53294
rect 27222 53058 31986 53294
rect 32222 53058 36986 53294
rect 37222 53058 40896 53294
rect 1056 53016 40896 53058
rect 1056 48954 40896 48996
rect 1056 48718 2646 48954
rect 2882 48718 7646 48954
rect 7882 48718 12646 48954
rect 12882 48718 17646 48954
rect 17882 48718 22646 48954
rect 22882 48718 27646 48954
rect 27882 48718 32646 48954
rect 32882 48718 37646 48954
rect 37882 48718 40896 48954
rect 1056 48676 40896 48718
rect 1056 48294 40896 48336
rect 1056 48058 1986 48294
rect 2222 48058 6986 48294
rect 7222 48058 11986 48294
rect 12222 48058 16986 48294
rect 17222 48058 21986 48294
rect 22222 48058 26986 48294
rect 27222 48058 31986 48294
rect 32222 48058 36986 48294
rect 37222 48058 40896 48294
rect 1056 48016 40896 48058
rect 1056 43954 40896 43996
rect 1056 43718 2646 43954
rect 2882 43718 7646 43954
rect 7882 43718 12646 43954
rect 12882 43718 17646 43954
rect 17882 43718 22646 43954
rect 22882 43718 27646 43954
rect 27882 43718 32646 43954
rect 32882 43718 37646 43954
rect 37882 43718 40896 43954
rect 1056 43676 40896 43718
rect 1056 43294 40896 43336
rect 1056 43058 1986 43294
rect 2222 43058 6986 43294
rect 7222 43058 11986 43294
rect 12222 43058 16986 43294
rect 17222 43058 21986 43294
rect 22222 43058 26986 43294
rect 27222 43058 31986 43294
rect 32222 43058 36986 43294
rect 37222 43058 40896 43294
rect 1056 43016 40896 43058
rect 1056 38954 40896 38996
rect 1056 38718 2646 38954
rect 2882 38718 7646 38954
rect 7882 38718 12646 38954
rect 12882 38718 17646 38954
rect 17882 38718 22646 38954
rect 22882 38718 27646 38954
rect 27882 38718 32646 38954
rect 32882 38718 37646 38954
rect 37882 38718 40896 38954
rect 1056 38676 40896 38718
rect 1056 38294 40896 38336
rect 1056 38058 1986 38294
rect 2222 38058 6986 38294
rect 7222 38058 11986 38294
rect 12222 38058 16986 38294
rect 17222 38058 21986 38294
rect 22222 38058 26986 38294
rect 27222 38058 31986 38294
rect 32222 38058 36986 38294
rect 37222 38058 40896 38294
rect 1056 38016 40896 38058
rect 1056 33954 40896 33996
rect 1056 33718 2646 33954
rect 2882 33718 7646 33954
rect 7882 33718 12646 33954
rect 12882 33718 17646 33954
rect 17882 33718 22646 33954
rect 22882 33718 27646 33954
rect 27882 33718 32646 33954
rect 32882 33718 37646 33954
rect 37882 33718 40896 33954
rect 1056 33676 40896 33718
rect 1056 33294 40896 33336
rect 1056 33058 1986 33294
rect 2222 33058 6986 33294
rect 7222 33058 11986 33294
rect 12222 33058 16986 33294
rect 17222 33058 21986 33294
rect 22222 33058 26986 33294
rect 27222 33058 31986 33294
rect 32222 33058 36986 33294
rect 37222 33058 40896 33294
rect 1056 33016 40896 33058
rect 1056 28954 40896 28996
rect 1056 28718 2646 28954
rect 2882 28718 7646 28954
rect 7882 28718 12646 28954
rect 12882 28718 17646 28954
rect 17882 28718 22646 28954
rect 22882 28718 27646 28954
rect 27882 28718 32646 28954
rect 32882 28718 37646 28954
rect 37882 28718 40896 28954
rect 1056 28676 40896 28718
rect 1056 28294 40896 28336
rect 1056 28058 1986 28294
rect 2222 28058 6986 28294
rect 7222 28058 11986 28294
rect 12222 28058 16986 28294
rect 17222 28058 21986 28294
rect 22222 28058 26986 28294
rect 27222 28058 31986 28294
rect 32222 28058 36986 28294
rect 37222 28058 40896 28294
rect 1056 28016 40896 28058
rect 1056 23954 40896 23996
rect 1056 23718 2646 23954
rect 2882 23718 7646 23954
rect 7882 23718 12646 23954
rect 12882 23718 17646 23954
rect 17882 23718 22646 23954
rect 22882 23718 27646 23954
rect 27882 23718 32646 23954
rect 32882 23718 37646 23954
rect 37882 23718 40896 23954
rect 1056 23676 40896 23718
rect 1056 23294 40896 23336
rect 1056 23058 1986 23294
rect 2222 23058 6986 23294
rect 7222 23058 11986 23294
rect 12222 23058 16986 23294
rect 17222 23058 21986 23294
rect 22222 23058 26986 23294
rect 27222 23058 31986 23294
rect 32222 23058 36986 23294
rect 37222 23058 40896 23294
rect 1056 23016 40896 23058
rect 1056 18954 40896 18996
rect 1056 18718 2646 18954
rect 2882 18718 7646 18954
rect 7882 18718 12646 18954
rect 12882 18718 17646 18954
rect 17882 18718 22646 18954
rect 22882 18718 27646 18954
rect 27882 18718 32646 18954
rect 32882 18718 37646 18954
rect 37882 18718 40896 18954
rect 1056 18676 40896 18718
rect 1056 18294 40896 18336
rect 1056 18058 1986 18294
rect 2222 18058 6986 18294
rect 7222 18058 11986 18294
rect 12222 18058 16986 18294
rect 17222 18058 21986 18294
rect 22222 18058 26986 18294
rect 27222 18058 31986 18294
rect 32222 18058 36986 18294
rect 37222 18058 40896 18294
rect 1056 18016 40896 18058
rect 1056 13954 40896 13996
rect 1056 13718 2646 13954
rect 2882 13718 7646 13954
rect 7882 13718 12646 13954
rect 12882 13718 17646 13954
rect 17882 13718 22646 13954
rect 22882 13718 27646 13954
rect 27882 13718 32646 13954
rect 32882 13718 37646 13954
rect 37882 13718 40896 13954
rect 1056 13676 40896 13718
rect 1056 13294 40896 13336
rect 1056 13058 1986 13294
rect 2222 13058 6986 13294
rect 7222 13058 11986 13294
rect 12222 13058 16986 13294
rect 17222 13058 21986 13294
rect 22222 13058 26986 13294
rect 27222 13058 31986 13294
rect 32222 13058 36986 13294
rect 37222 13058 40896 13294
rect 1056 13016 40896 13058
rect 1056 8954 40896 8996
rect 1056 8718 2646 8954
rect 2882 8718 7646 8954
rect 7882 8718 12646 8954
rect 12882 8718 17646 8954
rect 17882 8718 22646 8954
rect 22882 8718 27646 8954
rect 27882 8718 32646 8954
rect 32882 8718 37646 8954
rect 37882 8718 40896 8954
rect 1056 8676 40896 8718
rect 1056 8294 40896 8336
rect 1056 8058 1986 8294
rect 2222 8058 6986 8294
rect 7222 8058 11986 8294
rect 12222 8058 16986 8294
rect 17222 8058 21986 8294
rect 22222 8058 26986 8294
rect 27222 8058 31986 8294
rect 32222 8058 36986 8294
rect 37222 8058 40896 8294
rect 1056 8016 40896 8058
rect 1056 3954 40896 3996
rect 1056 3718 2646 3954
rect 2882 3718 7646 3954
rect 7882 3718 12646 3954
rect 12882 3718 17646 3954
rect 17882 3718 22646 3954
rect 22882 3718 27646 3954
rect 27882 3718 32646 3954
rect 32882 3718 37646 3954
rect 37882 3718 40896 3954
rect 1056 3676 40896 3718
rect 1056 3294 40896 3336
rect 1056 3058 1986 3294
rect 2222 3058 6986 3294
rect 7222 3058 11986 3294
rect 12222 3058 16986 3294
rect 17222 3058 21986 3294
rect 22222 3058 26986 3294
rect 27222 3058 31986 3294
rect 32222 3058 36986 3294
rect 37222 3058 40896 3294
rect 1056 3016 40896 3058
use sky130_fd_sc_hd__and3_4  _162_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 22632 0 -1 65280
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _163_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 39928 0 -1 58752
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_4  _164_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 34132 0 -1 10880
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_2  _165_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 36984 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_4  _166_
timestamp 1704896540
transform -1 0 25852 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _167_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2116 0 1 47872
box -38 -48 866 592
use sky130_fd_sc_hd__o2bb2a_2  _168_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 34684 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _169_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 20608 0 1 63104
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _170_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2116 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_2  _171_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 17940 0 -1 54400
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _172_
timestamp 1704896540
transform -1 0 33028 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _173_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 39836 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _174_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 39744 0 1 54400
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _175_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 25116 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _176_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 22356 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__and4_4  _177_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 24380 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__and4_2  _178_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 5704 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__and2_4  _179_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 18124 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and4_2  _180_
timestamp 1704896540
transform 1 0 16468 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _181_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 37536 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_2  _182_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 35972 0 1 68544
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_1  _183_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 32844 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_2  _184_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 31188 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__and4_4  _185_
timestamp 1704896540
transform -1 0 3680 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__o211ai_4  _186_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6624 0 -1 41344
box -38 -48 1602 592
use sky130_fd_sc_hd__a21bo_4  _187_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 15272 0 -1 67456
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _188_
timestamp 1704896540
transform -1 0 7268 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _189_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_2  _190_
timestamp 1704896540
transform -1 0 29440 0 -1 50048
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _191_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 37996 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _192_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 37628 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _193_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 33396 0 1 48960
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _194_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 33120 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_2  _195_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9476 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _196_
timestamp 1704896540
transform -1 0 14628 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _197_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 33672 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _198_
timestamp 1704896540
transform 1 0 2024 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _199_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 11224 0 -1 65280
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _200_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 26312 0 1 64192
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _201_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 33028 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_8  _202_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 7360 0 -1 29376
box -38 -48 1050 592
use sky130_fd_sc_hd__nand2_2  _203_
timestamp 1704896540
transform 1 0 23552 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _204_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 24840 0 1 67456
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _205_
timestamp 1704896540
transform -1 0 38180 0 1 59840
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _206_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 13892 0 1 53312
box -38 -48 958 592
use sky130_fd_sc_hd__a21oi_1  _207_
timestamp 1704896540
transform 1 0 13984 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__and3_4  _208_
timestamp 1704896540
transform -1 0 26128 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__nor3_1  _209_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 13156 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _210_
timestamp 1704896540
transform -1 0 28980 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_4  _211_
timestamp 1704896540
transform -1 0 36984 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__and3_2  _212_
timestamp 1704896540
transform -1 0 4784 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _213_
timestamp 1704896540
transform -1 0 15548 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _214_
timestamp 1704896540
transform -1 0 6348 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_4  _215_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1656 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__or2_2  _216_
timestamp 1704896540
transform 1 0 38548 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _217_
timestamp 1704896540
transform 1 0 17020 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _218_
timestamp 1704896540
transform -1 0 33948 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _219_
timestamp 1704896540
transform -1 0 18952 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _220_
timestamp 1704896540
transform -1 0 11960 0 1 64192
box -38 -48 1234 592
use sky130_fd_sc_hd__and4_4  _221_
timestamp 1704896540
transform 1 0 18492 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__nor3_2  _222_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 19964 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _223_
timestamp 1704896540
transform 1 0 11684 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _224_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 21804 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and3_2  _225_
timestamp 1704896540
transform 1 0 28796 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _226_
timestamp 1704896540
transform 1 0 30636 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__a21oi_2  _227_
timestamp 1704896540
transform -1 0 19872 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and3_4  _228_
timestamp 1704896540
transform -1 0 11592 0 1 51136
box -38 -48 866 592
use sky130_fd_sc_hd__nor3_2  _229_
timestamp 1704896540
transform -1 0 3588 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _230_
timestamp 1704896540
transform 1 0 29164 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _231_
timestamp 1704896540
transform 1 0 31372 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and3_2  _232_
timestamp 1704896540
transform -1 0 34224 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _233_
timestamp 1704896540
transform 1 0 5704 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_2  _234_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 28520 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_4  _235_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2392 0 1 40256
box -38 -48 1326 592
use sky130_fd_sc_hd__and3_2  _236_
timestamp 1704896540
transform 1 0 8924 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _237_
timestamp 1704896540
transform -1 0 23000 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _238_
timestamp 1704896540
transform -1 0 29808 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _239_
timestamp 1704896540
transform 1 0 3772 0 1 63104
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _240_
timestamp 1704896540
transform 1 0 23368 0 -1 66368
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _241_
timestamp 1704896540
transform -1 0 37352 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _242_
timestamp 1704896540
transform 1 0 24564 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _243_
timestamp 1704896540
transform -1 0 31556 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _244_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 19596 0 1 62016
box -38 -48 682 592
use sky130_fd_sc_hd__buf_8  _245_
timestamp 1704896540
transform 1 0 24932 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__a211oi_2  _246_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 24656 0 1 43520
box -38 -48 958 592
use sky130_fd_sc_hd__or2_2  _247_
timestamp 1704896540
transform 1 0 14260 0 -1 64192
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_4  _248_
timestamp 1704896540
transform 1 0 28612 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__and3_2  _249_
timestamp 1704896540
transform 1 0 39836 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _250_
timestamp 1704896540
transform 1 0 6440 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _251_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8924 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _252_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11132 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _253_
timestamp 1704896540
transform -1 0 30636 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_2  _254_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 31832 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _255_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 18124 0 -1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_2  _256_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2576 0 1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__and4_4  _257_
timestamp 1704896540
transform 1 0 5336 0 -1 57664
box -38 -48 866 592
use sky130_fd_sc_hd__and2_4  _258_
timestamp 1704896540
transform -1 0 18676 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _259_
timestamp 1704896540
transform -1 0 4876 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_2  _260_
timestamp 1704896540
transform 1 0 14628 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _261_
timestamp 1704896540
transform -1 0 21712 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _262_
timestamp 1704896540
transform 1 0 8924 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _263_
timestamp 1704896540
transform 1 0 36708 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _264_
timestamp 1704896540
transform 1 0 36432 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _265_
timestamp 1704896540
transform 1 0 1656 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _266_
timestamp 1704896540
transform 1 0 37812 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__and4_4  _267_
timestamp 1704896540
transform 1 0 6348 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a211oi_4  _268_
timestamp 1704896540
transform -1 0 33948 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__or2_2  _269_
timestamp 1704896540
transform -1 0 32568 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_4  _270_
timestamp 1704896540
transform -1 0 7544 0 -1 68544
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _271_
timestamp 1704896540
transform -1 0 24840 0 1 48960
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _272_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 22080 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _273_
timestamp 1704896540
transform -1 0 22080 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _274_
timestamp 1704896540
transform 1 0 33856 0 1 47872
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_4  _275_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7544 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__a21oi_4  _276_
timestamp 1704896540
transform -1 0 30728 0 1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__and3_4  _277_
timestamp 1704896540
transform 1 0 33488 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__nor3_2  _278_
timestamp 1704896540
transform -1 0 32844 0 -1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _279_
timestamp 1704896540
transform 1 0 34132 0 1 67456
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _280_
timestamp 1704896540
transform 1 0 20516 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__and3_2  _281_
timestamp 1704896540
transform -1 0 26588 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _282_
timestamp 1704896540
transform -1 0 3680 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _283_
timestamp 1704896540
transform 1 0 7176 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _284_
timestamp 1704896540
transform -1 0 17296 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_4  _285_
timestamp 1704896540
transform 1 0 20884 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_4  _286_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 38732 0 1 62016
box -38 -48 958 592
use sky130_fd_sc_hd__a2111o_4  _287_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 15824 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__nor2_1  _288_
timestamp 1704896540
transform -1 0 24196 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _289_
timestamp 1704896540
transform 1 0 34868 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__or3_4  _290_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10764 0 -1 52224
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _291_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 39100 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _292_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 39836 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _293_
timestamp 1704896540
transform -1 0 6440 0 1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__a21boi_2  _294_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 30452 0 -1 57664
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  _295_
timestamp 1704896540
transform -1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _296_
timestamp 1704896540
transform -1 0 26312 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _297_
timestamp 1704896540
transform -1 0 6532 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _298_
timestamp 1704896540
transform -1 0 25668 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _299_
timestamp 1704896540
transform -1 0 19596 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _300_
timestamp 1704896540
transform 1 0 6992 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _301_
timestamp 1704896540
transform 1 0 26956 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _302_
timestamp 1704896540
transform -1 0 21252 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _303_
timestamp 1704896540
transform 1 0 8924 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _304_
timestamp 1704896540
transform 1 0 7544 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _305_
timestamp 1704896540
transform 1 0 14536 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _306_
timestamp 1704896540
transform -1 0 11040 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _307_
timestamp 1704896540
transform 1 0 16468 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _308_
timestamp 1704896540
transform -1 0 27876 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _309_
timestamp 1704896540
transform -1 0 28152 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _310_
timestamp 1704896540
transform 1 0 32476 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _311_
timestamp 1704896540
transform -1 0 1932 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _312_
timestamp 1704896540
transform -1 0 14444 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _313_
timestamp 1704896540
transform 1 0 29532 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _314_
timestamp 1704896540
transform -1 0 8372 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _315_
timestamp 1704896540
transform -1 0 21068 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _316_
timestamp 1704896540
transform 1 0 4600 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _317_
timestamp 1704896540
transform -1 0 30636 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _318_
timestamp 1704896540
transform -1 0 31004 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _319_
timestamp 1704896540
transform -1 0 36524 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _320_
timestamp 1704896540
transform 1 0 15364 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _321_
timestamp 1704896540
transform -1 0 24932 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _322_
timestamp 1704896540
transform -1 0 10580 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _323_
timestamp 1704896540
transform -1 0 40020 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _324_
timestamp 1704896540
transform 1 0 19964 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _325_
timestamp 1704896540
transform 1 0 18584 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _326_
timestamp 1704896540
transform 1 0 40296 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _327_
timestamp 1704896540
transform -1 0 28704 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _328_
timestamp 1704896540
transform 1 0 10212 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _329_
timestamp 1704896540
transform -1 0 35328 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _330_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11868 0 1 25024
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _331_
timestamp 1704896540
transform -1 0 25024 0 -1 53312
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _332_
timestamp 1704896540
transform 1 0 5980 0 1 56576
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _333_
timestamp 1704896540
transform 1 0 7268 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _334_
timestamp 1704896540
transform 1 0 36892 0 1 41344
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _335_
timestamp 1704896540
transform -1 0 32200 0 1 53312
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _336_
timestamp 1704896540
transform -1 0 8096 0 1 29376
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _337_
timestamp 1704896540
transform -1 0 11960 0 1 30464
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _338_
timestamp 1704896540
transform 1 0 12604 0 -1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _339_
timestamp 1704896540
transform 1 0 37260 0 -1 56576
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _340_
timestamp 1704896540
transform 1 0 37260 0 -1 32640
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _341_
timestamp 1704896540
transform 1 0 24748 0 1 41344
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _342_
timestamp 1704896540
transform 1 0 22540 0 -1 21760
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _343_
timestamp 1704896540
transform -1 0 17940 0 1 27200
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _344_
timestamp 1704896540
transform 1 0 37628 0 1 50048
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _345_
timestamp 1704896540
transform 1 0 3864 0 -1 29376
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _346_
timestamp 1704896540
transform 1 0 31096 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _347_
timestamp 1704896540
transform -1 0 5336 0 -1 57664
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _348_
timestamp 1704896540
transform 1 0 18216 0 -1 29376
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _349_
timestamp 1704896540
transform -1 0 21344 0 1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _350_
timestamp 1704896540
transform 1 0 6624 0 -1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _351_
timestamp 1704896540
transform 1 0 34132 0 -1 57664
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _352_
timestamp 1704896540
transform 1 0 23460 0 -1 25024
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _353_
timestamp 1704896540
transform 1 0 21804 0 -1 39168
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _354_
timestamp 1704896540
transform 1 0 7820 0 -1 36992
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _355_
timestamp 1704896540
transform 1 0 9568 0 1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _356_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 37720 0 1 53312
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _357_
timestamp 1704896540
transform 1 0 30820 0 1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _358_
timestamp 1704896540
transform -1 0 5060 0 -1 20672
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _359_
timestamp 1704896540
transform 1 0 8372 0 -1 54400
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _360_
timestamp 1704896540
transform 1 0 18860 0 -1 31552
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _361_
timestamp 1704896540
transform -1 0 3496 0 -1 45696
box -38 -48 2154 592
use sky130_fd_sc_hd__buf_2  _370_
timestamp 1704896540
transform -1 0 9292 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 11684 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1704896540
transform -1 0 3680 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1704896540
transform -1 0 30912 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1704896540
transform -1 0 24288 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1704896540
transform -1 0 7636 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1704896540
transform 1 0 33028 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1704896540
transform -1 0 7452 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1704896540
transform -1 0 7084 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1704896540
transform -1 0 36708 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1704896540
transform -1 0 15640 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1704896540
transform -1 0 9384 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1704896540
transform -1 0 2760 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1704896540
transform -1 0 3864 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1704896540
transform 1 0 5244 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1704896540
transform 1 0 18492 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1704896540
transform -1 0 19964 0 1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1704896540
transform 1 0 34316 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1704896540
transform 1 0 36248 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1704896540
transform 1 0 32752 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1704896540
transform -1 0 34040 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1704896540
transform -1 0 12788 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1704896540
transform 1 0 3864 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1704896540
transform -1 0 18492 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1704896540
transform 1 0 28796 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1704896540
transform 1 0 28796 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1704896540
transform -1 0 5520 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1704896540
transform 1 0 23000 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 1704896540
transform -1 0 36616 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp 1704896540
transform -1 0 39192 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp 1704896540
transform 1 0 6440 0 1 65280
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp 1704896540
transform 1 0 14260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp 1704896540
transform 1 0 33488 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_33
timestamp 1704896540
transform 1 0 36064 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_34
timestamp 1704896540
transform -1 0 25208 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_35
timestamp 1704896540
transform -1 0 3220 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_36
timestamp 1704896540
transform 1 0 38732 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_37
timestamp 1704896540
transform 1 0 29808 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_38
timestamp 1704896540
transform -1 0 35788 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_39
timestamp 1704896540
transform -1 0 16284 0 1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_40
timestamp 1704896540
transform -1 0 37168 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_41
timestamp 1704896540
transform 1 0 7360 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_42
timestamp 1704896540
transform -1 0 4416 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_43
timestamp 1704896540
transform 1 0 25944 0 1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_44
timestamp 1704896540
transform 1 0 39376 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_45
timestamp 1704896540
transform 1 0 28428 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_46
timestamp 1704896540
transform 1 0 39376 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_47
timestamp 1704896540
transform 1 0 36800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_48
timestamp 1704896540
transform -1 0 22448 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_49
timestamp 1704896540
transform 1 0 33120 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_50
timestamp 1704896540
transform -1 0 4416 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_51
timestamp 1704896540
transform 1 0 36616 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_52
timestamp 1704896540
transform -1 0 37904 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_53
timestamp 1704896540
transform 1 0 4600 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 19596 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1704896540
transform -1 0 11132 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1704896540
transform 1 0 24564 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1704896540
transform 1 0 14536 0 1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1704896540
transform 1 0 28796 0 -1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  clkload0
timestamp 1704896540
transform 1 0 24564 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  clkload1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 14168 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  clkload2
timestamp 1704896540
transform 1 0 28796 0 1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2484 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_20 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2944 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1704896540
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1704896540
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1704896540
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_69 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_73 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7820 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_77 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_83
timestamp 1704896540
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1704896540
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1704896540
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1704896540
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1704896540
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_125
timestamp 1704896540
transform 1 0 12604 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_134
timestamp 1704896540
transform 1 0 13432 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1704896540
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1704896540
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1704896540
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1704896540
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_181
timestamp 1704896540
transform 1 0 17756 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_187
timestamp 1704896540
transform 1 0 18308 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_191
timestamp 1704896540
transform 1 0 18676 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_195
timestamp 1704896540
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1704896540
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 1704896540
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1704896540
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1704896540
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_237
timestamp 1704896540
transform 1 0 22908 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_248
timestamp 1704896540
transform 1 0 23920 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1704896540
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 1704896540
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 1704896540
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 1704896540
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_293
timestamp 1704896540
transform 1 0 28060 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_301
timestamp 1704896540
transform 1 0 28796 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 1704896540
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 1704896540
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_321
timestamp 1704896540
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_333
timestamp 1704896540
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_337
timestamp 1704896540
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_349
timestamp 1704896540
transform 1 0 33212 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_357
timestamp 1704896540
transform 1 0 33948 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_362
timestamp 1704896540
transform 1 0 34408 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_365
timestamp 1704896540
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_377
timestamp 1704896540
transform 1 0 35788 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_385
timestamp 1704896540
transform 1 0 36524 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_393
timestamp 1704896540
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_405
timestamp 1704896540
transform 1 0 38364 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_411
timestamp 1704896540
transform 1 0 38916 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_419
timestamp 1704896540
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_424
timestamp 1704896540
transform 1 0 40112 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_428
timestamp 1704896540
transform 1 0 40480 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1704896540
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1704896540
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1704896540
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1704896540
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1704896540
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1704896540
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1704896540
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_69
timestamp 1704896540
transform 1 0 7452 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_99
timestamp 1704896540
transform 1 0 10212 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1704896540
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1704896540
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1704896540
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_137
timestamp 1704896540
transform 1 0 13708 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_145
timestamp 1704896540
transform 1 0 14444 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_153
timestamp 1704896540
transform 1 0 15180 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_165
timestamp 1704896540
transform 1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1704896540
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1704896540
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1704896540
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1704896540
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 1704896540
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1704896540
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1704896540
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1704896540
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1704896540
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 1704896540
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 1704896540
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1704896540
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1704896540
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1704896540
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 1704896540
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_317
timestamp 1704896540
transform 1 0 30268 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_331
timestamp 1704896540
transform 1 0 31556 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 1704896540
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_337
timestamp 1704896540
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_349
timestamp 1704896540
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_361
timestamp 1704896540
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_373
timestamp 1704896540
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_385
timestamp 1704896540
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_391
timestamp 1704896540
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_393
timestamp 1704896540
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_405
timestamp 1704896540
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_417
timestamp 1704896540
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_3
timestamp 1704896540
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_22
timestamp 1704896540
transform 1 0 3128 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1704896540
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1704896540
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_53
timestamp 1704896540
transform 1 0 5980 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_61
timestamp 1704896540
transform 1 0 6716 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_67
timestamp 1704896540
transform 1 0 7268 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_79
timestamp 1704896540
transform 1 0 8372 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1704896540
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1704896540
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1704896540
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1704896540
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1704896540
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1704896540
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1704896540
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1704896540
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1704896540
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1704896540
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1704896540
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1704896540
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1704896540
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1704896540
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1704896540
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1704896540
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1704896540
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 1704896540
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1704896540
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1704896540
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1704896540
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1704896540
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 1704896540
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 1704896540
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1704896540
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1704896540
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 1704896540
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_333
timestamp 1704896540
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_345
timestamp 1704896540
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_357
timestamp 1704896540
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_363
timestamp 1704896540
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_365
timestamp 1704896540
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_377
timestamp 1704896540
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_389
timestamp 1704896540
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_401
timestamp 1704896540
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_413
timestamp 1704896540
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_419
timestamp 1704896540
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_421
timestamp 1704896540
transform 1 0 39836 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1704896540
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1704896540
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1704896540
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1704896540
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1704896540
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1704896540
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1704896540
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1704896540
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1704896540
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1704896540
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1704896540
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1704896540
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1704896540
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1704896540
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1704896540
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1704896540
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1704896540
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1704896540
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1704896540
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1704896540
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1704896540
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1704896540
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1704896540
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1704896540
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1704896540
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1704896540
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1704896540
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1704896540
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 1704896540
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1704896540
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1704896540
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1704896540
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1704896540
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 1704896540
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_329
timestamp 1704896540
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_335
timestamp 1704896540
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 1704896540
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 1704896540
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_361
timestamp 1704896540
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_373
timestamp 1704896540
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_385
timestamp 1704896540
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_391
timestamp 1704896540
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_393
timestamp 1704896540
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_405
timestamp 1704896540
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_417
timestamp 1704896540
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_3
timestamp 1704896540
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_9
timestamp 1704896540
transform 1 0 1932 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_21
timestamp 1704896540
transform 1 0 3036 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1704896540
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1704896540
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1704896540
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_53
timestamp 1704896540
transform 1 0 5980 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_57
timestamp 1704896540
transform 1 0 6348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_69
timestamp 1704896540
transform 1 0 7452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_81
timestamp 1704896540
transform 1 0 8556 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1704896540
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1704896540
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1704896540
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1704896540
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1704896540
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1704896540
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1704896540
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1704896540
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1704896540
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1704896540
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1704896540
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1704896540
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1704896540
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1704896540
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1704896540
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1704896540
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1704896540
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1704896540
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_253
timestamp 1704896540
transform 1 0 24380 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_261
timestamp 1704896540
transform 1 0 25116 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_272
timestamp 1704896540
transform 1 0 26128 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_284
timestamp 1704896540
transform 1 0 27232 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_296
timestamp 1704896540
transform 1 0 28336 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1704896540
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 1704896540
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_333
timestamp 1704896540
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_345
timestamp 1704896540
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_357
timestamp 1704896540
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_363
timestamp 1704896540
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_365
timestamp 1704896540
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_377
timestamp 1704896540
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_389
timestamp 1704896540
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_401
timestamp 1704896540
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_413
timestamp 1704896540
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_419
timestamp 1704896540
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_421
timestamp 1704896540
transform 1 0 39836 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1704896540
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1704896540
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1704896540
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1704896540
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1704896540
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1704896540
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1704896540
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1704896540
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1704896540
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1704896540
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1704896540
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1704896540
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1704896540
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1704896540
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1704896540
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1704896540
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1704896540
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1704896540
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1704896540
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1704896540
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1704896540
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_205
timestamp 1704896540
transform 1 0 19964 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_213
timestamp 1704896540
transform 1 0 20700 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_219
timestamp 1704896540
transform 1 0 21252 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1704896540
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1704896540
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1704896540
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1704896540
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1704896540
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1704896540
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1704896540
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1704896540
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1704896540
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1704896540
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 1704896540
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_329
timestamp 1704896540
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 1704896540
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 1704896540
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_349
timestamp 1704896540
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_361
timestamp 1704896540
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_373
timestamp 1704896540
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_385
timestamp 1704896540
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_391
timestamp 1704896540
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_393
timestamp 1704896540
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_405
timestamp 1704896540
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_417
timestamp 1704896540
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1704896540
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1704896540
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1704896540
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1704896540
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1704896540
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1704896540
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1704896540
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1704896540
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1704896540
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1704896540
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1704896540
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1704896540
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1704896540
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1704896540
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1704896540
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1704896540
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1704896540
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1704896540
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1704896540
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1704896540
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1704896540
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1704896540
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1704896540
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1704896540
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1704896540
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1704896540
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1704896540
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1704896540
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1704896540
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1704896540
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1704896540
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1704896540
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1704896540
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1704896540
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 1704896540
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_333
timestamp 1704896540
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_345
timestamp 1704896540
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_357
timestamp 1704896540
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_363
timestamp 1704896540
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_365
timestamp 1704896540
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_377
timestamp 1704896540
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_389
timestamp 1704896540
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_401
timestamp 1704896540
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_413
timestamp 1704896540
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_419
timestamp 1704896540
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_421
timestamp 1704896540
transform 1 0 39836 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1704896540
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1704896540
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1704896540
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1704896540
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1704896540
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1704896540
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1704896540
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1704896540
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1704896540
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1704896540
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1704896540
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1704896540
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1704896540
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1704896540
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1704896540
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1704896540
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1704896540
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1704896540
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1704896540
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1704896540
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1704896540
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1704896540
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1704896540
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1704896540
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1704896540
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1704896540
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1704896540
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1704896540
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 1704896540
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1704896540
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1704896540
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1704896540
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1704896540
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1704896540
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_329
timestamp 1704896540
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_335
timestamp 1704896540
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_337
timestamp 1704896540
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_349
timestamp 1704896540
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_361
timestamp 1704896540
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_373
timestamp 1704896540
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_385
timestamp 1704896540
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_391
timestamp 1704896540
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_393
timestamp 1704896540
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_405
timestamp 1704896540
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_417
timestamp 1704896540
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1704896540
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1704896540
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1704896540
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1704896540
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1704896540
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1704896540
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1704896540
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1704896540
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1704896540
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1704896540
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1704896540
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1704896540
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1704896540
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1704896540
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1704896540
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1704896540
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1704896540
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1704896540
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1704896540
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1704896540
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1704896540
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1704896540
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1704896540
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1704896540
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1704896540
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 1704896540
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1704896540
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1704896540
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1704896540
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1704896540
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 1704896540
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 1704896540
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 1704896540
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1704896540
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_321
timestamp 1704896540
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_333
timestamp 1704896540
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_345
timestamp 1704896540
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_357
timestamp 1704896540
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_363
timestamp 1704896540
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_365
timestamp 1704896540
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_377
timestamp 1704896540
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_389
timestamp 1704896540
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_401
timestamp 1704896540
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_413
timestamp 1704896540
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_419
timestamp 1704896540
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_421
timestamp 1704896540
transform 1 0 39836 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1704896540
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1704896540
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1704896540
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1704896540
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1704896540
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1704896540
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1704896540
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1704896540
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1704896540
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1704896540
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1704896540
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1704896540
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1704896540
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1704896540
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1704896540
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1704896540
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1704896540
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1704896540
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1704896540
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1704896540
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 1704896540
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_205
timestamp 1704896540
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 1704896540
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1704896540
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1704896540
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 1704896540
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 1704896540
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 1704896540
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_273
timestamp 1704896540
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1704896540
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1704896540
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 1704896540
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_305
timestamp 1704896540
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_317
timestamp 1704896540
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_329
timestamp 1704896540
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_335
timestamp 1704896540
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_337
timestamp 1704896540
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_349
timestamp 1704896540
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_361
timestamp 1704896540
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_373
timestamp 1704896540
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_385
timestamp 1704896540
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_391
timestamp 1704896540
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_393
timestamp 1704896540
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_405
timestamp 1704896540
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_417
timestamp 1704896540
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1704896540
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1704896540
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1704896540
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1704896540
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1704896540
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1704896540
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1704896540
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1704896540
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1704896540
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_88
timestamp 1704896540
transform 1 0 9200 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_100
timestamp 1704896540
transform 1 0 10304 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_112
timestamp 1704896540
transform 1 0 11408 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_124
timestamp 1704896540
transform 1 0 12512 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_136
timestamp 1704896540
transform 1 0 13616 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1704896540
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1704896540
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1704896540
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_177
timestamp 1704896540
transform 1 0 17388 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_185
timestamp 1704896540
transform 1 0 18124 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_189
timestamp 1704896540
transform 1 0 18492 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_194
timestamp 1704896540
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1704896540
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1704896540
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 1704896540
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_233
timestamp 1704896540
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_245
timestamp 1704896540
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1704896540
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1704896540
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 1704896540
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_277
timestamp 1704896540
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_289
timestamp 1704896540
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_301
timestamp 1704896540
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 1704896540
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 1704896540
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_321
timestamp 1704896540
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_333
timestamp 1704896540
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_345
timestamp 1704896540
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_357
timestamp 1704896540
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_363
timestamp 1704896540
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_365
timestamp 1704896540
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_377
timestamp 1704896540
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_389
timestamp 1704896540
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_401
timestamp 1704896540
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_413
timestamp 1704896540
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_419
timestamp 1704896540
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_421
timestamp 1704896540
transform 1 0 39836 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1704896540
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1704896540
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1704896540
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1704896540
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1704896540
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1704896540
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1704896540
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1704896540
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1704896540
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1704896540
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1704896540
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1704896540
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1704896540
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1704896540
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 1704896540
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 1704896540
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 1704896540
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1704896540
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 1704896540
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_181
timestamp 1704896540
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_193
timestamp 1704896540
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_205
timestamp 1704896540
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_217
timestamp 1704896540
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1704896540
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1704896540
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_237
timestamp 1704896540
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_249
timestamp 1704896540
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_261
timestamp 1704896540
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_273
timestamp 1704896540
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 1704896540
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 1704896540
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 1704896540
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_305
timestamp 1704896540
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_317
timestamp 1704896540
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_329
timestamp 1704896540
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_335
timestamp 1704896540
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_337
timestamp 1704896540
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_349
timestamp 1704896540
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_361
timestamp 1704896540
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_373
timestamp 1704896540
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_385
timestamp 1704896540
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_391
timestamp 1704896540
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_393
timestamp 1704896540
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_405
timestamp 1704896540
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_417
timestamp 1704896540
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1704896540
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1704896540
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1704896540
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1704896540
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1704896540
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1704896540
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_65
timestamp 1704896540
transform 1 0 7084 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_69
timestamp 1704896540
transform 1 0 7452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_81
timestamp 1704896540
transform 1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1704896540
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1704896540
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 1704896540
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 1704896540
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1704896540
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1704896540
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1704896540
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 1704896540
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 1704896540
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_177
timestamp 1704896540
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_189
timestamp 1704896540
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1704896540
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 1704896540
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_209
timestamp 1704896540
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_221
timestamp 1704896540
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_233
timestamp 1704896540
transform 1 0 22540 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_238
timestamp 1704896540
transform 1 0 23000 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_250
timestamp 1704896540
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 1704896540
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_265
timestamp 1704896540
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_277
timestamp 1704896540
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_289
timestamp 1704896540
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_301
timestamp 1704896540
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 1704896540
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 1704896540
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_321
timestamp 1704896540
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_333
timestamp 1704896540
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_345
timestamp 1704896540
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_357
timestamp 1704896540
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_363
timestamp 1704896540
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_365
timestamp 1704896540
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_377
timestamp 1704896540
transform 1 0 35788 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_385
timestamp 1704896540
transform 1 0 36524 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_390
timestamp 1704896540
transform 1 0 36984 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_397
timestamp 1704896540
transform 1 0 37628 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_409
timestamp 1704896540
transform 1 0 38732 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_417
timestamp 1704896540
transform 1 0 39468 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_421
timestamp 1704896540
transform 1 0 39836 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1704896540
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1704896540
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1704896540
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1704896540
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1704896540
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1704896540
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_57
timestamp 1704896540
transform 1 0 6348 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_65
timestamp 1704896540
transform 1 0 7084 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_90
timestamp 1704896540
transform 1 0 9384 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_102
timestamp 1704896540
transform 1 0 10488 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_110
timestamp 1704896540
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 1704896540
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 1704896540
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_137
timestamp 1704896540
transform 1 0 13708 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_145
timestamp 1704896540
transform 1 0 14444 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_149
timestamp 1704896540
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_161
timestamp 1704896540
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1704896540
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 1704896540
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_181
timestamp 1704896540
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_193
timestamp 1704896540
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_205
timestamp 1704896540
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_217
timestamp 1704896540
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 1704896540
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_225
timestamp 1704896540
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_237
timestamp 1704896540
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_249
timestamp 1704896540
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_261
timestamp 1704896540
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_273
timestamp 1704896540
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_279
timestamp 1704896540
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_281
timestamp 1704896540
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_293
timestamp 1704896540
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_305
timestamp 1704896540
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_317
timestamp 1704896540
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_329
timestamp 1704896540
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_335
timestamp 1704896540
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_337
timestamp 1704896540
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_349
timestamp 1704896540
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_361
timestamp 1704896540
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_373
timestamp 1704896540
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_385
timestamp 1704896540
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_391
timestamp 1704896540
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_393
timestamp 1704896540
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_405
timestamp 1704896540
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_417
timestamp 1704896540
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1704896540
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1704896540
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1704896540
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1704896540
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1704896540
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1704896540
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 1704896540
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 1704896540
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1704896540
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1704896540
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 1704896540
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_109
timestamp 1704896540
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_121
timestamp 1704896540
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 1704896540
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1704896540
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 1704896540
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_153
timestamp 1704896540
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_165
timestamp 1704896540
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_177
timestamp 1704896540
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_189
timestamp 1704896540
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 1704896540
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_197
timestamp 1704896540
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_209
timestamp 1704896540
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_221
timestamp 1704896540
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_233
timestamp 1704896540
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_245
timestamp 1704896540
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_251
timestamp 1704896540
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_253
timestamp 1704896540
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_265
timestamp 1704896540
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_277
timestamp 1704896540
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_289
timestamp 1704896540
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_301
timestamp 1704896540
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_307
timestamp 1704896540
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_309
timestamp 1704896540
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_321
timestamp 1704896540
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_333
timestamp 1704896540
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_345
timestamp 1704896540
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_357
timestamp 1704896540
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_363
timestamp 1704896540
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_365
timestamp 1704896540
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_377
timestamp 1704896540
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_389
timestamp 1704896540
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_401
timestamp 1704896540
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_413
timestamp 1704896540
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_419
timestamp 1704896540
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_421
timestamp 1704896540
transform 1 0 39836 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1704896540
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1704896540
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1704896540
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_39
timestamp 1704896540
transform 1 0 4692 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_45
timestamp 1704896540
transform 1 0 5244 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_48
timestamp 1704896540
transform 1 0 5520 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_53
timestamp 1704896540
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1704896540
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 1704896540
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_81
timestamp 1704896540
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_93
timestamp 1704896540
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 1704896540
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1704896540
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1704896540
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 1704896540
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_137
timestamp 1704896540
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_149
timestamp 1704896540
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_161
timestamp 1704896540
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1704896540
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_169
timestamp 1704896540
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_181
timestamp 1704896540
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_193
timestamp 1704896540
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_205
timestamp 1704896540
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_217
timestamp 1704896540
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_223
timestamp 1704896540
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_225
timestamp 1704896540
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_237
timestamp 1704896540
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_249
timestamp 1704896540
transform 1 0 24012 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_259
timestamp 1704896540
transform 1 0 24932 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_271
timestamp 1704896540
transform 1 0 26036 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_279
timestamp 1704896540
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_281
timestamp 1704896540
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_293
timestamp 1704896540
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_305
timestamp 1704896540
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_317
timestamp 1704896540
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_329
timestamp 1704896540
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_335
timestamp 1704896540
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_359
timestamp 1704896540
transform 1 0 34132 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_371
timestamp 1704896540
transform 1 0 35236 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_383
timestamp 1704896540
transform 1 0 36340 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_391
timestamp 1704896540
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_393
timestamp 1704896540
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_405
timestamp 1704896540
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_417
timestamp 1704896540
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1704896540
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1704896540
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1704896540
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1704896540
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1704896540
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 1704896540
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 1704896540
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 1704896540
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1704896540
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1704896540
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_97
timestamp 1704896540
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_109
timestamp 1704896540
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_121
timestamp 1704896540
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_133
timestamp 1704896540
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1704896540
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_141
timestamp 1704896540
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_153
timestamp 1704896540
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_165
timestamp 1704896540
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_177
timestamp 1704896540
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_189
timestamp 1704896540
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 1704896540
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_197
timestamp 1704896540
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_209
timestamp 1704896540
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_221
timestamp 1704896540
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_233
timestamp 1704896540
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_245
timestamp 1704896540
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_251
timestamp 1704896540
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_253
timestamp 1704896540
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_265
timestamp 1704896540
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_277
timestamp 1704896540
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_289
timestamp 1704896540
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_301
timestamp 1704896540
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_307
timestamp 1704896540
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_309
timestamp 1704896540
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_321
timestamp 1704896540
transform 1 0 30636 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_324
timestamp 1704896540
transform 1 0 30912 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_349
timestamp 1704896540
transform 1 0 33212 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_361
timestamp 1704896540
transform 1 0 34316 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_365
timestamp 1704896540
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_377
timestamp 1704896540
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_389
timestamp 1704896540
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_401
timestamp 1704896540
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_413
timestamp 1704896540
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_419
timestamp 1704896540
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_421
timestamp 1704896540
transform 1 0 39836 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1704896540
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1704896540
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1704896540
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 1704896540
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 1704896540
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1704896540
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1704896540
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1704896540
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 1704896540
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_93
timestamp 1704896540
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_105
timestamp 1704896540
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1704896540
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 1704896540
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_125
timestamp 1704896540
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_137
timestamp 1704896540
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_149
timestamp 1704896540
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_161
timestamp 1704896540
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp 1704896540
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_169
timestamp 1704896540
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_181
timestamp 1704896540
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_193
timestamp 1704896540
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_205
timestamp 1704896540
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_217
timestamp 1704896540
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_223
timestamp 1704896540
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_225
timestamp 1704896540
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_237
timestamp 1704896540
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_249
timestamp 1704896540
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_261
timestamp 1704896540
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_273
timestamp 1704896540
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_279
timestamp 1704896540
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_281
timestamp 1704896540
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_293
timestamp 1704896540
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_305
timestamp 1704896540
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_317
timestamp 1704896540
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_329
timestamp 1704896540
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_335
timestamp 1704896540
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_337
timestamp 1704896540
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_349
timestamp 1704896540
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_361
timestamp 1704896540
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_373
timestamp 1704896540
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_385
timestamp 1704896540
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_391
timestamp 1704896540
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_393
timestamp 1704896540
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_405
timestamp 1704896540
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_417
timestamp 1704896540
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1704896540
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1704896540
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1704896540
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_29
timestamp 1704896540
transform 1 0 3772 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_37
timestamp 1704896540
transform 1 0 4508 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1704896540
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 1704896540
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_65
timestamp 1704896540
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_77
timestamp 1704896540
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1704896540
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1704896540
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_97
timestamp 1704896540
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_109
timestamp 1704896540
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_121
timestamp 1704896540
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_133
timestamp 1704896540
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1704896540
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 1704896540
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_153
timestamp 1704896540
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_165
timestamp 1704896540
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_177
timestamp 1704896540
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_189
timestamp 1704896540
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_195
timestamp 1704896540
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_197
timestamp 1704896540
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_209
timestamp 1704896540
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_221
timestamp 1704896540
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_233
timestamp 1704896540
transform 1 0 22540 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_241
timestamp 1704896540
transform 1 0 23276 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_249
timestamp 1704896540
transform 1 0 24012 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_253
timestamp 1704896540
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_265
timestamp 1704896540
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_277
timestamp 1704896540
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_289
timestamp 1704896540
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_301
timestamp 1704896540
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_307
timestamp 1704896540
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_309
timestamp 1704896540
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_321
timestamp 1704896540
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_333
timestamp 1704896540
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_345
timestamp 1704896540
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_357
timestamp 1704896540
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_363
timestamp 1704896540
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_365
timestamp 1704896540
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_377
timestamp 1704896540
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_389
timestamp 1704896540
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_401
timestamp 1704896540
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_413
timestamp 1704896540
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_419
timestamp 1704896540
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_421
timestamp 1704896540
transform 1 0 39836 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1704896540
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1704896540
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1704896540
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 1704896540
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 1704896540
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1704896540
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 1704896540
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_69
timestamp 1704896540
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_81
timestamp 1704896540
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_93
timestamp 1704896540
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_105
timestamp 1704896540
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1704896540
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_113
timestamp 1704896540
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_125
timestamp 1704896540
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_137
timestamp 1704896540
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_149
timestamp 1704896540
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_161
timestamp 1704896540
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 1704896540
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_169
timestamp 1704896540
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_181
timestamp 1704896540
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_193
timestamp 1704896540
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_205
timestamp 1704896540
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_217
timestamp 1704896540
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_223
timestamp 1704896540
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_225
timestamp 1704896540
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_237
timestamp 1704896540
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_249
timestamp 1704896540
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_261
timestamp 1704896540
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_273
timestamp 1704896540
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_279
timestamp 1704896540
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_281
timestamp 1704896540
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_293
timestamp 1704896540
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_305
timestamp 1704896540
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_317
timestamp 1704896540
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_329
timestamp 1704896540
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_335
timestamp 1704896540
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_337
timestamp 1704896540
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_349
timestamp 1704896540
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_361
timestamp 1704896540
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_373
timestamp 1704896540
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_385
timestamp 1704896540
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_391
timestamp 1704896540
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_393
timestamp 1704896540
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_405
timestamp 1704896540
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_417
timestamp 1704896540
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1704896540
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1704896540
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1704896540
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1704896540
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1704896540
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_53
timestamp 1704896540
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_65
timestamp 1704896540
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_77
timestamp 1704896540
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1704896540
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 1704896540
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_97
timestamp 1704896540
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_109
timestamp 1704896540
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_121
timestamp 1704896540
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_133
timestamp 1704896540
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 1704896540
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 1704896540
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_153
timestamp 1704896540
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_165
timestamp 1704896540
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_177
timestamp 1704896540
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_189
timestamp 1704896540
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 1704896540
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_197
timestamp 1704896540
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_209
timestamp 1704896540
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_221
timestamp 1704896540
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_233
timestamp 1704896540
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_245
timestamp 1704896540
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_251
timestamp 1704896540
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_253
timestamp 1704896540
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_265
timestamp 1704896540
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_277
timestamp 1704896540
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_289
timestamp 1704896540
transform 1 0 27692 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_294
timestamp 1704896540
transform 1 0 28152 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_306
timestamp 1704896540
transform 1 0 29256 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_309
timestamp 1704896540
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_321
timestamp 1704896540
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_333
timestamp 1704896540
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_345
timestamp 1704896540
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_357
timestamp 1704896540
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_363
timestamp 1704896540
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_365
timestamp 1704896540
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_377
timestamp 1704896540
transform 1 0 35788 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_390
timestamp 1704896540
transform 1 0 36984 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_402
timestamp 1704896540
transform 1 0 38088 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_414
timestamp 1704896540
transform 1 0 39192 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_421
timestamp 1704896540
transform 1 0 39836 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1704896540
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1704896540
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 1704896540
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_39
timestamp 1704896540
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 1704896540
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1704896540
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1704896540
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 1704896540
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_81
timestamp 1704896540
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_93
timestamp 1704896540
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_105
timestamp 1704896540
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1704896540
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1704896540
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_148
timestamp 1704896540
transform 1 0 14720 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_160
timestamp 1704896540
transform 1 0 15824 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp 1704896540
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_181
timestamp 1704896540
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_193
timestamp 1704896540
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_205
timestamp 1704896540
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_217
timestamp 1704896540
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp 1704896540
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_225
timestamp 1704896540
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_237
timestamp 1704896540
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_249
timestamp 1704896540
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_261
timestamp 1704896540
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_273
timestamp 1704896540
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_279
timestamp 1704896540
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_281
timestamp 1704896540
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_293
timestamp 1704896540
transform 1 0 28060 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_300
timestamp 1704896540
transform 1 0 28704 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_312
timestamp 1704896540
transform 1 0 29808 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_324
timestamp 1704896540
transform 1 0 30912 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_337
timestamp 1704896540
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_349
timestamp 1704896540
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_361
timestamp 1704896540
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_373
timestamp 1704896540
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_385
timestamp 1704896540
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_391
timestamp 1704896540
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_393
timestamp 1704896540
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_405
timestamp 1704896540
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_417
timestamp 1704896540
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1704896540
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1704896540
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1704896540
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1704896540
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1704896540
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 1704896540
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_65
timestamp 1704896540
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_77
timestamp 1704896540
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 1704896540
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 1704896540
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_97
timestamp 1704896540
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_109
timestamp 1704896540
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_121
timestamp 1704896540
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_133
timestamp 1704896540
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1704896540
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 1704896540
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_153
timestamp 1704896540
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_165
timestamp 1704896540
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_177
timestamp 1704896540
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_189
timestamp 1704896540
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 1704896540
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_197
timestamp 1704896540
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_209
timestamp 1704896540
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_221
timestamp 1704896540
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_233
timestamp 1704896540
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_245
timestamp 1704896540
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_251
timestamp 1704896540
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_253
timestamp 1704896540
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_265
timestamp 1704896540
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_277
timestamp 1704896540
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_289
timestamp 1704896540
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_301
timestamp 1704896540
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_307
timestamp 1704896540
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_309
timestamp 1704896540
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_321
timestamp 1704896540
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_333
timestamp 1704896540
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_345
timestamp 1704896540
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_357
timestamp 1704896540
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_363
timestamp 1704896540
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_365
timestamp 1704896540
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_377
timestamp 1704896540
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_389
timestamp 1704896540
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_401
timestamp 1704896540
transform 1 0 37996 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_412
timestamp 1704896540
transform 1 0 39008 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_421
timestamp 1704896540
transform 1 0 39836 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1704896540
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1704896540
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 1704896540
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 1704896540
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 1704896540
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1704896540
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1704896540
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_69
timestamp 1704896540
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_81
timestamp 1704896540
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_93
timestamp 1704896540
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_105
timestamp 1704896540
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1704896540
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 1704896540
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_125
timestamp 1704896540
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_137
timestamp 1704896540
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_149
timestamp 1704896540
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_161
timestamp 1704896540
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 1704896540
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_169
timestamp 1704896540
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_181
timestamp 1704896540
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_193
timestamp 1704896540
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_205
timestamp 1704896540
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_217
timestamp 1704896540
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 1704896540
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_225
timestamp 1704896540
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_237
timestamp 1704896540
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_249
timestamp 1704896540
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_261
timestamp 1704896540
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_273
timestamp 1704896540
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_279
timestamp 1704896540
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_281
timestamp 1704896540
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_293
timestamp 1704896540
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_305
timestamp 1704896540
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_317
timestamp 1704896540
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_329
timestamp 1704896540
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_335
timestamp 1704896540
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_342
timestamp 1704896540
transform 1 0 32568 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_354
timestamp 1704896540
transform 1 0 33672 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_366
timestamp 1704896540
transform 1 0 34776 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_378
timestamp 1704896540
transform 1 0 35880 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_390
timestamp 1704896540
transform 1 0 36984 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_393
timestamp 1704896540
transform 1 0 37260 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_406
timestamp 1704896540
transform 1 0 38456 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_418
timestamp 1704896540
transform 1 0 39560 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_426
timestamp 1704896540
transform 1 0 40296 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1704896540
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1704896540
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1704896540
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1704896540
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 1704896540
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_53
timestamp 1704896540
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_65
timestamp 1704896540
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_77
timestamp 1704896540
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1704896540
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1704896540
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_97
timestamp 1704896540
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_109
timestamp 1704896540
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_121
timestamp 1704896540
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_133
timestamp 1704896540
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1704896540
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_147
timestamp 1704896540
transform 1 0 14628 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_159
timestamp 1704896540
transform 1 0 15732 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_171
timestamp 1704896540
transform 1 0 16836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_183
timestamp 1704896540
transform 1 0 17940 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_195
timestamp 1704896540
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_197
timestamp 1704896540
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_209
timestamp 1704896540
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_221
timestamp 1704896540
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_233
timestamp 1704896540
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_245
timestamp 1704896540
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_251
timestamp 1704896540
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_253
timestamp 1704896540
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_265
timestamp 1704896540
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_277
timestamp 1704896540
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_289
timestamp 1704896540
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_301
timestamp 1704896540
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_307
timestamp 1704896540
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_309
timestamp 1704896540
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_321
timestamp 1704896540
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_333
timestamp 1704896540
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_345
timestamp 1704896540
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_357
timestamp 1704896540
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_363
timestamp 1704896540
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_365
timestamp 1704896540
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_377
timestamp 1704896540
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_389
timestamp 1704896540
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_401
timestamp 1704896540
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_413
timestamp 1704896540
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_419
timestamp 1704896540
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_421
timestamp 1704896540
transform 1 0 39836 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1704896540
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 1704896540
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 1704896540
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_39
timestamp 1704896540
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp 1704896540
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1704896540
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1704896540
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 1704896540
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_81
timestamp 1704896540
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_93
timestamp 1704896540
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_105
timestamp 1704896540
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1704896540
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 1704896540
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_125
timestamp 1704896540
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_137
timestamp 1704896540
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_149
timestamp 1704896540
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_161
timestamp 1704896540
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 1704896540
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 1704896540
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_181
timestamp 1704896540
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_193
timestamp 1704896540
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_205
timestamp 1704896540
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_217
timestamp 1704896540
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 1704896540
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_225
timestamp 1704896540
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_237
timestamp 1704896540
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_249
timestamp 1704896540
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_261
timestamp 1704896540
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_273
timestamp 1704896540
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_279
timestamp 1704896540
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_281
timestamp 1704896540
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_293
timestamp 1704896540
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_305
timestamp 1704896540
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_317
timestamp 1704896540
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_329
timestamp 1704896540
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_335
timestamp 1704896540
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_337
timestamp 1704896540
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_349
timestamp 1704896540
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_361
timestamp 1704896540
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_373
timestamp 1704896540
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_385
timestamp 1704896540
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_391
timestamp 1704896540
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_393
timestamp 1704896540
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_405
timestamp 1704896540
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_417
timestamp 1704896540
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1704896540
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1704896540
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1704896540
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1704896540
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 1704896540
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_53
timestamp 1704896540
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_65
timestamp 1704896540
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_77
timestamp 1704896540
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1704896540
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 1704896540
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_97
timestamp 1704896540
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_109
timestamp 1704896540
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_121
timestamp 1704896540
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_133
timestamp 1704896540
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1704896540
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_141
timestamp 1704896540
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_160
timestamp 1704896540
transform 1 0 15824 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_172
timestamp 1704896540
transform 1 0 16928 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_184
timestamp 1704896540
transform 1 0 18032 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_197
timestamp 1704896540
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_209
timestamp 1704896540
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_221
timestamp 1704896540
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_233
timestamp 1704896540
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_245
timestamp 1704896540
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_251
timestamp 1704896540
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_253
timestamp 1704896540
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_265
timestamp 1704896540
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_277
timestamp 1704896540
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_289
timestamp 1704896540
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_301
timestamp 1704896540
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_307
timestamp 1704896540
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_309
timestamp 1704896540
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_321
timestamp 1704896540
transform 1 0 30636 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_346
timestamp 1704896540
transform 1 0 32936 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_358
timestamp 1704896540
transform 1 0 34040 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_365
timestamp 1704896540
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_377
timestamp 1704896540
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_389
timestamp 1704896540
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_401
timestamp 1704896540
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_413
timestamp 1704896540
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_419
timestamp 1704896540
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_421
timestamp 1704896540
transform 1 0 39836 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1704896540
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_15
timestamp 1704896540
transform 1 0 2484 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_28
timestamp 1704896540
transform 1 0 3680 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_32
timestamp 1704896540
transform 1 0 4048 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_40
timestamp 1704896540
transform 1 0 4784 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_52
timestamp 1704896540
transform 1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1704896540
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_69
timestamp 1704896540
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_81
timestamp 1704896540
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_93
timestamp 1704896540
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_105
timestamp 1704896540
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 1704896540
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_113
timestamp 1704896540
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_125
timestamp 1704896540
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_137
timestamp 1704896540
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_149
timestamp 1704896540
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_161
timestamp 1704896540
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1704896540
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 1704896540
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_181
timestamp 1704896540
transform 1 0 17756 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_201
timestamp 1704896540
transform 1 0 19596 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_213
timestamp 1704896540
transform 1 0 20700 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_221
timestamp 1704896540
transform 1 0 21436 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_225
timestamp 1704896540
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_237
timestamp 1704896540
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_249
timestamp 1704896540
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_261
timestamp 1704896540
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_273
timestamp 1704896540
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_279
timestamp 1704896540
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_281
timestamp 1704896540
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_293
timestamp 1704896540
transform 1 0 28060 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_297
timestamp 1704896540
transform 1 0 28428 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_303
timestamp 1704896540
transform 1 0 28980 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_315
timestamp 1704896540
transform 1 0 30084 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_327
timestamp 1704896540
transform 1 0 31188 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_332
timestamp 1704896540
transform 1 0 31648 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_337
timestamp 1704896540
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_349
timestamp 1704896540
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_361
timestamp 1704896540
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_373
timestamp 1704896540
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_385
timestamp 1704896540
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_391
timestamp 1704896540
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_393
timestamp 1704896540
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_405
timestamp 1704896540
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_417
timestamp 1704896540
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1704896540
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1704896540
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1704896540
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1704896540
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp 1704896540
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_53
timestamp 1704896540
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_65
timestamp 1704896540
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_77
timestamp 1704896540
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 1704896540
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_85
timestamp 1704896540
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_97
timestamp 1704896540
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_109
timestamp 1704896540
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_121
timestamp 1704896540
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_133
timestamp 1704896540
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 1704896540
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_141
timestamp 1704896540
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_153
timestamp 1704896540
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_165
timestamp 1704896540
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_177
timestamp 1704896540
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_189
timestamp 1704896540
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 1704896540
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_197
timestamp 1704896540
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_209
timestamp 1704896540
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_221
timestamp 1704896540
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_233
timestamp 1704896540
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_245
timestamp 1704896540
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_251
timestamp 1704896540
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_253
timestamp 1704896540
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_265
timestamp 1704896540
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_277
timestamp 1704896540
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_289
timestamp 1704896540
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_301
timestamp 1704896540
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_307
timestamp 1704896540
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_309
timestamp 1704896540
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_321
timestamp 1704896540
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_333
timestamp 1704896540
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_345
timestamp 1704896540
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_357
timestamp 1704896540
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_363
timestamp 1704896540
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_365
timestamp 1704896540
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_377
timestamp 1704896540
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_389
timestamp 1704896540
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_401
timestamp 1704896540
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_413
timestamp 1704896540
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_419
timestamp 1704896540
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_421
timestamp 1704896540
transform 1 0 39836 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1704896540
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 1704896540
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_27
timestamp 1704896540
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_39
timestamp 1704896540
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_51
timestamp 1704896540
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 1704896540
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 1704896540
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_69
timestamp 1704896540
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_81
timestamp 1704896540
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_93
timestamp 1704896540
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_105
timestamp 1704896540
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 1704896540
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_113
timestamp 1704896540
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_125
timestamp 1704896540
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_137
timestamp 1704896540
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_149
timestamp 1704896540
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_161
timestamp 1704896540
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 1704896540
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_169
timestamp 1704896540
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_181
timestamp 1704896540
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_193
timestamp 1704896540
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_205
timestamp 1704896540
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_217
timestamp 1704896540
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_223
timestamp 1704896540
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_225
timestamp 1704896540
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_237
timestamp 1704896540
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_249
timestamp 1704896540
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_261
timestamp 1704896540
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_273
timestamp 1704896540
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_279
timestamp 1704896540
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_281
timestamp 1704896540
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_293
timestamp 1704896540
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_305
timestamp 1704896540
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_317
timestamp 1704896540
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_329
timestamp 1704896540
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_335
timestamp 1704896540
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_337
timestamp 1704896540
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_349
timestamp 1704896540
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_361
timestamp 1704896540
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_373
timestamp 1704896540
transform 1 0 35420 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_379
timestamp 1704896540
transform 1 0 35972 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_382
timestamp 1704896540
transform 1 0 36248 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_390
timestamp 1704896540
transform 1 0 36984 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_393
timestamp 1704896540
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_405
timestamp 1704896540
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_417
timestamp 1704896540
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1704896540
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_15
timestamp 1704896540
transform 1 0 2484 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_23
timestamp 1704896540
transform 1 0 3220 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1704896540
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_41
timestamp 1704896540
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_53
timestamp 1704896540
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_65
timestamp 1704896540
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_77
timestamp 1704896540
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1704896540
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_85
timestamp 1704896540
transform 1 0 8924 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_90
timestamp 1704896540
transform 1 0 9384 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_115
timestamp 1704896540
transform 1 0 11684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_127
timestamp 1704896540
transform 1 0 12788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 1704896540
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 1704896540
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_153
timestamp 1704896540
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_165
timestamp 1704896540
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_177
timestamp 1704896540
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_189
timestamp 1704896540
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_195
timestamp 1704896540
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_197
timestamp 1704896540
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_209
timestamp 1704896540
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_221
timestamp 1704896540
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_233
timestamp 1704896540
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_245
timestamp 1704896540
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 1704896540
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_253
timestamp 1704896540
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_265
timestamp 1704896540
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_277
timestamp 1704896540
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_289
timestamp 1704896540
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_301
timestamp 1704896540
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_307
timestamp 1704896540
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_309
timestamp 1704896540
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_321
timestamp 1704896540
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_333
timestamp 1704896540
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_345
timestamp 1704896540
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_357
timestamp 1704896540
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_363
timestamp 1704896540
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_365
timestamp 1704896540
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_377
timestamp 1704896540
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_389
timestamp 1704896540
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_401
timestamp 1704896540
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_413
timestamp 1704896540
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_419
timestamp 1704896540
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_421
timestamp 1704896540
transform 1 0 39836 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1704896540
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 1704896540
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_27
timestamp 1704896540
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_39
timestamp 1704896540
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_51
timestamp 1704896540
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 1704896540
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_57
timestamp 1704896540
transform 1 0 6348 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_83
timestamp 1704896540
transform 1 0 8740 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_95
timestamp 1704896540
transform 1 0 9844 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_107
timestamp 1704896540
transform 1 0 10948 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 1704896540
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_113
timestamp 1704896540
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_125
timestamp 1704896540
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_137
timestamp 1704896540
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_149
timestamp 1704896540
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_161
timestamp 1704896540
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 1704896540
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_169
timestamp 1704896540
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_181
timestamp 1704896540
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_193
timestamp 1704896540
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_205
timestamp 1704896540
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_217
timestamp 1704896540
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_223
timestamp 1704896540
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_225
timestamp 1704896540
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_237
timestamp 1704896540
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_249
timestamp 1704896540
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_261
timestamp 1704896540
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_273
timestamp 1704896540
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_279
timestamp 1704896540
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_281
timestamp 1704896540
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_293
timestamp 1704896540
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_305
timestamp 1704896540
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_317
timestamp 1704896540
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_329
timestamp 1704896540
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_335
timestamp 1704896540
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_337
timestamp 1704896540
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_349
timestamp 1704896540
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_361
timestamp 1704896540
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_373
timestamp 1704896540
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_385
timestamp 1704896540
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_391
timestamp 1704896540
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_393
timestamp 1704896540
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_405
timestamp 1704896540
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_417
timestamp 1704896540
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1704896540
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 1704896540
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1704896540
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 1704896540
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_41
timestamp 1704896540
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_53
timestamp 1704896540
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_65
timestamp 1704896540
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_77
timestamp 1704896540
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 1704896540
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_85
timestamp 1704896540
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_97
timestamp 1704896540
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_109
timestamp 1704896540
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_121
timestamp 1704896540
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_133
timestamp 1704896540
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 1704896540
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_141
timestamp 1704896540
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_153
timestamp 1704896540
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_165
timestamp 1704896540
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_177
timestamp 1704896540
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_189
timestamp 1704896540
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 1704896540
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_220
timestamp 1704896540
transform 1 0 21344 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_224
timestamp 1704896540
transform 1 0 21712 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_228
timestamp 1704896540
transform 1 0 22080 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_240
timestamp 1704896540
transform 1 0 23184 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_253
timestamp 1704896540
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_265
timestamp 1704896540
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_277
timestamp 1704896540
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_289
timestamp 1704896540
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_301
timestamp 1704896540
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_307
timestamp 1704896540
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_309
timestamp 1704896540
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_321
timestamp 1704896540
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_333
timestamp 1704896540
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_345
timestamp 1704896540
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_357
timestamp 1704896540
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_363
timestamp 1704896540
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_365
timestamp 1704896540
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_377
timestamp 1704896540
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_389
timestamp 1704896540
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_401
timestamp 1704896540
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_413
timestamp 1704896540
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_419
timestamp 1704896540
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_421
timestamp 1704896540
transform 1 0 39836 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1704896540
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_15
timestamp 1704896540
transform 1 0 2484 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_18
timestamp 1704896540
transform 1 0 2760 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_43
timestamp 1704896540
transform 1 0 5060 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_47
timestamp 1704896540
transform 1 0 5428 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 1704896540
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 1704896540
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_69
timestamp 1704896540
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_81
timestamp 1704896540
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_93
timestamp 1704896540
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_105
timestamp 1704896540
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_111
timestamp 1704896540
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_113
timestamp 1704896540
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_125
timestamp 1704896540
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_137
timestamp 1704896540
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_149
timestamp 1704896540
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_161
timestamp 1704896540
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_167
timestamp 1704896540
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_169
timestamp 1704896540
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_181
timestamp 1704896540
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_193
timestamp 1704896540
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_205
timestamp 1704896540
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_217
timestamp 1704896540
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_223
timestamp 1704896540
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_225
timestamp 1704896540
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_237
timestamp 1704896540
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_249
timestamp 1704896540
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_261
timestamp 1704896540
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_273
timestamp 1704896540
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_279
timestamp 1704896540
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_281
timestamp 1704896540
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_293
timestamp 1704896540
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_305
timestamp 1704896540
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_317
timestamp 1704896540
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_329
timestamp 1704896540
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_335
timestamp 1704896540
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_337
timestamp 1704896540
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_349
timestamp 1704896540
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_361
timestamp 1704896540
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_373
timestamp 1704896540
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_385
timestamp 1704896540
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_391
timestamp 1704896540
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_393
timestamp 1704896540
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_405
timestamp 1704896540
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_417
timestamp 1704896540
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 1704896540
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_15
timestamp 1704896540
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1704896540
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_29
timestamp 1704896540
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_41
timestamp 1704896540
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_53
timestamp 1704896540
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_65
timestamp 1704896540
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_77
timestamp 1704896540
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_83
timestamp 1704896540
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_85
timestamp 1704896540
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_97
timestamp 1704896540
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_109
timestamp 1704896540
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_121
timestamp 1704896540
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_133
timestamp 1704896540
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_139
timestamp 1704896540
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_141
timestamp 1704896540
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_153
timestamp 1704896540
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_165
timestamp 1704896540
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_177
timestamp 1704896540
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_189
timestamp 1704896540
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_195
timestamp 1704896540
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_197
timestamp 1704896540
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_209
timestamp 1704896540
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_221
timestamp 1704896540
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_233
timestamp 1704896540
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_245
timestamp 1704896540
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_251
timestamp 1704896540
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_253
timestamp 1704896540
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_265
timestamp 1704896540
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_277
timestamp 1704896540
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_289
timestamp 1704896540
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_301
timestamp 1704896540
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_307
timestamp 1704896540
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_309
timestamp 1704896540
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_321
timestamp 1704896540
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_333
timestamp 1704896540
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_345
timestamp 1704896540
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_357
timestamp 1704896540
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_363
timestamp 1704896540
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_365
timestamp 1704896540
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_377
timestamp 1704896540
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_389
timestamp 1704896540
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_401
timestamp 1704896540
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_413
timestamp 1704896540
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_419
timestamp 1704896540
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_421
timestamp 1704896540
transform 1 0 39836 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 1704896540
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_15
timestamp 1704896540
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_27
timestamp 1704896540
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_39
timestamp 1704896540
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_51
timestamp 1704896540
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 1704896540
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_57
timestamp 1704896540
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_69
timestamp 1704896540
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_81
timestamp 1704896540
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_93
timestamp 1704896540
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_105
timestamp 1704896540
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_111
timestamp 1704896540
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_113
timestamp 1704896540
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_125
timestamp 1704896540
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_137
timestamp 1704896540
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_149
timestamp 1704896540
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_161
timestamp 1704896540
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_167
timestamp 1704896540
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_169
timestamp 1704896540
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_181
timestamp 1704896540
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_193
timestamp 1704896540
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_205
timestamp 1704896540
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_217
timestamp 1704896540
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_223
timestamp 1704896540
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_225
timestamp 1704896540
transform 1 0 21804 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_256
timestamp 1704896540
transform 1 0 24656 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_268
timestamp 1704896540
transform 1 0 25760 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_281
timestamp 1704896540
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_293
timestamp 1704896540
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_305
timestamp 1704896540
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_317
timestamp 1704896540
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_329
timestamp 1704896540
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_335
timestamp 1704896540
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_337
timestamp 1704896540
transform 1 0 32108 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_357
timestamp 1704896540
transform 1 0 33948 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_369
timestamp 1704896540
transform 1 0 35052 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_381
timestamp 1704896540
transform 1 0 36156 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_389
timestamp 1704896540
transform 1 0 36892 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_393
timestamp 1704896540
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_405
timestamp 1704896540
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_417
timestamp 1704896540
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 1704896540
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_15
timestamp 1704896540
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1704896540
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_29
timestamp 1704896540
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_41
timestamp 1704896540
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_53
timestamp 1704896540
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_65
timestamp 1704896540
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_77
timestamp 1704896540
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_83
timestamp 1704896540
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_85
timestamp 1704896540
transform 1 0 8924 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_109
timestamp 1704896540
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_121
timestamp 1704896540
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_133
timestamp 1704896540
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_139
timestamp 1704896540
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_141
timestamp 1704896540
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_153
timestamp 1704896540
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_165
timestamp 1704896540
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_177
timestamp 1704896540
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_189
timestamp 1704896540
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_195
timestamp 1704896540
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_197
timestamp 1704896540
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_209
timestamp 1704896540
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_221
timestamp 1704896540
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_233
timestamp 1704896540
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_245
timestamp 1704896540
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_251
timestamp 1704896540
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_253
timestamp 1704896540
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_261
timestamp 1704896540
transform 1 0 25116 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_273
timestamp 1704896540
transform 1 0 26220 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_285
timestamp 1704896540
transform 1 0 27324 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_297
timestamp 1704896540
transform 1 0 28428 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_305
timestamp 1704896540
transform 1 0 29164 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_309
timestamp 1704896540
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_321
timestamp 1704896540
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_333
timestamp 1704896540
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_345
timestamp 1704896540
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_357
timestamp 1704896540
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_363
timestamp 1704896540
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_365
timestamp 1704896540
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_377
timestamp 1704896540
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_389
timestamp 1704896540
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_401
timestamp 1704896540
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_413
timestamp 1704896540
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_419
timestamp 1704896540
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_421
timestamp 1704896540
transform 1 0 39836 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 1704896540
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_15
timestamp 1704896540
transform 1 0 2484 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_27
timestamp 1704896540
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_39
timestamp 1704896540
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_51
timestamp 1704896540
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 1704896540
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_66
timestamp 1704896540
transform 1 0 7176 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_70
timestamp 1704896540
transform 1 0 7544 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_82
timestamp 1704896540
transform 1 0 8648 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_94
timestamp 1704896540
transform 1 0 9752 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_106
timestamp 1704896540
transform 1 0 10856 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_113
timestamp 1704896540
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_125
timestamp 1704896540
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_137
timestamp 1704896540
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_149
timestamp 1704896540
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_161
timestamp 1704896540
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_167
timestamp 1704896540
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_169
timestamp 1704896540
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_181
timestamp 1704896540
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_193
timestamp 1704896540
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_205
timestamp 1704896540
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_217
timestamp 1704896540
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_223
timestamp 1704896540
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_225
timestamp 1704896540
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_237
timestamp 1704896540
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_249
timestamp 1704896540
transform 1 0 24012 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_275
timestamp 1704896540
transform 1 0 26404 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_279
timestamp 1704896540
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_281
timestamp 1704896540
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_293
timestamp 1704896540
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_305
timestamp 1704896540
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_317
timestamp 1704896540
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_329
timestamp 1704896540
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_335
timestamp 1704896540
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_337
timestamp 1704896540
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_349
timestamp 1704896540
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_361
timestamp 1704896540
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_373
timestamp 1704896540
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_385
timestamp 1704896540
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_391
timestamp 1704896540
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_393
timestamp 1704896540
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_405
timestamp 1704896540
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_417
timestamp 1704896540
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 1704896540
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_15
timestamp 1704896540
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1704896540
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_29
timestamp 1704896540
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_41
timestamp 1704896540
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_53
timestamp 1704896540
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_65
timestamp 1704896540
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_77
timestamp 1704896540
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_83
timestamp 1704896540
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_85
timestamp 1704896540
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_97
timestamp 1704896540
transform 1 0 10028 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_102
timestamp 1704896540
transform 1 0 10488 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_114
timestamp 1704896540
transform 1 0 11592 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_126
timestamp 1704896540
transform 1 0 12696 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_138
timestamp 1704896540
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_141
timestamp 1704896540
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_153
timestamp 1704896540
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_165
timestamp 1704896540
transform 1 0 16284 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_170
timestamp 1704896540
transform 1 0 16744 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_182
timestamp 1704896540
transform 1 0 17848 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_194
timestamp 1704896540
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_197
timestamp 1704896540
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_209
timestamp 1704896540
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_221
timestamp 1704896540
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_233
timestamp 1704896540
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_245
timestamp 1704896540
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_251
timestamp 1704896540
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_253
timestamp 1704896540
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_265
timestamp 1704896540
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_277
timestamp 1704896540
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_289
timestamp 1704896540
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_301
timestamp 1704896540
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_307
timestamp 1704896540
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_309
timestamp 1704896540
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_321
timestamp 1704896540
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_333
timestamp 1704896540
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_345
timestamp 1704896540
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_357
timestamp 1704896540
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_363
timestamp 1704896540
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_365
timestamp 1704896540
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_377
timestamp 1704896540
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_389
timestamp 1704896540
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_401
timestamp 1704896540
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_413
timestamp 1704896540
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_419
timestamp 1704896540
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_421
timestamp 1704896540
transform 1 0 39836 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 1704896540
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_15
timestamp 1704896540
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_27
timestamp 1704896540
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_39
timestamp 1704896540
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_51
timestamp 1704896540
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_55
timestamp 1704896540
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_57
timestamp 1704896540
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_69
timestamp 1704896540
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_81
timestamp 1704896540
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_93
timestamp 1704896540
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_105
timestamp 1704896540
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_111
timestamp 1704896540
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_113
timestamp 1704896540
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_125
timestamp 1704896540
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_137
timestamp 1704896540
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_149
timestamp 1704896540
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_161
timestamp 1704896540
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_167
timestamp 1704896540
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_169
timestamp 1704896540
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_181
timestamp 1704896540
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_193
timestamp 1704896540
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_205
timestamp 1704896540
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_217
timestamp 1704896540
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_223
timestamp 1704896540
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_228
timestamp 1704896540
transform 1 0 22080 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_240
timestamp 1704896540
transform 1 0 23184 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_252
timestamp 1704896540
transform 1 0 24288 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_264
timestamp 1704896540
transform 1 0 25392 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_276
timestamp 1704896540
transform 1 0 26496 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_281
timestamp 1704896540
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_293
timestamp 1704896540
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_305
timestamp 1704896540
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_317
timestamp 1704896540
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_329
timestamp 1704896540
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_335
timestamp 1704896540
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_337
timestamp 1704896540
transform 1 0 32108 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_343
timestamp 1704896540
transform 1 0 32660 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_346
timestamp 1704896540
transform 1 0 32936 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_354
timestamp 1704896540
transform 1 0 33672 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_358
timestamp 1704896540
transform 1 0 34040 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_370
timestamp 1704896540
transform 1 0 35144 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_382
timestamp 1704896540
transform 1 0 36248 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_390
timestamp 1704896540
transform 1 0 36984 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_393
timestamp 1704896540
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_405
timestamp 1704896540
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_417
timestamp 1704896540
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_3
timestamp 1704896540
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_15
timestamp 1704896540
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1704896540
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_29
timestamp 1704896540
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_41
timestamp 1704896540
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_53
timestamp 1704896540
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_65
timestamp 1704896540
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_77
timestamp 1704896540
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_83
timestamp 1704896540
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_85
timestamp 1704896540
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_97
timestamp 1704896540
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_109
timestamp 1704896540
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_121
timestamp 1704896540
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_133
timestamp 1704896540
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_139
timestamp 1704896540
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_141
timestamp 1704896540
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_153
timestamp 1704896540
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_165
timestamp 1704896540
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_177
timestamp 1704896540
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_189
timestamp 1704896540
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_195
timestamp 1704896540
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_197
timestamp 1704896540
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_209
timestamp 1704896540
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_221
timestamp 1704896540
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_233
timestamp 1704896540
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_245
timestamp 1704896540
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_251
timestamp 1704896540
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_253
timestamp 1704896540
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_265
timestamp 1704896540
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_277
timestamp 1704896540
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_289
timestamp 1704896540
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_301
timestamp 1704896540
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_307
timestamp 1704896540
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_309
timestamp 1704896540
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_321
timestamp 1704896540
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_333
timestamp 1704896540
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_345
timestamp 1704896540
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_357
timestamp 1704896540
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_363
timestamp 1704896540
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_365
timestamp 1704896540
transform 1 0 34684 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_380
timestamp 1704896540
transform 1 0 36064 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_392
timestamp 1704896540
transform 1 0 37168 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_404
timestamp 1704896540
transform 1 0 38272 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_416
timestamp 1704896540
transform 1 0 39376 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_421
timestamp 1704896540
transform 1 0 39836 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_3
timestamp 1704896540
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_15
timestamp 1704896540
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_27
timestamp 1704896540
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_39
timestamp 1704896540
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_51
timestamp 1704896540
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_55
timestamp 1704896540
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_57
timestamp 1704896540
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_69
timestamp 1704896540
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_81
timestamp 1704896540
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_93
timestamp 1704896540
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_105
timestamp 1704896540
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_111
timestamp 1704896540
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_113
timestamp 1704896540
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_125
timestamp 1704896540
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_137
timestamp 1704896540
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_149
timestamp 1704896540
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_161
timestamp 1704896540
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_167
timestamp 1704896540
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_169
timestamp 1704896540
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_181
timestamp 1704896540
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_193
timestamp 1704896540
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_205
timestamp 1704896540
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_217
timestamp 1704896540
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_223
timestamp 1704896540
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_225
timestamp 1704896540
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_237
timestamp 1704896540
transform 1 0 22908 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_266
timestamp 1704896540
transform 1 0 25576 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_278
timestamp 1704896540
transform 1 0 26680 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_281
timestamp 1704896540
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_293
timestamp 1704896540
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_305
timestamp 1704896540
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_317
timestamp 1704896540
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_329
timestamp 1704896540
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_335
timestamp 1704896540
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_337
timestamp 1704896540
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_349
timestamp 1704896540
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_361
timestamp 1704896540
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_373
timestamp 1704896540
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_385
timestamp 1704896540
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_391
timestamp 1704896540
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_393
timestamp 1704896540
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_405
timestamp 1704896540
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_417
timestamp 1704896540
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_3
timestamp 1704896540
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_15
timestamp 1704896540
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 1704896540
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_29
timestamp 1704896540
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_41
timestamp 1704896540
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_53
timestamp 1704896540
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_65
timestamp 1704896540
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_77
timestamp 1704896540
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_83
timestamp 1704896540
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_85
timestamp 1704896540
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_97
timestamp 1704896540
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_109
timestamp 1704896540
transform 1 0 11132 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_115
timestamp 1704896540
transform 1 0 11684 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_141
timestamp 1704896540
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_153
timestamp 1704896540
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_165
timestamp 1704896540
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_177
timestamp 1704896540
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_189
timestamp 1704896540
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_195
timestamp 1704896540
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_197
timestamp 1704896540
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_209
timestamp 1704896540
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_221
timestamp 1704896540
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_233
timestamp 1704896540
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_245
timestamp 1704896540
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_251
timestamp 1704896540
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_253
timestamp 1704896540
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_265
timestamp 1704896540
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_277
timestamp 1704896540
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_289
timestamp 1704896540
transform 1 0 27692 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_297
timestamp 1704896540
transform 1 0 28428 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_305
timestamp 1704896540
transform 1 0 29164 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_309
timestamp 1704896540
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_321
timestamp 1704896540
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_333
timestamp 1704896540
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_345
timestamp 1704896540
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_357
timestamp 1704896540
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_363
timestamp 1704896540
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_365
timestamp 1704896540
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_377
timestamp 1704896540
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_389
timestamp 1704896540
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_401
timestamp 1704896540
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_413
timestamp 1704896540
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_419
timestamp 1704896540
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_421
timestamp 1704896540
transform 1 0 39836 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_3
timestamp 1704896540
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_15
timestamp 1704896540
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_27
timestamp 1704896540
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_39
timestamp 1704896540
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_51
timestamp 1704896540
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 1704896540
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_57
timestamp 1704896540
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_69
timestamp 1704896540
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_81
timestamp 1704896540
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_93
timestamp 1704896540
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_105
timestamp 1704896540
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_111
timestamp 1704896540
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_113
timestamp 1704896540
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_125
timestamp 1704896540
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_137
timestamp 1704896540
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_149
timestamp 1704896540
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_161
timestamp 1704896540
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_167
timestamp 1704896540
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_169
timestamp 1704896540
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_181
timestamp 1704896540
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_193
timestamp 1704896540
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_205
timestamp 1704896540
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_217
timestamp 1704896540
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_223
timestamp 1704896540
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_225
timestamp 1704896540
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_237
timestamp 1704896540
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_249
timestamp 1704896540
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_261
timestamp 1704896540
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_273
timestamp 1704896540
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_279
timestamp 1704896540
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_281
timestamp 1704896540
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_293
timestamp 1704896540
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_305
timestamp 1704896540
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_317
timestamp 1704896540
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_329
timestamp 1704896540
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_335
timestamp 1704896540
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_345
timestamp 1704896540
transform 1 0 32844 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_357
timestamp 1704896540
transform 1 0 33948 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_369
timestamp 1704896540
transform 1 0 35052 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_381
timestamp 1704896540
transform 1 0 36156 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_389
timestamp 1704896540
transform 1 0 36892 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_393
timestamp 1704896540
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_405
timestamp 1704896540
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_417
timestamp 1704896540
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_3
timestamp 1704896540
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_15
timestamp 1704896540
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 1704896540
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_29
timestamp 1704896540
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_41
timestamp 1704896540
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_53
timestamp 1704896540
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_65
timestamp 1704896540
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_77
timestamp 1704896540
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 1704896540
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_85
timestamp 1704896540
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_97
timestamp 1704896540
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_109
timestamp 1704896540
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_121
timestamp 1704896540
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_133
timestamp 1704896540
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_139
timestamp 1704896540
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_141
timestamp 1704896540
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_153
timestamp 1704896540
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_165
timestamp 1704896540
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_177
timestamp 1704896540
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_189
timestamp 1704896540
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_195
timestamp 1704896540
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_197
timestamp 1704896540
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_209
timestamp 1704896540
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_221
timestamp 1704896540
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_233
timestamp 1704896540
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_245
timestamp 1704896540
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_251
timestamp 1704896540
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_253
timestamp 1704896540
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_265
timestamp 1704896540
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_277
timestamp 1704896540
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_289
timestamp 1704896540
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_301
timestamp 1704896540
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_307
timestamp 1704896540
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_309
timestamp 1704896540
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_321
timestamp 1704896540
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_333
timestamp 1704896540
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_345
timestamp 1704896540
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_357
timestamp 1704896540
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_363
timestamp 1704896540
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_365
timestamp 1704896540
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_377
timestamp 1704896540
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_389
timestamp 1704896540
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_401
timestamp 1704896540
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_413
timestamp 1704896540
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_419
timestamp 1704896540
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_421
timestamp 1704896540
transform 1 0 39836 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 1704896540
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_15
timestamp 1704896540
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_27
timestamp 1704896540
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_39
timestamp 1704896540
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_51
timestamp 1704896540
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 1704896540
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_57
timestamp 1704896540
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_69
timestamp 1704896540
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_81
timestamp 1704896540
transform 1 0 8556 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_90
timestamp 1704896540
transform 1 0 9384 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_102
timestamp 1704896540
transform 1 0 10488 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_110
timestamp 1704896540
transform 1 0 11224 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_113
timestamp 1704896540
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_125
timestamp 1704896540
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_137
timestamp 1704896540
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_149
timestamp 1704896540
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_161
timestamp 1704896540
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_167
timestamp 1704896540
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_169
timestamp 1704896540
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_181
timestamp 1704896540
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_193
timestamp 1704896540
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_205
timestamp 1704896540
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_217
timestamp 1704896540
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_223
timestamp 1704896540
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_225
timestamp 1704896540
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_237
timestamp 1704896540
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_249
timestamp 1704896540
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_261
timestamp 1704896540
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_273
timestamp 1704896540
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_279
timestamp 1704896540
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_281
timestamp 1704896540
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_293
timestamp 1704896540
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_305
timestamp 1704896540
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_317
timestamp 1704896540
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_329
timestamp 1704896540
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_335
timestamp 1704896540
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_337
timestamp 1704896540
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_349
timestamp 1704896540
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_361
timestamp 1704896540
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_373
timestamp 1704896540
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_385
timestamp 1704896540
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_391
timestamp 1704896540
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_393
timestamp 1704896540
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_405
timestamp 1704896540
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_417
timestamp 1704896540
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_3
timestamp 1704896540
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_15
timestamp 1704896540
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 1704896540
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_29
timestamp 1704896540
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_41
timestamp 1704896540
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_53
timestamp 1704896540
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_65
timestamp 1704896540
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_77
timestamp 1704896540
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_83
timestamp 1704896540
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_85
timestamp 1704896540
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_97
timestamp 1704896540
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_109
timestamp 1704896540
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_121
timestamp 1704896540
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_133
timestamp 1704896540
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_139
timestamp 1704896540
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_141
timestamp 1704896540
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_153
timestamp 1704896540
transform 1 0 15180 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_158
timestamp 1704896540
transform 1 0 15640 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_183
timestamp 1704896540
transform 1 0 17940 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_195
timestamp 1704896540
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_197
timestamp 1704896540
transform 1 0 19228 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_213
timestamp 1704896540
transform 1 0 20700 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_225
timestamp 1704896540
transform 1 0 21804 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_237
timestamp 1704896540
transform 1 0 22908 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_249
timestamp 1704896540
transform 1 0 24012 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_253
timestamp 1704896540
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_265
timestamp 1704896540
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_277
timestamp 1704896540
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_289
timestamp 1704896540
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_301
timestamp 1704896540
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_307
timestamp 1704896540
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_309
timestamp 1704896540
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_321
timestamp 1704896540
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_333
timestamp 1704896540
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_345
timestamp 1704896540
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_357
timestamp 1704896540
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_363
timestamp 1704896540
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_365
timestamp 1704896540
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_377
timestamp 1704896540
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_389
timestamp 1704896540
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_401
timestamp 1704896540
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_413
timestamp 1704896540
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_419
timestamp 1704896540
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_421
timestamp 1704896540
transform 1 0 39836 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_3
timestamp 1704896540
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_15
timestamp 1704896540
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_27
timestamp 1704896540
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_39
timestamp 1704896540
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_51
timestamp 1704896540
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_55
timestamp 1704896540
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_57
timestamp 1704896540
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_69
timestamp 1704896540
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_81
timestamp 1704896540
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_93
timestamp 1704896540
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_105
timestamp 1704896540
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_111
timestamp 1704896540
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_113
timestamp 1704896540
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_125
timestamp 1704896540
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_137
timestamp 1704896540
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_149
timestamp 1704896540
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_161
timestamp 1704896540
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_167
timestamp 1704896540
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_169
timestamp 1704896540
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_181
timestamp 1704896540
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_193
timestamp 1704896540
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_205
timestamp 1704896540
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_217
timestamp 1704896540
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_223
timestamp 1704896540
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_228
timestamp 1704896540
transform 1 0 22080 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_232
timestamp 1704896540
transform 1 0 22448 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_244
timestamp 1704896540
transform 1 0 23552 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_256
timestamp 1704896540
transform 1 0 24656 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_268
timestamp 1704896540
transform 1 0 25760 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_281
timestamp 1704896540
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_293
timestamp 1704896540
transform 1 0 28060 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_303
timestamp 1704896540
transform 1 0 28980 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_310
timestamp 1704896540
transform 1 0 29624 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_314
timestamp 1704896540
transform 1 0 29992 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_326
timestamp 1704896540
transform 1 0 31096 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_334
timestamp 1704896540
transform 1 0 31832 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_337
timestamp 1704896540
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_349
timestamp 1704896540
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_361
timestamp 1704896540
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_373
timestamp 1704896540
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_385
timestamp 1704896540
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_391
timestamp 1704896540
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_393
timestamp 1704896540
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_405
timestamp 1704896540
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_417
timestamp 1704896540
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_3
timestamp 1704896540
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_15
timestamp 1704896540
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_27
timestamp 1704896540
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_29
timestamp 1704896540
transform 1 0 3772 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_37
timestamp 1704896540
transform 1 0 4508 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_41
timestamp 1704896540
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_53
timestamp 1704896540
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_65
timestamp 1704896540
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_77
timestamp 1704896540
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_83
timestamp 1704896540
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_85
timestamp 1704896540
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_97
timestamp 1704896540
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_109
timestamp 1704896540
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_121
timestamp 1704896540
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_133
timestamp 1704896540
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_139
timestamp 1704896540
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_141
timestamp 1704896540
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_153
timestamp 1704896540
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_165
timestamp 1704896540
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_177
timestamp 1704896540
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_189
timestamp 1704896540
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_195
timestamp 1704896540
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_204
timestamp 1704896540
transform 1 0 19872 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_216
timestamp 1704896540
transform 1 0 20976 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_228
timestamp 1704896540
transform 1 0 22080 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_240
timestamp 1704896540
transform 1 0 23184 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_253
timestamp 1704896540
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_265
timestamp 1704896540
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_277
timestamp 1704896540
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_289
timestamp 1704896540
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_301
timestamp 1704896540
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_307
timestamp 1704896540
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_322
timestamp 1704896540
transform 1 0 30728 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_334
timestamp 1704896540
transform 1 0 31832 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_346
timestamp 1704896540
transform 1 0 32936 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_358
timestamp 1704896540
transform 1 0 34040 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_365
timestamp 1704896540
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_377
timestamp 1704896540
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_389
timestamp 1704896540
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_401
timestamp 1704896540
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_413
timestamp 1704896540
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_419
timestamp 1704896540
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_421
timestamp 1704896540
transform 1 0 39836 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_3
timestamp 1704896540
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_15
timestamp 1704896540
transform 1 0 2484 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_23
timestamp 1704896540
transform 1 0 3220 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_28
timestamp 1704896540
transform 1 0 3680 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_53
timestamp 1704896540
transform 1 0 5980 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_68
timestamp 1704896540
transform 1 0 7360 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_80
timestamp 1704896540
transform 1 0 8464 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_92
timestamp 1704896540
transform 1 0 9568 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_104
timestamp 1704896540
transform 1 0 10672 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_113
timestamp 1704896540
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_125
timestamp 1704896540
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_137
timestamp 1704896540
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_149
timestamp 1704896540
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_161
timestamp 1704896540
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_167
timestamp 1704896540
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_169
timestamp 1704896540
transform 1 0 16652 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_178
timestamp 1704896540
transform 1 0 17480 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_209
timestamp 1704896540
transform 1 0 20332 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_221
timestamp 1704896540
transform 1 0 21436 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_225
timestamp 1704896540
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_237
timestamp 1704896540
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_249
timestamp 1704896540
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_261
timestamp 1704896540
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_273
timestamp 1704896540
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_279
timestamp 1704896540
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_281
timestamp 1704896540
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_293
timestamp 1704896540
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_305
timestamp 1704896540
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_317
timestamp 1704896540
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_329
timestamp 1704896540
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_335
timestamp 1704896540
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_337
timestamp 1704896540
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_349
timestamp 1704896540
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_361
timestamp 1704896540
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_373
timestamp 1704896540
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_385
timestamp 1704896540
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_391
timestamp 1704896540
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_393
timestamp 1704896540
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_405
timestamp 1704896540
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_3
timestamp 1704896540
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_15
timestamp 1704896540
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 1704896540
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_29
timestamp 1704896540
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_41
timestamp 1704896540
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_79
timestamp 1704896540
transform 1 0 8372 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_83
timestamp 1704896540
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_85
timestamp 1704896540
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_97
timestamp 1704896540
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_109
timestamp 1704896540
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_121
timestamp 1704896540
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_133
timestamp 1704896540
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_139
timestamp 1704896540
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_153
timestamp 1704896540
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_165
timestamp 1704896540
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_177
timestamp 1704896540
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_189
timestamp 1704896540
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_195
timestamp 1704896540
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_197
timestamp 1704896540
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_209
timestamp 1704896540
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_221
timestamp 1704896540
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_233
timestamp 1704896540
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_245
timestamp 1704896540
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_251
timestamp 1704896540
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_253
timestamp 1704896540
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_265
timestamp 1704896540
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_277
timestamp 1704896540
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_289
timestamp 1704896540
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_301
timestamp 1704896540
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_307
timestamp 1704896540
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_309
timestamp 1704896540
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_321
timestamp 1704896540
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_333
timestamp 1704896540
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_345
timestamp 1704896540
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_357
timestamp 1704896540
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_363
timestamp 1704896540
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_365
timestamp 1704896540
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_377
timestamp 1704896540
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_389
timestamp 1704896540
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_401
timestamp 1704896540
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_413
timestamp 1704896540
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_419
timestamp 1704896540
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_421
timestamp 1704896540
transform 1 0 39836 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_3
timestamp 1704896540
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_15
timestamp 1704896540
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_27
timestamp 1704896540
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_39
timestamp 1704896540
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_51
timestamp 1704896540
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_55
timestamp 1704896540
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_57
timestamp 1704896540
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_69
timestamp 1704896540
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_81
timestamp 1704896540
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_93
timestamp 1704896540
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_105
timestamp 1704896540
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_111
timestamp 1704896540
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_113
timestamp 1704896540
transform 1 0 11500 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_120
timestamp 1704896540
transform 1 0 12144 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_132
timestamp 1704896540
transform 1 0 13248 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_144
timestamp 1704896540
transform 1 0 14352 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_156
timestamp 1704896540
transform 1 0 15456 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_169
timestamp 1704896540
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_181
timestamp 1704896540
transform 1 0 17756 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_192
timestamp 1704896540
transform 1 0 18768 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_204
timestamp 1704896540
transform 1 0 19872 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_216
timestamp 1704896540
transform 1 0 20976 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_225
timestamp 1704896540
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_237
timestamp 1704896540
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_249
timestamp 1704896540
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_261
timestamp 1704896540
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_273
timestamp 1704896540
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_279
timestamp 1704896540
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_281
timestamp 1704896540
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_293
timestamp 1704896540
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_305
timestamp 1704896540
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_317
timestamp 1704896540
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_329
timestamp 1704896540
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_335
timestamp 1704896540
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_337
timestamp 1704896540
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_349
timestamp 1704896540
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_361
timestamp 1704896540
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_373
timestamp 1704896540
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_385
timestamp 1704896540
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_391
timestamp 1704896540
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_393
timestamp 1704896540
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_405
timestamp 1704896540
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_417
timestamp 1704896540
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_3
timestamp 1704896540
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_15
timestamp 1704896540
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_27
timestamp 1704896540
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_29
timestamp 1704896540
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_41
timestamp 1704896540
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_53
timestamp 1704896540
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_65
timestamp 1704896540
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_77
timestamp 1704896540
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_83
timestamp 1704896540
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_89
timestamp 1704896540
transform 1 0 9292 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_118
timestamp 1704896540
transform 1 0 11960 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_130
timestamp 1704896540
transform 1 0 13064 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_138
timestamp 1704896540
transform 1 0 13800 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_141
timestamp 1704896540
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_153
timestamp 1704896540
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_165
timestamp 1704896540
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_177
timestamp 1704896540
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_189
timestamp 1704896540
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_195
timestamp 1704896540
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_197
timestamp 1704896540
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_209
timestamp 1704896540
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_221
timestamp 1704896540
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_233
timestamp 1704896540
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_245
timestamp 1704896540
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_251
timestamp 1704896540
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_253
timestamp 1704896540
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_265
timestamp 1704896540
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_277
timestamp 1704896540
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_289
timestamp 1704896540
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_301
timestamp 1704896540
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_307
timestamp 1704896540
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_309
timestamp 1704896540
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_321
timestamp 1704896540
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_333
timestamp 1704896540
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_345
timestamp 1704896540
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_357
timestamp 1704896540
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_363
timestamp 1704896540
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_365
timestamp 1704896540
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_377
timestamp 1704896540
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_389
timestamp 1704896540
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_401
timestamp 1704896540
transform 1 0 37996 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_409
timestamp 1704896540
transform 1 0 38732 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_414
timestamp 1704896540
transform 1 0 39192 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_418
timestamp 1704896540
transform 1 0 39560 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_427
timestamp 1704896540
transform 1 0 40388 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_3
timestamp 1704896540
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_15
timestamp 1704896540
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_27
timestamp 1704896540
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_39
timestamp 1704896540
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_51
timestamp 1704896540
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_55
timestamp 1704896540
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_57
timestamp 1704896540
transform 1 0 6348 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_65
timestamp 1704896540
transform 1 0 7084 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_72
timestamp 1704896540
transform 1 0 7728 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_84
timestamp 1704896540
transform 1 0 8832 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_96
timestamp 1704896540
transform 1 0 9936 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_108
timestamp 1704896540
transform 1 0 11040 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_113
timestamp 1704896540
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_125
timestamp 1704896540
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_137
timestamp 1704896540
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_149
timestamp 1704896540
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_161
timestamp 1704896540
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_167
timestamp 1704896540
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_169
timestamp 1704896540
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_181
timestamp 1704896540
transform 1 0 17756 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_191
timestamp 1704896540
transform 1 0 18676 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_216
timestamp 1704896540
transform 1 0 20976 0 -1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_225
timestamp 1704896540
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_237
timestamp 1704896540
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_249
timestamp 1704896540
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_261
timestamp 1704896540
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_273
timestamp 1704896540
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_279
timestamp 1704896540
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_281
timestamp 1704896540
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_293
timestamp 1704896540
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_305
timestamp 1704896540
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_317
timestamp 1704896540
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_329
timestamp 1704896540
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_335
timestamp 1704896540
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_337
timestamp 1704896540
transform 1 0 32108 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_345
timestamp 1704896540
transform 1 0 32844 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_350
timestamp 1704896540
transform 1 0 33304 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_361
timestamp 1704896540
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_373
timestamp 1704896540
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_385
timestamp 1704896540
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_391
timestamp 1704896540
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_393
timestamp 1704896540
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_405
timestamp 1704896540
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_417
timestamp 1704896540
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_3
timestamp 1704896540
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_15
timestamp 1704896540
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_27
timestamp 1704896540
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_29
timestamp 1704896540
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_41
timestamp 1704896540
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_53
timestamp 1704896540
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_65
timestamp 1704896540
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_77
timestamp 1704896540
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_83
timestamp 1704896540
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_85
timestamp 1704896540
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_97
timestamp 1704896540
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_109
timestamp 1704896540
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_121
timestamp 1704896540
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_133
timestamp 1704896540
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_139
timestamp 1704896540
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_141
timestamp 1704896540
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_153
timestamp 1704896540
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_165
timestamp 1704896540
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_177
timestamp 1704896540
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_189
timestamp 1704896540
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_195
timestamp 1704896540
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_197
timestamp 1704896540
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_209
timestamp 1704896540
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_221
timestamp 1704896540
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_233
timestamp 1704896540
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_245
timestamp 1704896540
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_251
timestamp 1704896540
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_253
timestamp 1704896540
transform 1 0 24380 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_259
timestamp 1704896540
transform 1 0 24932 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_269
timestamp 1704896540
transform 1 0 25852 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_281
timestamp 1704896540
transform 1 0 26956 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_293
timestamp 1704896540
transform 1 0 28060 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_305
timestamp 1704896540
transform 1 0 29164 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_312
timestamp 1704896540
transform 1 0 29808 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_324
timestamp 1704896540
transform 1 0 30912 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_336
timestamp 1704896540
transform 1 0 32016 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_348
timestamp 1704896540
transform 1 0 33120 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_360
timestamp 1704896540
transform 1 0 34224 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_365
timestamp 1704896540
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_377
timestamp 1704896540
transform 1 0 35788 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_390
timestamp 1704896540
transform 1 0 36984 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_402
timestamp 1704896540
transform 1 0 38088 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_414
timestamp 1704896540
transform 1 0 39192 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_418
timestamp 1704896540
transform 1 0 39560 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_427
timestamp 1704896540
transform 1 0 40388 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_3
timestamp 1704896540
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_15
timestamp 1704896540
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_27
timestamp 1704896540
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_39
timestamp 1704896540
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_51
timestamp 1704896540
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_55
timestamp 1704896540
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_57
timestamp 1704896540
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_69
timestamp 1704896540
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_81
timestamp 1704896540
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_93
timestamp 1704896540
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_105
timestamp 1704896540
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_111
timestamp 1704896540
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_113
timestamp 1704896540
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_125
timestamp 1704896540
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_137
timestamp 1704896540
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_149
timestamp 1704896540
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_161
timestamp 1704896540
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_167
timestamp 1704896540
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_169
timestamp 1704896540
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_181
timestamp 1704896540
transform 1 0 17756 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_191
timestamp 1704896540
transform 1 0 18676 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_203
timestamp 1704896540
transform 1 0 19780 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_215
timestamp 1704896540
transform 1 0 20884 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_223
timestamp 1704896540
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_225
timestamp 1704896540
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_237
timestamp 1704896540
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_249
timestamp 1704896540
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_261
timestamp 1704896540
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_273
timestamp 1704896540
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_279
timestamp 1704896540
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_281
timestamp 1704896540
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_293
timestamp 1704896540
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_305
timestamp 1704896540
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_317
timestamp 1704896540
transform 1 0 30268 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_325
timestamp 1704896540
transform 1 0 31004 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_331
timestamp 1704896540
transform 1 0 31556 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_335
timestamp 1704896540
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_337
timestamp 1704896540
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_349
timestamp 1704896540
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_361
timestamp 1704896540
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_373
timestamp 1704896540
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_385
timestamp 1704896540
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_391
timestamp 1704896540
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_416
timestamp 1704896540
transform 1 0 39376 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_428
timestamp 1704896540
transform 1 0 40480 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_3
timestamp 1704896540
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_15
timestamp 1704896540
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_27
timestamp 1704896540
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_29
timestamp 1704896540
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_41
timestamp 1704896540
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_53
timestamp 1704896540
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_65
timestamp 1704896540
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_77
timestamp 1704896540
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_83
timestamp 1704896540
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_85
timestamp 1704896540
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_97
timestamp 1704896540
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_109
timestamp 1704896540
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_121
timestamp 1704896540
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_133
timestamp 1704896540
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_139
timestamp 1704896540
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_141
timestamp 1704896540
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_153
timestamp 1704896540
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_165
timestamp 1704896540
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_177
timestamp 1704896540
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_189
timestamp 1704896540
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_195
timestamp 1704896540
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_197
timestamp 1704896540
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_209
timestamp 1704896540
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_221
timestamp 1704896540
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_233
timestamp 1704896540
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_245
timestamp 1704896540
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_251
timestamp 1704896540
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_253
timestamp 1704896540
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_265
timestamp 1704896540
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_277
timestamp 1704896540
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_289
timestamp 1704896540
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_301
timestamp 1704896540
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_307
timestamp 1704896540
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_309
timestamp 1704896540
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_321
timestamp 1704896540
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_333
timestamp 1704896540
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_345
timestamp 1704896540
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_357
timestamp 1704896540
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_363
timestamp 1704896540
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_365
timestamp 1704896540
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_377
timestamp 1704896540
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_389
timestamp 1704896540
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_401
timestamp 1704896540
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_413
timestamp 1704896540
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_419
timestamp 1704896540
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_421
timestamp 1704896540
transform 1 0 39836 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_3
timestamp 1704896540
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_15
timestamp 1704896540
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_27
timestamp 1704896540
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_39
timestamp 1704896540
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_51
timestamp 1704896540
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_55
timestamp 1704896540
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_57
timestamp 1704896540
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_69
timestamp 1704896540
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_81
timestamp 1704896540
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_93
timestamp 1704896540
transform 1 0 9660 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_99
timestamp 1704896540
transform 1 0 10212 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_103
timestamp 1704896540
transform 1 0 10580 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_111
timestamp 1704896540
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_113
timestamp 1704896540
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_125
timestamp 1704896540
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_137
timestamp 1704896540
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_149
timestamp 1704896540
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_161
timestamp 1704896540
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_167
timestamp 1704896540
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_169
timestamp 1704896540
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_181
timestamp 1704896540
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_193
timestamp 1704896540
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_205
timestamp 1704896540
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_217
timestamp 1704896540
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_223
timestamp 1704896540
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_225
timestamp 1704896540
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_237
timestamp 1704896540
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_249
timestamp 1704896540
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_261
timestamp 1704896540
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_273
timestamp 1704896540
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_279
timestamp 1704896540
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_281
timestamp 1704896540
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_293
timestamp 1704896540
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_305
timestamp 1704896540
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_317
timestamp 1704896540
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_329
timestamp 1704896540
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_335
timestamp 1704896540
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_337
timestamp 1704896540
transform 1 0 32108 0 -1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_348
timestamp 1704896540
transform 1 0 33120 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_360
timestamp 1704896540
transform 1 0 34224 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_372
timestamp 1704896540
transform 1 0 35328 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_384
timestamp 1704896540
transform 1 0 36432 0 -1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_393
timestamp 1704896540
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_405
timestamp 1704896540
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_417
timestamp 1704896540
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_3
timestamp 1704896540
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_15
timestamp 1704896540
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_27
timestamp 1704896540
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_29
timestamp 1704896540
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_41
timestamp 1704896540
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_53
timestamp 1704896540
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_65
timestamp 1704896540
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_77
timestamp 1704896540
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_83
timestamp 1704896540
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_85
timestamp 1704896540
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_97
timestamp 1704896540
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_109
timestamp 1704896540
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_121
timestamp 1704896540
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_133
timestamp 1704896540
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_139
timestamp 1704896540
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_141
timestamp 1704896540
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_153
timestamp 1704896540
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_165
timestamp 1704896540
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_177
timestamp 1704896540
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_189
timestamp 1704896540
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_195
timestamp 1704896540
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_197
timestamp 1704896540
transform 1 0 19228 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_221
timestamp 1704896540
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_233
timestamp 1704896540
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_245
timestamp 1704896540
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_251
timestamp 1704896540
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_262
timestamp 1704896540
transform 1 0 25208 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_274
timestamp 1704896540
transform 1 0 26312 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_286
timestamp 1704896540
transform 1 0 27416 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_298
timestamp 1704896540
transform 1 0 28520 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_306
timestamp 1704896540
transform 1 0 29256 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_309
timestamp 1704896540
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_321
timestamp 1704896540
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_333
timestamp 1704896540
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_345
timestamp 1704896540
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_357
timestamp 1704896540
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_363
timestamp 1704896540
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_365
timestamp 1704896540
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_377
timestamp 1704896540
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_389
timestamp 1704896540
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_401
timestamp 1704896540
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_413
timestamp 1704896540
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_419
timestamp 1704896540
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_421
timestamp 1704896540
transform 1 0 39836 0 1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_3
timestamp 1704896540
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_15
timestamp 1704896540
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_27
timestamp 1704896540
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_39
timestamp 1704896540
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_51
timestamp 1704896540
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_55
timestamp 1704896540
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_57
timestamp 1704896540
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_69
timestamp 1704896540
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_81
timestamp 1704896540
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_93
timestamp 1704896540
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_105
timestamp 1704896540
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_111
timestamp 1704896540
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_113
timestamp 1704896540
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_125
timestamp 1704896540
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_137
timestamp 1704896540
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_149
timestamp 1704896540
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_161
timestamp 1704896540
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_167
timestamp 1704896540
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_169
timestamp 1704896540
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_181
timestamp 1704896540
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_193
timestamp 1704896540
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_205
timestamp 1704896540
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_217
timestamp 1704896540
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_223
timestamp 1704896540
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_225
timestamp 1704896540
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_237
timestamp 1704896540
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_249
timestamp 1704896540
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_261
timestamp 1704896540
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_273
timestamp 1704896540
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_279
timestamp 1704896540
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_281
timestamp 1704896540
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_293
timestamp 1704896540
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_305
timestamp 1704896540
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_317
timestamp 1704896540
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_329
timestamp 1704896540
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_335
timestamp 1704896540
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_337
timestamp 1704896540
transform 1 0 32108 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_341
timestamp 1704896540
transform 1 0 32476 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_347
timestamp 1704896540
transform 1 0 33028 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_359
timestamp 1704896540
transform 1 0 34132 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_371
timestamp 1704896540
transform 1 0 35236 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_383
timestamp 1704896540
transform 1 0 36340 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_391
timestamp 1704896540
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_393
timestamp 1704896540
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_405
timestamp 1704896540
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_417
timestamp 1704896540
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_3
timestamp 1704896540
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_15
timestamp 1704896540
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_27
timestamp 1704896540
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_29
timestamp 1704896540
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_41
timestamp 1704896540
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_53
timestamp 1704896540
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_65
timestamp 1704896540
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_77
timestamp 1704896540
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_83
timestamp 1704896540
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_85
timestamp 1704896540
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_97
timestamp 1704896540
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_109
timestamp 1704896540
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_121
timestamp 1704896540
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_133
timestamp 1704896540
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_139
timestamp 1704896540
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_141
timestamp 1704896540
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_153
timestamp 1704896540
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_165
timestamp 1704896540
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_177
timestamp 1704896540
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_189
timestamp 1704896540
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_195
timestamp 1704896540
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_197
timestamp 1704896540
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_209
timestamp 1704896540
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_221
timestamp 1704896540
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_233
timestamp 1704896540
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_245
timestamp 1704896540
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_251
timestamp 1704896540
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_253
timestamp 1704896540
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_265
timestamp 1704896540
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_277
timestamp 1704896540
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_289
timestamp 1704896540
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_301
timestamp 1704896540
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_307
timestamp 1704896540
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_309
timestamp 1704896540
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_321
timestamp 1704896540
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_333
timestamp 1704896540
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_345
timestamp 1704896540
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_357
timestamp 1704896540
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_363
timestamp 1704896540
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_365
timestamp 1704896540
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_377
timestamp 1704896540
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_389
timestamp 1704896540
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_401
timestamp 1704896540
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_413
timestamp 1704896540
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_419
timestamp 1704896540
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_421
timestamp 1704896540
transform 1 0 39836 0 1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_3
timestamp 1704896540
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_15
timestamp 1704896540
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_27
timestamp 1704896540
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_39
timestamp 1704896540
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_51
timestamp 1704896540
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_55
timestamp 1704896540
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_57
timestamp 1704896540
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_69
timestamp 1704896540
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_81
timestamp 1704896540
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_93
timestamp 1704896540
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_105
timestamp 1704896540
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_111
timestamp 1704896540
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_113
timestamp 1704896540
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_125
timestamp 1704896540
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_137
timestamp 1704896540
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_149
timestamp 1704896540
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_161
timestamp 1704896540
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_167
timestamp 1704896540
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_169
timestamp 1704896540
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_181
timestamp 1704896540
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_193
timestamp 1704896540
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_205
timestamp 1704896540
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_217
timestamp 1704896540
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_223
timestamp 1704896540
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_225
timestamp 1704896540
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_237
timestamp 1704896540
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_249
timestamp 1704896540
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_261
timestamp 1704896540
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_273
timestamp 1704896540
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_279
timestamp 1704896540
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_281
timestamp 1704896540
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_293
timestamp 1704896540
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_305
timestamp 1704896540
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_317
timestamp 1704896540
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_329
timestamp 1704896540
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_335
timestamp 1704896540
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_337
timestamp 1704896540
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_349
timestamp 1704896540
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_363
timestamp 1704896540
transform 1 0 34500 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_374
timestamp 1704896540
transform 1 0 35512 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_386
timestamp 1704896540
transform 1 0 36616 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_393
timestamp 1704896540
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_405
timestamp 1704896540
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_417
timestamp 1704896540
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_3
timestamp 1704896540
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_15
timestamp 1704896540
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_27
timestamp 1704896540
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_29
timestamp 1704896540
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_41
timestamp 1704896540
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_53
timestamp 1704896540
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_65
timestamp 1704896540
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_77
timestamp 1704896540
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_83
timestamp 1704896540
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_92
timestamp 1704896540
transform 1 0 9568 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_104
timestamp 1704896540
transform 1 0 10672 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_116
timestamp 1704896540
transform 1 0 11776 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_128
timestamp 1704896540
transform 1 0 12880 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_141
timestamp 1704896540
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_153
timestamp 1704896540
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_165
timestamp 1704896540
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_177
timestamp 1704896540
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_189
timestamp 1704896540
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_195
timestamp 1704896540
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_197
timestamp 1704896540
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_209
timestamp 1704896540
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_221
timestamp 1704896540
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_233
timestamp 1704896540
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_245
timestamp 1704896540
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_251
timestamp 1704896540
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_253
timestamp 1704896540
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_265
timestamp 1704896540
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_277
timestamp 1704896540
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_289
timestamp 1704896540
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_301
timestamp 1704896540
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_307
timestamp 1704896540
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_309
timestamp 1704896540
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_321
timestamp 1704896540
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_333
timestamp 1704896540
transform 1 0 31740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_341
timestamp 1704896540
transform 1 0 32476 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_353
timestamp 1704896540
transform 1 0 33580 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_361
timestamp 1704896540
transform 1 0 34316 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_365
timestamp 1704896540
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_377
timestamp 1704896540
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_389
timestamp 1704896540
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_401
timestamp 1704896540
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_413
timestamp 1704896540
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_419
timestamp 1704896540
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_421
timestamp 1704896540
transform 1 0 39836 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_3
timestamp 1704896540
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_15
timestamp 1704896540
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_27
timestamp 1704896540
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_39
timestamp 1704896540
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_51
timestamp 1704896540
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_55
timestamp 1704896540
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_57
timestamp 1704896540
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_71
timestamp 1704896540
transform 1 0 7636 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_96
timestamp 1704896540
transform 1 0 9936 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_108
timestamp 1704896540
transform 1 0 11040 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_113
timestamp 1704896540
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_125
timestamp 1704896540
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_137
timestamp 1704896540
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_149
timestamp 1704896540
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_161
timestamp 1704896540
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_167
timestamp 1704896540
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_169
timestamp 1704896540
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_181
timestamp 1704896540
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_193
timestamp 1704896540
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_205
timestamp 1704896540
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_217
timestamp 1704896540
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_223
timestamp 1704896540
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_225
timestamp 1704896540
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_237
timestamp 1704896540
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_249
timestamp 1704896540
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_261
timestamp 1704896540
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_273
timestamp 1704896540
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_279
timestamp 1704896540
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_284
timestamp 1704896540
transform 1 0 27232 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_296
timestamp 1704896540
transform 1 0 28336 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_308
timestamp 1704896540
transform 1 0 29440 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_320
timestamp 1704896540
transform 1 0 30544 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_332
timestamp 1704896540
transform 1 0 31648 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_337
timestamp 1704896540
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_349
timestamp 1704896540
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_361
timestamp 1704896540
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_373
timestamp 1704896540
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_385
timestamp 1704896540
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_391
timestamp 1704896540
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_393
timestamp 1704896540
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_405
timestamp 1704896540
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_417
timestamp 1704896540
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_3
timestamp 1704896540
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_15
timestamp 1704896540
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_27
timestamp 1704896540
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_29
timestamp 1704896540
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_41
timestamp 1704896540
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_53
timestamp 1704896540
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_65
timestamp 1704896540
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_77
timestamp 1704896540
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_83
timestamp 1704896540
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_85
timestamp 1704896540
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_97
timestamp 1704896540
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_109
timestamp 1704896540
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_121
timestamp 1704896540
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_133
timestamp 1704896540
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_139
timestamp 1704896540
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_141
timestamp 1704896540
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_153
timestamp 1704896540
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_165
timestamp 1704896540
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_177
timestamp 1704896540
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_189
timestamp 1704896540
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_195
timestamp 1704896540
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_197
timestamp 1704896540
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_209
timestamp 1704896540
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_221
timestamp 1704896540
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_233
timestamp 1704896540
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_245
timestamp 1704896540
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_251
timestamp 1704896540
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_253
timestamp 1704896540
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_265
timestamp 1704896540
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_277
timestamp 1704896540
transform 1 0 26588 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_285
timestamp 1704896540
transform 1 0 27324 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_291
timestamp 1704896540
transform 1 0 27876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_303
timestamp 1704896540
transform 1 0 28980 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_307
timestamp 1704896540
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_309
timestamp 1704896540
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_321
timestamp 1704896540
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_333
timestamp 1704896540
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_345
timestamp 1704896540
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_357
timestamp 1704896540
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_363
timestamp 1704896540
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_365
timestamp 1704896540
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_377
timestamp 1704896540
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_389
timestamp 1704896540
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_401
timestamp 1704896540
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_413
timestamp 1704896540
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_419
timestamp 1704896540
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_421
timestamp 1704896540
transform 1 0 39836 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_3
timestamp 1704896540
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_15
timestamp 1704896540
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_27
timestamp 1704896540
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_39
timestamp 1704896540
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_51
timestamp 1704896540
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_55
timestamp 1704896540
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_57
timestamp 1704896540
transform 1 0 6348 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_63
timestamp 1704896540
transform 1 0 6900 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_67
timestamp 1704896540
transform 1 0 7268 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_79
timestamp 1704896540
transform 1 0 8372 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_91
timestamp 1704896540
transform 1 0 9476 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_103
timestamp 1704896540
transform 1 0 10580 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_111
timestamp 1704896540
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_113
timestamp 1704896540
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_125
timestamp 1704896540
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_137
timestamp 1704896540
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_149
timestamp 1704896540
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_161
timestamp 1704896540
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_167
timestamp 1704896540
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_169
timestamp 1704896540
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_181
timestamp 1704896540
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_193
timestamp 1704896540
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_205
timestamp 1704896540
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_217
timestamp 1704896540
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_223
timestamp 1704896540
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_225
timestamp 1704896540
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_237
timestamp 1704896540
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_249
timestamp 1704896540
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_261
timestamp 1704896540
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_273
timestamp 1704896540
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_279
timestamp 1704896540
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_281
timestamp 1704896540
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_293
timestamp 1704896540
transform 1 0 28060 0 -1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_308
timestamp 1704896540
transform 1 0 29440 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_320
timestamp 1704896540
transform 1 0 30544 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_332
timestamp 1704896540
transform 1 0 31648 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_337
timestamp 1704896540
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_349
timestamp 1704896540
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_361
timestamp 1704896540
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_373
timestamp 1704896540
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_385
timestamp 1704896540
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_391
timestamp 1704896540
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_393
timestamp 1704896540
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_405
timestamp 1704896540
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_417
timestamp 1704896540
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_3
timestamp 1704896540
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_15
timestamp 1704896540
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_27
timestamp 1704896540
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_29
timestamp 1704896540
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_41
timestamp 1704896540
transform 1 0 4876 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_47
timestamp 1704896540
transform 1 0 5428 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_58
timestamp 1704896540
transform 1 0 6440 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_70
timestamp 1704896540
transform 1 0 7544 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_82
timestamp 1704896540
transform 1 0 8648 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_85
timestamp 1704896540
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_97
timestamp 1704896540
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_109
timestamp 1704896540
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_121
timestamp 1704896540
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_133
timestamp 1704896540
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_139
timestamp 1704896540
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_141
timestamp 1704896540
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_153
timestamp 1704896540
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_165
timestamp 1704896540
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_177
timestamp 1704896540
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_189
timestamp 1704896540
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_195
timestamp 1704896540
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_197
timestamp 1704896540
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_209
timestamp 1704896540
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_221
timestamp 1704896540
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_233
timestamp 1704896540
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_245
timestamp 1704896540
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_251
timestamp 1704896540
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_253
timestamp 1704896540
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_265
timestamp 1704896540
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_277
timestamp 1704896540
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_289
timestamp 1704896540
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_301
timestamp 1704896540
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_307
timestamp 1704896540
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_309
timestamp 1704896540
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_321
timestamp 1704896540
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_333
timestamp 1704896540
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_345
timestamp 1704896540
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_357
timestamp 1704896540
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_363
timestamp 1704896540
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_365
timestamp 1704896540
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_377
timestamp 1704896540
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_389
timestamp 1704896540
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_401
timestamp 1704896540
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_413
timestamp 1704896540
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_419
timestamp 1704896540
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_421
timestamp 1704896540
transform 1 0 39836 0 1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_3
timestamp 1704896540
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_15
timestamp 1704896540
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_27
timestamp 1704896540
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_39
timestamp 1704896540
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_51
timestamp 1704896540
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_55
timestamp 1704896540
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_57
timestamp 1704896540
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_69
timestamp 1704896540
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_81
timestamp 1704896540
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_93
timestamp 1704896540
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_105
timestamp 1704896540
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_111
timestamp 1704896540
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_113
timestamp 1704896540
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_125
timestamp 1704896540
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_137
timestamp 1704896540
transform 1 0 13708 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_144
timestamp 1704896540
transform 1 0 14352 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_156
timestamp 1704896540
transform 1 0 15456 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_169
timestamp 1704896540
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_181
timestamp 1704896540
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_193
timestamp 1704896540
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_205
timestamp 1704896540
transform 1 0 19964 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_213
timestamp 1704896540
transform 1 0 20700 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_248
timestamp 1704896540
transform 1 0 23920 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_252
timestamp 1704896540
transform 1 0 24288 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_264
timestamp 1704896540
transform 1 0 25392 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_276
timestamp 1704896540
transform 1 0 26496 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_281
timestamp 1704896540
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_293
timestamp 1704896540
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_305
timestamp 1704896540
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_317
timestamp 1704896540
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_329
timestamp 1704896540
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_335
timestamp 1704896540
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_337
timestamp 1704896540
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_349
timestamp 1704896540
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_361
timestamp 1704896540
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_373
timestamp 1704896540
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_385
timestamp 1704896540
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_391
timestamp 1704896540
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_393
timestamp 1704896540
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_405
timestamp 1704896540
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_417
timestamp 1704896540
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_3
timestamp 1704896540
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_15
timestamp 1704896540
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_27
timestamp 1704896540
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_29
timestamp 1704896540
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_41
timestamp 1704896540
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_53
timestamp 1704896540
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_65
timestamp 1704896540
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_77
timestamp 1704896540
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_83
timestamp 1704896540
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_85
timestamp 1704896540
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_97
timestamp 1704896540
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_109
timestamp 1704896540
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_121
timestamp 1704896540
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_133
timestamp 1704896540
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_139
timestamp 1704896540
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_141
timestamp 1704896540
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_153
timestamp 1704896540
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_165
timestamp 1704896540
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_177
timestamp 1704896540
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_189
timestamp 1704896540
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_195
timestamp 1704896540
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_197
timestamp 1704896540
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_209
timestamp 1704896540
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_221
timestamp 1704896540
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_233
timestamp 1704896540
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_245
timestamp 1704896540
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_251
timestamp 1704896540
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_253
timestamp 1704896540
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_265
timestamp 1704896540
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_277
timestamp 1704896540
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_289
timestamp 1704896540
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_301
timestamp 1704896540
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_307
timestamp 1704896540
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_309
timestamp 1704896540
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_321
timestamp 1704896540
transform 1 0 30636 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_325
timestamp 1704896540
transform 1 0 31004 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_337
timestamp 1704896540
transform 1 0 32108 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_349
timestamp 1704896540
transform 1 0 33212 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_361
timestamp 1704896540
transform 1 0 34316 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_365
timestamp 1704896540
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_377
timestamp 1704896540
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_389
timestamp 1704896540
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_401
timestamp 1704896540
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_413
timestamp 1704896540
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_419
timestamp 1704896540
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_421
timestamp 1704896540
transform 1 0 39836 0 1 39168
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_3
timestamp 1704896540
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_15
timestamp 1704896540
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_27
timestamp 1704896540
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_39
timestamp 1704896540
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_51
timestamp 1704896540
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_55
timestamp 1704896540
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_57
timestamp 1704896540
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_69
timestamp 1704896540
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_81
timestamp 1704896540
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_93
timestamp 1704896540
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_105
timestamp 1704896540
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_111
timestamp 1704896540
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_113
timestamp 1704896540
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_125
timestamp 1704896540
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_137
timestamp 1704896540
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_149
timestamp 1704896540
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_161
timestamp 1704896540
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_167
timestamp 1704896540
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_169
timestamp 1704896540
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_181
timestamp 1704896540
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_193
timestamp 1704896540
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_205
timestamp 1704896540
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_217
timestamp 1704896540
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_223
timestamp 1704896540
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_225
timestamp 1704896540
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_237
timestamp 1704896540
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_249
timestamp 1704896540
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_261
timestamp 1704896540
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_273
timestamp 1704896540
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_279
timestamp 1704896540
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_281
timestamp 1704896540
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_293
timestamp 1704896540
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_305
timestamp 1704896540
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_317
timestamp 1704896540
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_329
timestamp 1704896540
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_335
timestamp 1704896540
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_337
timestamp 1704896540
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_349
timestamp 1704896540
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_361
timestamp 1704896540
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_373
timestamp 1704896540
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_385
timestamp 1704896540
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_391
timestamp 1704896540
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_393
timestamp 1704896540
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_405
timestamp 1704896540
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_417
timestamp 1704896540
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_3
timestamp 1704896540
transform 1 0 1380 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_70_11
timestamp 1704896540
transform 1 0 2116 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_29
timestamp 1704896540
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_41
timestamp 1704896540
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_53
timestamp 1704896540
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_65
timestamp 1704896540
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_77
timestamp 1704896540
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_83
timestamp 1704896540
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_85
timestamp 1704896540
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_97
timestamp 1704896540
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_109
timestamp 1704896540
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_121
timestamp 1704896540
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_133
timestamp 1704896540
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_139
timestamp 1704896540
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_141
timestamp 1704896540
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_153
timestamp 1704896540
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_165
timestamp 1704896540
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_177
timestamp 1704896540
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_189
timestamp 1704896540
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_195
timestamp 1704896540
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_197
timestamp 1704896540
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_209
timestamp 1704896540
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_221
timestamp 1704896540
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_233
timestamp 1704896540
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_245
timestamp 1704896540
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_251
timestamp 1704896540
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_253
timestamp 1704896540
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_265
timestamp 1704896540
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_277
timestamp 1704896540
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_289
timestamp 1704896540
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_301
timestamp 1704896540
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_307
timestamp 1704896540
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_309
timestamp 1704896540
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_321
timestamp 1704896540
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_333
timestamp 1704896540
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_345
timestamp 1704896540
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_357
timestamp 1704896540
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_363
timestamp 1704896540
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_365
timestamp 1704896540
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_377
timestamp 1704896540
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_389
timestamp 1704896540
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_401
timestamp 1704896540
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_413
timestamp 1704896540
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_419
timestamp 1704896540
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_421
timestamp 1704896540
transform 1 0 39836 0 1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_3
timestamp 1704896540
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_15
timestamp 1704896540
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_27
timestamp 1704896540
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_39
timestamp 1704896540
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71_51
timestamp 1704896540
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_55
timestamp 1704896540
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_71_57
timestamp 1704896540
transform 1 0 6348 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_77
timestamp 1704896540
transform 1 0 8188 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_89
timestamp 1704896540
transform 1 0 9292 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_71_101
timestamp 1704896540
transform 1 0 10396 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_71_109
timestamp 1704896540
transform 1 0 11132 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_113
timestamp 1704896540
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_125
timestamp 1704896540
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_137
timestamp 1704896540
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_149
timestamp 1704896540
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_161
timestamp 1704896540
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_167
timestamp 1704896540
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_169
timestamp 1704896540
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_181
timestamp 1704896540
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_193
timestamp 1704896540
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_205
timestamp 1704896540
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_217
timestamp 1704896540
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_223
timestamp 1704896540
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_225
timestamp 1704896540
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_237
timestamp 1704896540
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_249
timestamp 1704896540
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_71_261
timestamp 1704896540
transform 1 0 25116 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_267
timestamp 1704896540
transform 1 0 25668 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_279
timestamp 1704896540
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_281
timestamp 1704896540
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_293
timestamp 1704896540
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_305
timestamp 1704896540
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_317
timestamp 1704896540
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_329
timestamp 1704896540
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_335
timestamp 1704896540
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_337
timestamp 1704896540
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_349
timestamp 1704896540
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_361
timestamp 1704896540
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_373
timestamp 1704896540
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_385
timestamp 1704896540
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_391
timestamp 1704896540
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_393
timestamp 1704896540
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_405
timestamp 1704896540
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_417
timestamp 1704896540
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_3
timestamp 1704896540
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_15
timestamp 1704896540
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_27
timestamp 1704896540
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_29
timestamp 1704896540
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_41
timestamp 1704896540
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_53
timestamp 1704896540
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_65
timestamp 1704896540
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_77
timestamp 1704896540
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_83
timestamp 1704896540
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_85
timestamp 1704896540
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_97
timestamp 1704896540
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_109
timestamp 1704896540
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_121
timestamp 1704896540
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_133
timestamp 1704896540
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_139
timestamp 1704896540
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_141
timestamp 1704896540
transform 1 0 14076 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72_145
timestamp 1704896540
transform 1 0 14444 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_153
timestamp 1704896540
transform 1 0 15180 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_158
timestamp 1704896540
transform 1 0 15640 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_170
timestamp 1704896540
transform 1 0 16744 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_182
timestamp 1704896540
transform 1 0 17848 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_194
timestamp 1704896540
transform 1 0 18952 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_197
timestamp 1704896540
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_209
timestamp 1704896540
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_221
timestamp 1704896540
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_233
timestamp 1704896540
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_245
timestamp 1704896540
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_251
timestamp 1704896540
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72_253
timestamp 1704896540
transform 1 0 24380 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_280
timestamp 1704896540
transform 1 0 26864 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_292
timestamp 1704896540
transform 1 0 27968 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72_304
timestamp 1704896540
transform 1 0 29072 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_309
timestamp 1704896540
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_321
timestamp 1704896540
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_333
timestamp 1704896540
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_345
timestamp 1704896540
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_357
timestamp 1704896540
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_363
timestamp 1704896540
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_365
timestamp 1704896540
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72_377
timestamp 1704896540
transform 1 0 35788 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_387
timestamp 1704896540
transform 1 0 36708 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72_412
timestamp 1704896540
transform 1 0 39008 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72_421
timestamp 1704896540
transform 1 0 39836 0 1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_3
timestamp 1704896540
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_15
timestamp 1704896540
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_27
timestamp 1704896540
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_39
timestamp 1704896540
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73_51
timestamp 1704896540
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_55
timestamp 1704896540
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_57
timestamp 1704896540
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_69
timestamp 1704896540
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_81
timestamp 1704896540
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_93
timestamp 1704896540
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_105
timestamp 1704896540
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_111
timestamp 1704896540
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_113
timestamp 1704896540
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_125
timestamp 1704896540
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_137
timestamp 1704896540
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_149
timestamp 1704896540
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_161
timestamp 1704896540
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_167
timestamp 1704896540
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_169
timestamp 1704896540
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_181
timestamp 1704896540
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_193
timestamp 1704896540
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_205
timestamp 1704896540
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_217
timestamp 1704896540
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_223
timestamp 1704896540
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_225
timestamp 1704896540
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_237
timestamp 1704896540
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_249
timestamp 1704896540
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_261
timestamp 1704896540
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_273
timestamp 1704896540
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_279
timestamp 1704896540
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_281
timestamp 1704896540
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_293
timestamp 1704896540
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_305
timestamp 1704896540
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_317
timestamp 1704896540
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_329
timestamp 1704896540
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_335
timestamp 1704896540
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_337
timestamp 1704896540
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_349
timestamp 1704896540
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_361
timestamp 1704896540
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_373
timestamp 1704896540
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_385
timestamp 1704896540
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_391
timestamp 1704896540
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_393
timestamp 1704896540
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_405
timestamp 1704896540
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_417
timestamp 1704896540
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_3
timestamp 1704896540
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_15
timestamp 1704896540
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_27
timestamp 1704896540
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_29
timestamp 1704896540
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_41
timestamp 1704896540
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_53
timestamp 1704896540
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_65
timestamp 1704896540
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_77
timestamp 1704896540
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_83
timestamp 1704896540
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_85
timestamp 1704896540
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_97
timestamp 1704896540
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_109
timestamp 1704896540
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_121
timestamp 1704896540
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_133
timestamp 1704896540
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_139
timestamp 1704896540
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_141
timestamp 1704896540
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_153
timestamp 1704896540
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_165
timestamp 1704896540
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_177
timestamp 1704896540
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_189
timestamp 1704896540
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_195
timestamp 1704896540
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_197
timestamp 1704896540
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_209
timestamp 1704896540
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_221
timestamp 1704896540
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_233
timestamp 1704896540
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_245
timestamp 1704896540
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_251
timestamp 1704896540
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_253
timestamp 1704896540
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_265
timestamp 1704896540
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_277
timestamp 1704896540
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_289
timestamp 1704896540
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_301
timestamp 1704896540
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_307
timestamp 1704896540
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_309
timestamp 1704896540
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_321
timestamp 1704896540
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_333
timestamp 1704896540
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_345
timestamp 1704896540
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_357
timestamp 1704896540
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_363
timestamp 1704896540
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_365
timestamp 1704896540
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_377
timestamp 1704896540
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_389
timestamp 1704896540
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_401
timestamp 1704896540
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_413
timestamp 1704896540
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_419
timestamp 1704896540
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_74_421
timestamp 1704896540
transform 1 0 39836 0 1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_3
timestamp 1704896540
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_15
timestamp 1704896540
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_27
timestamp 1704896540
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_39
timestamp 1704896540
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75_51
timestamp 1704896540
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_55
timestamp 1704896540
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_57
timestamp 1704896540
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_69
timestamp 1704896540
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_81
timestamp 1704896540
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_93
timestamp 1704896540
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_105
timestamp 1704896540
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_111
timestamp 1704896540
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_113
timestamp 1704896540
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_125
timestamp 1704896540
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_137
timestamp 1704896540
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_149
timestamp 1704896540
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_161
timestamp 1704896540
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_167
timestamp 1704896540
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_169
timestamp 1704896540
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_181
timestamp 1704896540
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_193
timestamp 1704896540
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_205
timestamp 1704896540
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_217
timestamp 1704896540
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_223
timestamp 1704896540
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_225
timestamp 1704896540
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_237
timestamp 1704896540
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_249
timestamp 1704896540
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_261
timestamp 1704896540
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_273
timestamp 1704896540
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_279
timestamp 1704896540
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_281
timestamp 1704896540
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_293
timestamp 1704896540
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_305
timestamp 1704896540
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_317
timestamp 1704896540
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_329
timestamp 1704896540
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_335
timestamp 1704896540
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_337
timestamp 1704896540
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_349
timestamp 1704896540
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_361
timestamp 1704896540
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_373
timestamp 1704896540
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_385
timestamp 1704896540
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_391
timestamp 1704896540
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_393
timestamp 1704896540
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_405
timestamp 1704896540
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_417
timestamp 1704896540
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_3
timestamp 1704896540
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_15
timestamp 1704896540
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_27
timestamp 1704896540
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_29
timestamp 1704896540
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_41
timestamp 1704896540
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_53
timestamp 1704896540
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_65
timestamp 1704896540
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_77
timestamp 1704896540
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_83
timestamp 1704896540
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_85
timestamp 1704896540
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_97
timestamp 1704896540
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_109
timestamp 1704896540
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_121
timestamp 1704896540
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_133
timestamp 1704896540
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_139
timestamp 1704896540
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_141
timestamp 1704896540
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_153
timestamp 1704896540
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_165
timestamp 1704896540
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_177
timestamp 1704896540
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_189
timestamp 1704896540
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_195
timestamp 1704896540
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_197
timestamp 1704896540
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_209
timestamp 1704896540
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_221
timestamp 1704896540
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_233
timestamp 1704896540
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_245
timestamp 1704896540
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_251
timestamp 1704896540
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_76_253
timestamp 1704896540
transform 1 0 24380 0 1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_266
timestamp 1704896540
transform 1 0 25576 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_278
timestamp 1704896540
transform 1 0 26680 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_290
timestamp 1704896540
transform 1 0 27784 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_302
timestamp 1704896540
transform 1 0 28888 0 1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_309
timestamp 1704896540
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_321
timestamp 1704896540
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_333
timestamp 1704896540
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_345
timestamp 1704896540
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_357
timestamp 1704896540
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_363
timestamp 1704896540
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_365
timestamp 1704896540
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_377
timestamp 1704896540
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_389
timestamp 1704896540
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_401
timestamp 1704896540
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_413
timestamp 1704896540
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_419
timestamp 1704896540
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76_421
timestamp 1704896540
transform 1 0 39836 0 1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_3
timestamp 1704896540
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_15
timestamp 1704896540
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_27
timestamp 1704896540
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_39
timestamp 1704896540
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_77_51
timestamp 1704896540
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_55
timestamp 1704896540
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_57
timestamp 1704896540
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_69
timestamp 1704896540
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_81
timestamp 1704896540
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_93
timestamp 1704896540
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_105
timestamp 1704896540
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_111
timestamp 1704896540
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_113
timestamp 1704896540
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_125
timestamp 1704896540
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_137
timestamp 1704896540
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_149
timestamp 1704896540
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_161
timestamp 1704896540
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_167
timestamp 1704896540
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_169
timestamp 1704896540
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_181
timestamp 1704896540
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_193
timestamp 1704896540
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_205
timestamp 1704896540
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_217
timestamp 1704896540
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_223
timestamp 1704896540
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_225
timestamp 1704896540
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_237
timestamp 1704896540
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_249
timestamp 1704896540
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_261
timestamp 1704896540
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_273
timestamp 1704896540
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_279
timestamp 1704896540
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_281
timestamp 1704896540
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_293
timestamp 1704896540
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_305
timestamp 1704896540
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_317
timestamp 1704896540
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_329
timestamp 1704896540
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_335
timestamp 1704896540
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_337
timestamp 1704896540
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_349
timestamp 1704896540
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_361
timestamp 1704896540
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_373
timestamp 1704896540
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_385
timestamp 1704896540
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_391
timestamp 1704896540
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_393
timestamp 1704896540
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_405
timestamp 1704896540
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_417
timestamp 1704896540
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_3
timestamp 1704896540
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_15
timestamp 1704896540
transform 1 0 2484 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_78_25
timestamp 1704896540
transform 1 0 3404 0 1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_29
timestamp 1704896540
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_41
timestamp 1704896540
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_53
timestamp 1704896540
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_65
timestamp 1704896540
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_77
timestamp 1704896540
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_83
timestamp 1704896540
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_85
timestamp 1704896540
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_97
timestamp 1704896540
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_109
timestamp 1704896540
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_121
timestamp 1704896540
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_133
timestamp 1704896540
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_139
timestamp 1704896540
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_141
timestamp 1704896540
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_153
timestamp 1704896540
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_165
timestamp 1704896540
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_177
timestamp 1704896540
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_189
timestamp 1704896540
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_195
timestamp 1704896540
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_197
timestamp 1704896540
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_209
timestamp 1704896540
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_78_221
timestamp 1704896540
transform 1 0 21436 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_78_229
timestamp 1704896540
transform 1 0 22172 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_237
timestamp 1704896540
transform 1 0 22908 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_78_249
timestamp 1704896540
transform 1 0 24012 0 1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_253
timestamp 1704896540
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_265
timestamp 1704896540
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_277
timestamp 1704896540
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_289
timestamp 1704896540
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_301
timestamp 1704896540
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_307
timestamp 1704896540
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_309
timestamp 1704896540
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_321
timestamp 1704896540
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_333
timestamp 1704896540
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_345
timestamp 1704896540
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_357
timestamp 1704896540
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_363
timestamp 1704896540
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_365
timestamp 1704896540
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_377
timestamp 1704896540
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_389
timestamp 1704896540
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_401
timestamp 1704896540
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_413
timestamp 1704896540
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_419
timestamp 1704896540
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_78_421
timestamp 1704896540
transform 1 0 39836 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_79_26
timestamp 1704896540
transform 1 0 3496 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_30
timestamp 1704896540
transform 1 0 3864 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_42
timestamp 1704896540
transform 1 0 4968 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_79_54
timestamp 1704896540
transform 1 0 6072 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_57
timestamp 1704896540
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_69
timestamp 1704896540
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_81
timestamp 1704896540
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_93
timestamp 1704896540
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_105
timestamp 1704896540
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_111
timestamp 1704896540
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_113
timestamp 1704896540
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_125
timestamp 1704896540
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_137
timestamp 1704896540
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_149
timestamp 1704896540
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_161
timestamp 1704896540
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_167
timestamp 1704896540
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_169
timestamp 1704896540
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_181
timestamp 1704896540
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_193
timestamp 1704896540
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_205
timestamp 1704896540
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_217
timestamp 1704896540
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_223
timestamp 1704896540
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_225
timestamp 1704896540
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_237
timestamp 1704896540
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_79_249
timestamp 1704896540
transform 1 0 24012 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_257
timestamp 1704896540
transform 1 0 24748 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_261
timestamp 1704896540
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_273
timestamp 1704896540
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_279
timestamp 1704896540
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_281
timestamp 1704896540
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_293
timestamp 1704896540
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_305
timestamp 1704896540
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_317
timestamp 1704896540
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_329
timestamp 1704896540
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_335
timestamp 1704896540
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_337
timestamp 1704896540
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_349
timestamp 1704896540
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_361
timestamp 1704896540
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_373
timestamp 1704896540
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_385
timestamp 1704896540
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_391
timestamp 1704896540
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_393
timestamp 1704896540
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_405
timestamp 1704896540
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_417
timestamp 1704896540
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_3
timestamp 1704896540
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_15
timestamp 1704896540
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_27
timestamp 1704896540
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_29
timestamp 1704896540
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_41
timestamp 1704896540
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_53
timestamp 1704896540
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_65
timestamp 1704896540
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_77
timestamp 1704896540
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_83
timestamp 1704896540
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_85
timestamp 1704896540
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_97
timestamp 1704896540
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_109
timestamp 1704896540
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_121
timestamp 1704896540
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_133
timestamp 1704896540
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_139
timestamp 1704896540
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_141
timestamp 1704896540
transform 1 0 14076 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_166
timestamp 1704896540
transform 1 0 16376 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_178
timestamp 1704896540
transform 1 0 17480 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_80_193
timestamp 1704896540
transform 1 0 18860 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_197
timestamp 1704896540
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_209
timestamp 1704896540
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_221
timestamp 1704896540
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_233
timestamp 1704896540
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_245
timestamp 1704896540
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_251
timestamp 1704896540
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_253
timestamp 1704896540
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_265
timestamp 1704896540
transform 1 0 25484 0 1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_277
timestamp 1704896540
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_289
timestamp 1704896540
transform 1 0 27692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_307
timestamp 1704896540
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_309
timestamp 1704896540
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_321
timestamp 1704896540
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_333
timestamp 1704896540
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_345
timestamp 1704896540
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_357
timestamp 1704896540
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_363
timestamp 1704896540
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_365
timestamp 1704896540
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_377
timestamp 1704896540
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_389
timestamp 1704896540
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_401
timestamp 1704896540
transform 1 0 37996 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_413
timestamp 1704896540
transform 1 0 39100 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_419
timestamp 1704896540
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_80_421
timestamp 1704896540
transform 1 0 39836 0 1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_3
timestamp 1704896540
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_15
timestamp 1704896540
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_27
timestamp 1704896540
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_39
timestamp 1704896540
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_81_51
timestamp 1704896540
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_55
timestamp 1704896540
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_57
timestamp 1704896540
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_69
timestamp 1704896540
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_81
timestamp 1704896540
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_93
timestamp 1704896540
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_105
timestamp 1704896540
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_111
timestamp 1704896540
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_113
timestamp 1704896540
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_125
timestamp 1704896540
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_137
timestamp 1704896540
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_149
timestamp 1704896540
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_161
timestamp 1704896540
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_167
timestamp 1704896540
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_169
timestamp 1704896540
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_181
timestamp 1704896540
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_193
timestamp 1704896540
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_205
timestamp 1704896540
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_217
timestamp 1704896540
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_223
timestamp 1704896540
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_225
timestamp 1704896540
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_237
timestamp 1704896540
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_249
timestamp 1704896540
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_261
timestamp 1704896540
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_273
timestamp 1704896540
transform 1 0 26220 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_279
timestamp 1704896540
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_281
timestamp 1704896540
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_81_293
timestamp 1704896540
transform 1 0 28060 0 -1 46784
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_321
timestamp 1704896540
transform 1 0 30636 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81_333
timestamp 1704896540
transform 1 0 31740 0 -1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_337
timestamp 1704896540
transform 1 0 32108 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_349
timestamp 1704896540
transform 1 0 33212 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_361
timestamp 1704896540
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_373
timestamp 1704896540
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_385
timestamp 1704896540
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_391
timestamp 1704896540
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_393
timestamp 1704896540
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_405
timestamp 1704896540
transform 1 0 38364 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_417
timestamp 1704896540
transform 1 0 39468 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_82_3
timestamp 1704896540
transform 1 0 1380 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_9
timestamp 1704896540
transform 1 0 1932 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_21
timestamp 1704896540
transform 1 0 3036 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_27
timestamp 1704896540
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_29
timestamp 1704896540
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_41
timestamp 1704896540
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_53
timestamp 1704896540
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_65
timestamp 1704896540
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_77
timestamp 1704896540
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_83
timestamp 1704896540
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_82_85
timestamp 1704896540
transform 1 0 8924 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_82_93
timestamp 1704896540
transform 1 0 9660 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_108
timestamp 1704896540
transform 1 0 11040 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_120
timestamp 1704896540
transform 1 0 12144 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_82_132
timestamp 1704896540
transform 1 0 13248 0 1 46784
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_141
timestamp 1704896540
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_153
timestamp 1704896540
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_165
timestamp 1704896540
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_177
timestamp 1704896540
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_189
timestamp 1704896540
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_195
timestamp 1704896540
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_197
timestamp 1704896540
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_209
timestamp 1704896540
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_221
timestamp 1704896540
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_233
timestamp 1704896540
transform 1 0 22540 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_245
timestamp 1704896540
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_251
timestamp 1704896540
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_253
timestamp 1704896540
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_265
timestamp 1704896540
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_277
timestamp 1704896540
transform 1 0 26588 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_289
timestamp 1704896540
transform 1 0 27692 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_301
timestamp 1704896540
transform 1 0 28796 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_307
timestamp 1704896540
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_309
timestamp 1704896540
transform 1 0 29532 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_321
timestamp 1704896540
transform 1 0 30636 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_333
timestamp 1704896540
transform 1 0 31740 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_345
timestamp 1704896540
transform 1 0 32844 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_357
timestamp 1704896540
transform 1 0 33948 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_363
timestamp 1704896540
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_365
timestamp 1704896540
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_82_377
timestamp 1704896540
transform 1 0 35788 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_381
timestamp 1704896540
transform 1 0 36156 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82_384
timestamp 1704896540
transform 1 0 36432 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82_388
timestamp 1704896540
transform 1 0 36800 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82_396
timestamp 1704896540
transform 1 0 37536 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_400
timestamp 1704896540
transform 1 0 37904 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_82_412
timestamp 1704896540
transform 1 0 39008 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_82_421
timestamp 1704896540
transform 1 0 39836 0 1 46784
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_3
timestamp 1704896540
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_15
timestamp 1704896540
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_27
timestamp 1704896540
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_39
timestamp 1704896540
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_83_51
timestamp 1704896540
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_55
timestamp 1704896540
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_57
timestamp 1704896540
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_69
timestamp 1704896540
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_81
timestamp 1704896540
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_93
timestamp 1704896540
transform 1 0 9660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_105
timestamp 1704896540
transform 1 0 10764 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_111
timestamp 1704896540
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_113
timestamp 1704896540
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_125
timestamp 1704896540
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_137
timestamp 1704896540
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_149
timestamp 1704896540
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_161
timestamp 1704896540
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_167
timestamp 1704896540
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_169
timestamp 1704896540
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_181
timestamp 1704896540
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_193
timestamp 1704896540
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_205
timestamp 1704896540
transform 1 0 19964 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_217
timestamp 1704896540
transform 1 0 21068 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_223
timestamp 1704896540
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_225
timestamp 1704896540
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_237
timestamp 1704896540
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_249
timestamp 1704896540
transform 1 0 24012 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_261
timestamp 1704896540
transform 1 0 25116 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_273
timestamp 1704896540
transform 1 0 26220 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_279
timestamp 1704896540
transform 1 0 26772 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_281
timestamp 1704896540
transform 1 0 26956 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_293
timestamp 1704896540
transform 1 0 28060 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_305
timestamp 1704896540
transform 1 0 29164 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_317
timestamp 1704896540
transform 1 0 30268 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_329
timestamp 1704896540
transform 1 0 31372 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_335
timestamp 1704896540
transform 1 0 31924 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_337
timestamp 1704896540
transform 1 0 32108 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_349
timestamp 1704896540
transform 1 0 33212 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_83_361
timestamp 1704896540
transform 1 0 34316 0 -1 47872
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_372
timestamp 1704896540
transform 1 0 35328 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_83_384
timestamp 1704896540
transform 1 0 36432 0 -1 47872
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_393
timestamp 1704896540
transform 1 0 37260 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_405
timestamp 1704896540
transform 1 0 38364 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_417
timestamp 1704896540
transform 1 0 39468 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_84_3
timestamp 1704896540
transform 1 0 1380 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_84_20
timestamp 1704896540
transform 1 0 2944 0 1 47872
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_29
timestamp 1704896540
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_41
timestamp 1704896540
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_53
timestamp 1704896540
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_65
timestamp 1704896540
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_77
timestamp 1704896540
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_83
timestamp 1704896540
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_85
timestamp 1704896540
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_97
timestamp 1704896540
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_109
timestamp 1704896540
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_121
timestamp 1704896540
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_133
timestamp 1704896540
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_139
timestamp 1704896540
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_141
timestamp 1704896540
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_153
timestamp 1704896540
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_165
timestamp 1704896540
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_177
timestamp 1704896540
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_189
timestamp 1704896540
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_195
timestamp 1704896540
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_197
timestamp 1704896540
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_209
timestamp 1704896540
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_221
timestamp 1704896540
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_233
timestamp 1704896540
transform 1 0 22540 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_245
timestamp 1704896540
transform 1 0 23644 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_251
timestamp 1704896540
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_253
timestamp 1704896540
transform 1 0 24380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_265
timestamp 1704896540
transform 1 0 25484 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_277
timestamp 1704896540
transform 1 0 26588 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_289
timestamp 1704896540
transform 1 0 27692 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_301
timestamp 1704896540
transform 1 0 28796 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_307
timestamp 1704896540
transform 1 0 29348 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_321
timestamp 1704896540
transform 1 0 30636 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_333
timestamp 1704896540
transform 1 0 31740 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_345
timestamp 1704896540
transform 1 0 32844 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_351
timestamp 1704896540
transform 1 0 33396 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_84_354
timestamp 1704896540
transform 1 0 33672 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_363
timestamp 1704896540
transform 1 0 34500 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_365
timestamp 1704896540
transform 1 0 34684 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_377
timestamp 1704896540
transform 1 0 35788 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_389
timestamp 1704896540
transform 1 0 36892 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_401
timestamp 1704896540
transform 1 0 37996 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_413
timestamp 1704896540
transform 1 0 39100 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_419
timestamp 1704896540
transform 1 0 39652 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_84_421
timestamp 1704896540
transform 1 0 39836 0 1 47872
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_3
timestamp 1704896540
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_15
timestamp 1704896540
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_27
timestamp 1704896540
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_39
timestamp 1704896540
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85_51
timestamp 1704896540
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_55
timestamp 1704896540
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_57
timestamp 1704896540
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_69
timestamp 1704896540
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_81
timestamp 1704896540
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_93
timestamp 1704896540
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85_105
timestamp 1704896540
transform 1 0 10764 0 -1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_113
timestamp 1704896540
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_125
timestamp 1704896540
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_137
timestamp 1704896540
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_149
timestamp 1704896540
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_161
timestamp 1704896540
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_167
timestamp 1704896540
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_169
timestamp 1704896540
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_181
timestamp 1704896540
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_193
timestamp 1704896540
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_205
timestamp 1704896540
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85_217
timestamp 1704896540
transform 1 0 21068 0 -1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_225
timestamp 1704896540
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_237
timestamp 1704896540
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_249
timestamp 1704896540
transform 1 0 24012 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_261
timestamp 1704896540
transform 1 0 25116 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_273
timestamp 1704896540
transform 1 0 26220 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_279
timestamp 1704896540
transform 1 0 26772 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_281
timestamp 1704896540
transform 1 0 26956 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_293
timestamp 1704896540
transform 1 0 28060 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_305
timestamp 1704896540
transform 1 0 29164 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_317
timestamp 1704896540
transform 1 0 30268 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_329
timestamp 1704896540
transform 1 0 31372 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_335
timestamp 1704896540
transform 1 0 31924 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_337
timestamp 1704896540
transform 1 0 32108 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_349
timestamp 1704896540
transform 1 0 33212 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_361
timestamp 1704896540
transform 1 0 34316 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_373
timestamp 1704896540
transform 1 0 35420 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_385
timestamp 1704896540
transform 1 0 36524 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_391
timestamp 1704896540
transform 1 0 37076 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_393
timestamp 1704896540
transform 1 0 37260 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_405
timestamp 1704896540
transform 1 0 38364 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_417
timestamp 1704896540
transform 1 0 39468 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_3
timestamp 1704896540
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_15
timestamp 1704896540
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_27
timestamp 1704896540
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_29
timestamp 1704896540
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_41
timestamp 1704896540
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_53
timestamp 1704896540
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_65
timestamp 1704896540
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_77
timestamp 1704896540
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_83
timestamp 1704896540
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_85
timestamp 1704896540
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_97
timestamp 1704896540
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_109
timestamp 1704896540
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_121
timestamp 1704896540
transform 1 0 12236 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_133
timestamp 1704896540
transform 1 0 13340 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_139
timestamp 1704896540
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_141
timestamp 1704896540
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_153
timestamp 1704896540
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_165
timestamp 1704896540
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_177
timestamp 1704896540
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_189
timestamp 1704896540
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_195
timestamp 1704896540
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_197
timestamp 1704896540
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_209
timestamp 1704896540
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_221
timestamp 1704896540
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_233
timestamp 1704896540
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_245
timestamp 1704896540
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_251
timestamp 1704896540
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_86_258
timestamp 1704896540
transform 1 0 24840 0 1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_262
timestamp 1704896540
transform 1 0 25208 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_274
timestamp 1704896540
transform 1 0 26312 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_286
timestamp 1704896540
transform 1 0 27416 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_86_298
timestamp 1704896540
transform 1 0 28520 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_86_306
timestamp 1704896540
transform 1 0 29256 0 1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_309
timestamp 1704896540
transform 1 0 29532 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_321
timestamp 1704896540
transform 1 0 30636 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_333
timestamp 1704896540
transform 1 0 31740 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_345
timestamp 1704896540
transform 1 0 32844 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_351
timestamp 1704896540
transform 1 0 33396 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_363
timestamp 1704896540
transform 1 0 34500 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_365
timestamp 1704896540
transform 1 0 34684 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_377
timestamp 1704896540
transform 1 0 35788 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_389
timestamp 1704896540
transform 1 0 36892 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_401
timestamp 1704896540
transform 1 0 37996 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_413
timestamp 1704896540
transform 1 0 39100 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_419
timestamp 1704896540
transform 1 0 39652 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_86_421
timestamp 1704896540
transform 1 0 39836 0 1 48960
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_3
timestamp 1704896540
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_15
timestamp 1704896540
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_27
timestamp 1704896540
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_39
timestamp 1704896540
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_87_51
timestamp 1704896540
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_55
timestamp 1704896540
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_57
timestamp 1704896540
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_69
timestamp 1704896540
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_81
timestamp 1704896540
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_93
timestamp 1704896540
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_105
timestamp 1704896540
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_111
timestamp 1704896540
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_113
timestamp 1704896540
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_125
timestamp 1704896540
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_137
timestamp 1704896540
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_149
timestamp 1704896540
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_161
timestamp 1704896540
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_167
timestamp 1704896540
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_169
timestamp 1704896540
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_181
timestamp 1704896540
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_193
timestamp 1704896540
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_205
timestamp 1704896540
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_217
timestamp 1704896540
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_223
timestamp 1704896540
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_225
timestamp 1704896540
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_237
timestamp 1704896540
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_249
timestamp 1704896540
transform 1 0 24012 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_261
timestamp 1704896540
transform 1 0 25116 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_273
timestamp 1704896540
transform 1 0 26220 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_279
timestamp 1704896540
transform 1 0 26772 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_281
timestamp 1704896540
transform 1 0 26956 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_87_293
timestamp 1704896540
transform 1 0 28060 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_87_301
timestamp 1704896540
transform 1 0 28796 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_308
timestamp 1704896540
transform 1 0 29440 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_320
timestamp 1704896540
transform 1 0 30544 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_87_332
timestamp 1704896540
transform 1 0 31648 0 -1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_337
timestamp 1704896540
transform 1 0 32108 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_349
timestamp 1704896540
transform 1 0 33212 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_361
timestamp 1704896540
transform 1 0 34316 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_373
timestamp 1704896540
transform 1 0 35420 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_385
timestamp 1704896540
transform 1 0 36524 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_391
timestamp 1704896540
transform 1 0 37076 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_393
timestamp 1704896540
transform 1 0 37260 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_405
timestamp 1704896540
transform 1 0 38364 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_417
timestamp 1704896540
transform 1 0 39468 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_3
timestamp 1704896540
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_15
timestamp 1704896540
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_27
timestamp 1704896540
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_29
timestamp 1704896540
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_41
timestamp 1704896540
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_53
timestamp 1704896540
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_65
timestamp 1704896540
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_77
timestamp 1704896540
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_83
timestamp 1704896540
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_85
timestamp 1704896540
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_97
timestamp 1704896540
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_109
timestamp 1704896540
transform 1 0 11132 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_121
timestamp 1704896540
transform 1 0 12236 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_133
timestamp 1704896540
transform 1 0 13340 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_139
timestamp 1704896540
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_141
timestamp 1704896540
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_153
timestamp 1704896540
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_165
timestamp 1704896540
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_177
timestamp 1704896540
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_189
timestamp 1704896540
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_195
timestamp 1704896540
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_197
timestamp 1704896540
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_209
timestamp 1704896540
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_221
timestamp 1704896540
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_233
timestamp 1704896540
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_245
timestamp 1704896540
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_251
timestamp 1704896540
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_253
timestamp 1704896540
transform 1 0 24380 0 1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_271
timestamp 1704896540
transform 1 0 26036 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_283
timestamp 1704896540
transform 1 0 27140 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_295
timestamp 1704896540
transform 1 0 28244 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_307
timestamp 1704896540
transform 1 0 29348 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_309
timestamp 1704896540
transform 1 0 29532 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_321
timestamp 1704896540
transform 1 0 30636 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_333
timestamp 1704896540
transform 1 0 31740 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_88_345
timestamp 1704896540
transform 1 0 32844 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_353
timestamp 1704896540
transform 1 0 33580 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_88_360
timestamp 1704896540
transform 1 0 34224 0 1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_365
timestamp 1704896540
transform 1 0 34684 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_377
timestamp 1704896540
transform 1 0 35788 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_88_389
timestamp 1704896540
transform 1 0 36892 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_88_421
timestamp 1704896540
transform 1 0 39836 0 1 50048
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_3
timestamp 1704896540
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_15
timestamp 1704896540
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_27
timestamp 1704896540
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_39
timestamp 1704896540
transform 1 0 4692 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_89_51
timestamp 1704896540
transform 1 0 5796 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_55
timestamp 1704896540
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_57
timestamp 1704896540
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_69
timestamp 1704896540
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_81
timestamp 1704896540
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_93
timestamp 1704896540
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_105
timestamp 1704896540
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_111
timestamp 1704896540
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_113
timestamp 1704896540
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_89_125
timestamp 1704896540
transform 1 0 12604 0 -1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_131
timestamp 1704896540
transform 1 0 13156 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_143
timestamp 1704896540
transform 1 0 14260 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_155
timestamp 1704896540
transform 1 0 15364 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_167
timestamp 1704896540
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_169
timestamp 1704896540
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_181
timestamp 1704896540
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_193
timestamp 1704896540
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_205
timestamp 1704896540
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_217
timestamp 1704896540
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_223
timestamp 1704896540
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_225
timestamp 1704896540
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_237
timestamp 1704896540
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_249
timestamp 1704896540
transform 1 0 24012 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_261
timestamp 1704896540
transform 1 0 25116 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_273
timestamp 1704896540
transform 1 0 26220 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_279
timestamp 1704896540
transform 1 0 26772 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_281
timestamp 1704896540
transform 1 0 26956 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_293
timestamp 1704896540
transform 1 0 28060 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_305
timestamp 1704896540
transform 1 0 29164 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_317
timestamp 1704896540
transform 1 0 30268 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_329
timestamp 1704896540
transform 1 0 31372 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_335
timestamp 1704896540
transform 1 0 31924 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_337
timestamp 1704896540
transform 1 0 32108 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_349
timestamp 1704896540
transform 1 0 33212 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_361
timestamp 1704896540
transform 1 0 34316 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_373
timestamp 1704896540
transform 1 0 35420 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_385
timestamp 1704896540
transform 1 0 36524 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_391
timestamp 1704896540
transform 1 0 37076 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_393
timestamp 1704896540
transform 1 0 37260 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_405
timestamp 1704896540
transform 1 0 38364 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_417
timestamp 1704896540
transform 1 0 39468 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_3
timestamp 1704896540
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_15
timestamp 1704896540
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_27
timestamp 1704896540
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_29
timestamp 1704896540
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_41
timestamp 1704896540
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_53
timestamp 1704896540
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_65
timestamp 1704896540
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_77
timestamp 1704896540
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_83
timestamp 1704896540
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_85
timestamp 1704896540
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_90_97
timestamp 1704896540
transform 1 0 10028 0 1 51136
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_114
timestamp 1704896540
transform 1 0 11592 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_126
timestamp 1704896540
transform 1 0 12696 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_90_138
timestamp 1704896540
transform 1 0 13800 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_141
timestamp 1704896540
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_153
timestamp 1704896540
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_90_165
timestamp 1704896540
transform 1 0 16284 0 1 51136
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_176
timestamp 1704896540
transform 1 0 17296 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_90_188
timestamp 1704896540
transform 1 0 18400 0 1 51136
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_197
timestamp 1704896540
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_209
timestamp 1704896540
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_221
timestamp 1704896540
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_233
timestamp 1704896540
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_245
timestamp 1704896540
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_251
timestamp 1704896540
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_253
timestamp 1704896540
transform 1 0 24380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_265
timestamp 1704896540
transform 1 0 25484 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_277
timestamp 1704896540
transform 1 0 26588 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_289
timestamp 1704896540
transform 1 0 27692 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_301
timestamp 1704896540
transform 1 0 28796 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_307
timestamp 1704896540
transform 1 0 29348 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_309
timestamp 1704896540
transform 1 0 29532 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_321
timestamp 1704896540
transform 1 0 30636 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_333
timestamp 1704896540
transform 1 0 31740 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_90_345
timestamp 1704896540
transform 1 0 32844 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_349
timestamp 1704896540
transform 1 0 33212 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_90_361
timestamp 1704896540
transform 1 0 34316 0 1 51136
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_365
timestamp 1704896540
transform 1 0 34684 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_377
timestamp 1704896540
transform 1 0 35788 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_389
timestamp 1704896540
transform 1 0 36892 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_401
timestamp 1704896540
transform 1 0 37996 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_413
timestamp 1704896540
transform 1 0 39100 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_419
timestamp 1704896540
transform 1 0 39652 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_90_421
timestamp 1704896540
transform 1 0 39836 0 1 51136
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_3
timestamp 1704896540
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_15
timestamp 1704896540
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_27
timestamp 1704896540
transform 1 0 3588 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_33
timestamp 1704896540
transform 1 0 4140 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_36
timestamp 1704896540
transform 1 0 4416 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_91_48
timestamp 1704896540
transform 1 0 5520 0 -1 52224
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_57
timestamp 1704896540
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_69
timestamp 1704896540
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_81
timestamp 1704896540
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_91_93
timestamp 1704896540
transform 1 0 9660 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_105
timestamp 1704896540
transform 1 0 10764 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_111
timestamp 1704896540
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_113
timestamp 1704896540
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_125
timestamp 1704896540
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_137
timestamp 1704896540
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_149
timestamp 1704896540
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_161
timestamp 1704896540
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_167
timestamp 1704896540
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_169
timestamp 1704896540
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_181
timestamp 1704896540
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_193
timestamp 1704896540
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_205
timestamp 1704896540
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_217
timestamp 1704896540
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_223
timestamp 1704896540
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_225
timestamp 1704896540
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_237
timestamp 1704896540
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_249
timestamp 1704896540
transform 1 0 24012 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_261
timestamp 1704896540
transform 1 0 25116 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_273
timestamp 1704896540
transform 1 0 26220 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_279
timestamp 1704896540
transform 1 0 26772 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_281
timestamp 1704896540
transform 1 0 26956 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_293
timestamp 1704896540
transform 1 0 28060 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_305
timestamp 1704896540
transform 1 0 29164 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_91_317
timestamp 1704896540
transform 1 0 30268 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_91_325
timestamp 1704896540
transform 1 0 31004 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_335
timestamp 1704896540
transform 1 0 31924 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_91_337
timestamp 1704896540
transform 1 0 32108 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_91_345
timestamp 1704896540
transform 1 0 32844 0 -1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_351
timestamp 1704896540
transform 1 0 33396 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_363
timestamp 1704896540
transform 1 0 34500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_375
timestamp 1704896540
transform 1 0 35604 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_91_387
timestamp 1704896540
transform 1 0 36708 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_391
timestamp 1704896540
transform 1 0 37076 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_393
timestamp 1704896540
transform 1 0 37260 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_405
timestamp 1704896540
transform 1 0 38364 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_417
timestamp 1704896540
transform 1 0 39468 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_3
timestamp 1704896540
transform 1 0 1380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_15
timestamp 1704896540
transform 1 0 2484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_27
timestamp 1704896540
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_92_29
timestamp 1704896540
transform 1 0 3772 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_33
timestamp 1704896540
transform 1 0 4140 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_92_36
timestamp 1704896540
transform 1 0 4416 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_92_40
timestamp 1704896540
transform 1 0 4784 0 1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_50
timestamp 1704896540
transform 1 0 5704 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_62
timestamp 1704896540
transform 1 0 6808 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_92_74
timestamp 1704896540
transform 1 0 7912 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_92_82
timestamp 1704896540
transform 1 0 8648 0 1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_85
timestamp 1704896540
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_97
timestamp 1704896540
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_109
timestamp 1704896540
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_121
timestamp 1704896540
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_133
timestamp 1704896540
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_139
timestamp 1704896540
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_141
timestamp 1704896540
transform 1 0 14076 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_153
timestamp 1704896540
transform 1 0 15180 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_165
timestamp 1704896540
transform 1 0 16284 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_177
timestamp 1704896540
transform 1 0 17388 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_189
timestamp 1704896540
transform 1 0 18492 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_195
timestamp 1704896540
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_197
timestamp 1704896540
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_209
timestamp 1704896540
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_221
timestamp 1704896540
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_233
timestamp 1704896540
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_92_245
timestamp 1704896540
transform 1 0 23644 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_251
timestamp 1704896540
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_253
timestamp 1704896540
transform 1 0 24380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_265
timestamp 1704896540
transform 1 0 25484 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_277
timestamp 1704896540
transform 1 0 26588 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_289
timestamp 1704896540
transform 1 0 27692 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_301
timestamp 1704896540
transform 1 0 28796 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_307
timestamp 1704896540
transform 1 0 29348 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_309
timestamp 1704896540
transform 1 0 29532 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_321
timestamp 1704896540
transform 1 0 30636 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_333
timestamp 1704896540
transform 1 0 31740 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_345
timestamp 1704896540
transform 1 0 32844 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_357
timestamp 1704896540
transform 1 0 33948 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_363
timestamp 1704896540
transform 1 0 34500 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_365
timestamp 1704896540
transform 1 0 34684 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_377
timestamp 1704896540
transform 1 0 35788 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_383
timestamp 1704896540
transform 1 0 36340 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_92_386
timestamp 1704896540
transform 1 0 36616 0 1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_394
timestamp 1704896540
transform 1 0 37352 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_406
timestamp 1704896540
transform 1 0 38456 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_92_418
timestamp 1704896540
transform 1 0 39560 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_92_421
timestamp 1704896540
transform 1 0 39836 0 1 52224
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_3
timestamp 1704896540
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_15
timestamp 1704896540
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_27
timestamp 1704896540
transform 1 0 3588 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_39
timestamp 1704896540
transform 1 0 4692 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_93_51
timestamp 1704896540
transform 1 0 5796 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_55
timestamp 1704896540
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_57
timestamp 1704896540
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_69
timestamp 1704896540
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_81
timestamp 1704896540
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_93
timestamp 1704896540
transform 1 0 9660 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_105
timestamp 1704896540
transform 1 0 10764 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_111
timestamp 1704896540
transform 1 0 11316 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_113
timestamp 1704896540
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_125
timestamp 1704896540
transform 1 0 12604 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_137
timestamp 1704896540
transform 1 0 13708 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_149
timestamp 1704896540
transform 1 0 14812 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_161
timestamp 1704896540
transform 1 0 15916 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_167
timestamp 1704896540
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_169
timestamp 1704896540
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_181
timestamp 1704896540
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_193
timestamp 1704896540
transform 1 0 18860 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_205
timestamp 1704896540
transform 1 0 19964 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_217
timestamp 1704896540
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_223
timestamp 1704896540
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_225
timestamp 1704896540
transform 1 0 21804 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_260
timestamp 1704896540
transform 1 0 25024 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_93_272
timestamp 1704896540
transform 1 0 26128 0 -1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_281
timestamp 1704896540
transform 1 0 26956 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_293
timestamp 1704896540
transform 1 0 28060 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_305
timestamp 1704896540
transform 1 0 29164 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_317
timestamp 1704896540
transform 1 0 30268 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_329
timestamp 1704896540
transform 1 0 31372 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_335
timestamp 1704896540
transform 1 0 31924 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_337
timestamp 1704896540
transform 1 0 32108 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_349
timestamp 1704896540
transform 1 0 33212 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_361
timestamp 1704896540
transform 1 0 34316 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_373
timestamp 1704896540
transform 1 0 35420 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_385
timestamp 1704896540
transform 1 0 36524 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_391
timestamp 1704896540
transform 1 0 37076 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_393
timestamp 1704896540
transform 1 0 37260 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_405
timestamp 1704896540
transform 1 0 38364 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_417
timestamp 1704896540
transform 1 0 39468 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_3
timestamp 1704896540
transform 1 0 1380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_15
timestamp 1704896540
transform 1 0 2484 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_27
timestamp 1704896540
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_29
timestamp 1704896540
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_41
timestamp 1704896540
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_53
timestamp 1704896540
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_65
timestamp 1704896540
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_77
timestamp 1704896540
transform 1 0 8188 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_83
timestamp 1704896540
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_85
timestamp 1704896540
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_97
timestamp 1704896540
transform 1 0 10028 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_109
timestamp 1704896540
transform 1 0 11132 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_94_121
timestamp 1704896540
transform 1 0 12236 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_94_127
timestamp 1704896540
transform 1 0 12788 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_139
timestamp 1704896540
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_141
timestamp 1704896540
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_153
timestamp 1704896540
transform 1 0 15180 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_165
timestamp 1704896540
transform 1 0 16284 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_177
timestamp 1704896540
transform 1 0 17388 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_189
timestamp 1704896540
transform 1 0 18492 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_195
timestamp 1704896540
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_197
timestamp 1704896540
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_209
timestamp 1704896540
transform 1 0 20332 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_221
timestamp 1704896540
transform 1 0 21436 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_233
timestamp 1704896540
transform 1 0 22540 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_245
timestamp 1704896540
transform 1 0 23644 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_251
timestamp 1704896540
transform 1 0 24196 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_253
timestamp 1704896540
transform 1 0 24380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_265
timestamp 1704896540
transform 1 0 25484 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_277
timestamp 1704896540
transform 1 0 26588 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_289
timestamp 1704896540
transform 1 0 27692 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_301
timestamp 1704896540
transform 1 0 28796 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_307
timestamp 1704896540
transform 1 0 29348 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_309
timestamp 1704896540
transform 1 0 29532 0 1 53312
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_338
timestamp 1704896540
transform 1 0 32200 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_350
timestamp 1704896540
transform 1 0 33304 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_94_362
timestamp 1704896540
transform 1 0 34408 0 1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_365
timestamp 1704896540
transform 1 0 34684 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_398
timestamp 1704896540
transform 1 0 37720 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_94_410
timestamp 1704896540
transform 1 0 38824 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_94_418
timestamp 1704896540
transform 1 0 39560 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_94_421
timestamp 1704896540
transform 1 0 39836 0 1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_3
timestamp 1704896540
transform 1 0 1380 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_15
timestamp 1704896540
transform 1 0 2484 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_27
timestamp 1704896540
transform 1 0 3588 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_39
timestamp 1704896540
transform 1 0 4692 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_95_51
timestamp 1704896540
transform 1 0 5796 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_55
timestamp 1704896540
transform 1 0 6164 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_57
timestamp 1704896540
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_95_69
timestamp 1704896540
transform 1 0 7452 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_95_77
timestamp 1704896540
transform 1 0 8188 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_95_102
timestamp 1704896540
transform 1 0 10488 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_95_110
timestamp 1704896540
transform 1 0 11224 0 -1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_113
timestamp 1704896540
transform 1 0 11500 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_125
timestamp 1704896540
transform 1 0 12604 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_137
timestamp 1704896540
transform 1 0 13708 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_149
timestamp 1704896540
transform 1 0 14812 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_161
timestamp 1704896540
transform 1 0 15916 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_167
timestamp 1704896540
transform 1 0 16468 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_169
timestamp 1704896540
transform 1 0 16652 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_175
timestamp 1704896540
transform 1 0 17204 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_183
timestamp 1704896540
transform 1 0 17940 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_195
timestamp 1704896540
transform 1 0 19044 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_207
timestamp 1704896540
transform 1 0 20148 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_95_219
timestamp 1704896540
transform 1 0 21252 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_223
timestamp 1704896540
transform 1 0 21620 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_225
timestamp 1704896540
transform 1 0 21804 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_237
timestamp 1704896540
transform 1 0 22908 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_249
timestamp 1704896540
transform 1 0 24012 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_261
timestamp 1704896540
transform 1 0 25116 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_273
timestamp 1704896540
transform 1 0 26220 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_279
timestamp 1704896540
transform 1 0 26772 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_281
timestamp 1704896540
transform 1 0 26956 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_293
timestamp 1704896540
transform 1 0 28060 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_305
timestamp 1704896540
transform 1 0 29164 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_317
timestamp 1704896540
transform 1 0 30268 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_329
timestamp 1704896540
transform 1 0 31372 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_335
timestamp 1704896540
transform 1 0 31924 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_337
timestamp 1704896540
transform 1 0 32108 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_349
timestamp 1704896540
transform 1 0 33212 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_361
timestamp 1704896540
transform 1 0 34316 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_373
timestamp 1704896540
transform 1 0 35420 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_385
timestamp 1704896540
transform 1 0 36524 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_391
timestamp 1704896540
transform 1 0 37076 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_393
timestamp 1704896540
transform 1 0 37260 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_405
timestamp 1704896540
transform 1 0 38364 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_417
timestamp 1704896540
transform 1 0 39468 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_3
timestamp 1704896540
transform 1 0 1380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_15
timestamp 1704896540
transform 1 0 2484 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_27
timestamp 1704896540
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_29
timestamp 1704896540
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_41
timestamp 1704896540
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_53
timestamp 1704896540
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_65
timestamp 1704896540
transform 1 0 7084 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_77
timestamp 1704896540
transform 1 0 8188 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_83
timestamp 1704896540
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_85
timestamp 1704896540
transform 1 0 8924 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_97
timestamp 1704896540
transform 1 0 10028 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_109
timestamp 1704896540
transform 1 0 11132 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_121
timestamp 1704896540
transform 1 0 12236 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_133
timestamp 1704896540
transform 1 0 13340 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_139
timestamp 1704896540
transform 1 0 13892 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_141
timestamp 1704896540
transform 1 0 14076 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_153
timestamp 1704896540
transform 1 0 15180 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_165
timestamp 1704896540
transform 1 0 16284 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_177
timestamp 1704896540
transform 1 0 17388 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_189
timestamp 1704896540
transform 1 0 18492 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_195
timestamp 1704896540
transform 1 0 19044 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_197
timestamp 1704896540
transform 1 0 19228 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_209
timestamp 1704896540
transform 1 0 20332 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_221
timestamp 1704896540
transform 1 0 21436 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_233
timestamp 1704896540
transform 1 0 22540 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_245
timestamp 1704896540
transform 1 0 23644 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_251
timestamp 1704896540
transform 1 0 24196 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_253
timestamp 1704896540
transform 1 0 24380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_265
timestamp 1704896540
transform 1 0 25484 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_277
timestamp 1704896540
transform 1 0 26588 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_289
timestamp 1704896540
transform 1 0 27692 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_301
timestamp 1704896540
transform 1 0 28796 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_307
timestamp 1704896540
transform 1 0 29348 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_309
timestamp 1704896540
transform 1 0 29532 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_321
timestamp 1704896540
transform 1 0 30636 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_333
timestamp 1704896540
transform 1 0 31740 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_345
timestamp 1704896540
transform 1 0 32844 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_357
timestamp 1704896540
transform 1 0 33948 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_363
timestamp 1704896540
transform 1 0 34500 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_365
timestamp 1704896540
transform 1 0 34684 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_377
timestamp 1704896540
transform 1 0 35788 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_389
timestamp 1704896540
transform 1 0 36892 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_401
timestamp 1704896540
transform 1 0 37996 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_96_421
timestamp 1704896540
transform 1 0 39836 0 1 54400
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_3
timestamp 1704896540
transform 1 0 1380 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_15
timestamp 1704896540
transform 1 0 2484 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_27
timestamp 1704896540
transform 1 0 3588 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_39
timestamp 1704896540
transform 1 0 4692 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_97_51
timestamp 1704896540
transform 1 0 5796 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_55
timestamp 1704896540
transform 1 0 6164 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_57
timestamp 1704896540
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_69
timestamp 1704896540
transform 1 0 7452 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_81
timestamp 1704896540
transform 1 0 8556 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_93
timestamp 1704896540
transform 1 0 9660 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_105
timestamp 1704896540
transform 1 0 10764 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_111
timestamp 1704896540
transform 1 0 11316 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_113
timestamp 1704896540
transform 1 0 11500 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_125
timestamp 1704896540
transform 1 0 12604 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_137
timestamp 1704896540
transform 1 0 13708 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_149
timestamp 1704896540
transform 1 0 14812 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_161
timestamp 1704896540
transform 1 0 15916 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_167
timestamp 1704896540
transform 1 0 16468 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_169
timestamp 1704896540
transform 1 0 16652 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_181
timestamp 1704896540
transform 1 0 17756 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_193
timestamp 1704896540
transform 1 0 18860 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_205
timestamp 1704896540
transform 1 0 19964 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_97_214
timestamp 1704896540
transform 1 0 20792 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_97_222
timestamp 1704896540
transform 1 0 21528 0 -1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_225
timestamp 1704896540
transform 1 0 21804 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_237
timestamp 1704896540
transform 1 0 22908 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_249
timestamp 1704896540
transform 1 0 24012 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_261
timestamp 1704896540
transform 1 0 25116 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_273
timestamp 1704896540
transform 1 0 26220 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_279
timestamp 1704896540
transform 1 0 26772 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_281
timestamp 1704896540
transform 1 0 26956 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_293
timestamp 1704896540
transform 1 0 28060 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_305
timestamp 1704896540
transform 1 0 29164 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_317
timestamp 1704896540
transform 1 0 30268 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_321
timestamp 1704896540
transform 1 0 30636 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_97_333
timestamp 1704896540
transform 1 0 31740 0 -1 55488
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_337
timestamp 1704896540
transform 1 0 32108 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_349
timestamp 1704896540
transform 1 0 33212 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_361
timestamp 1704896540
transform 1 0 34316 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_373
timestamp 1704896540
transform 1 0 35420 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_385
timestamp 1704896540
transform 1 0 36524 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_391
timestamp 1704896540
transform 1 0 37076 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_393
timestamp 1704896540
transform 1 0 37260 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_405
timestamp 1704896540
transform 1 0 38364 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_97_417
timestamp 1704896540
transform 1 0 39468 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_423
timestamp 1704896540
transform 1 0 40020 0 -1 55488
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_3
timestamp 1704896540
transform 1 0 1380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_15
timestamp 1704896540
transform 1 0 2484 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_27
timestamp 1704896540
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_29
timestamp 1704896540
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_41
timestamp 1704896540
transform 1 0 4876 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_53
timestamp 1704896540
transform 1 0 5980 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_65
timestamp 1704896540
transform 1 0 7084 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_77
timestamp 1704896540
transform 1 0 8188 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_83
timestamp 1704896540
transform 1 0 8740 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_85
timestamp 1704896540
transform 1 0 8924 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_97
timestamp 1704896540
transform 1 0 10028 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_109
timestamp 1704896540
transform 1 0 11132 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_121
timestamp 1704896540
transform 1 0 12236 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_133
timestamp 1704896540
transform 1 0 13340 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_139
timestamp 1704896540
transform 1 0 13892 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_141
timestamp 1704896540
transform 1 0 14076 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_153
timestamp 1704896540
transform 1 0 15180 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_165
timestamp 1704896540
transform 1 0 16284 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_177
timestamp 1704896540
transform 1 0 17388 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_189
timestamp 1704896540
transform 1 0 18492 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_195
timestamp 1704896540
transform 1 0 19044 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_197
timestamp 1704896540
transform 1 0 19228 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_209
timestamp 1704896540
transform 1 0 20332 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_221
timestamp 1704896540
transform 1 0 21436 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_233
timestamp 1704896540
transform 1 0 22540 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_245
timestamp 1704896540
transform 1 0 23644 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_251
timestamp 1704896540
transform 1 0 24196 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_253
timestamp 1704896540
transform 1 0 24380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_265
timestamp 1704896540
transform 1 0 25484 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_277
timestamp 1704896540
transform 1 0 26588 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_289
timestamp 1704896540
transform 1 0 27692 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_98_303
timestamp 1704896540
transform 1 0 28980 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_307
timestamp 1704896540
transform 1 0 29348 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_312
timestamp 1704896540
transform 1 0 29808 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_324
timestamp 1704896540
transform 1 0 30912 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_336
timestamp 1704896540
transform 1 0 32016 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_348
timestamp 1704896540
transform 1 0 33120 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_98_360
timestamp 1704896540
transform 1 0 34224 0 1 55488
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_365
timestamp 1704896540
transform 1 0 34684 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_377
timestamp 1704896540
transform 1 0 35788 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_389
timestamp 1704896540
transform 1 0 36892 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_401
timestamp 1704896540
transform 1 0 37996 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_413
timestamp 1704896540
transform 1 0 39100 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_419
timestamp 1704896540
transform 1 0 39652 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_98_421
timestamp 1704896540
transform 1 0 39836 0 1 55488
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_3
timestamp 1704896540
transform 1 0 1380 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_15
timestamp 1704896540
transform 1 0 2484 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_27
timestamp 1704896540
transform 1 0 3588 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_39
timestamp 1704896540
transform 1 0 4692 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_99_51
timestamp 1704896540
transform 1 0 5796 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_55
timestamp 1704896540
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_57
timestamp 1704896540
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_69
timestamp 1704896540
transform 1 0 7452 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_81
timestamp 1704896540
transform 1 0 8556 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_93
timestamp 1704896540
transform 1 0 9660 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_105
timestamp 1704896540
transform 1 0 10764 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_111
timestamp 1704896540
transform 1 0 11316 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_113
timestamp 1704896540
transform 1 0 11500 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_125
timestamp 1704896540
transform 1 0 12604 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_137
timestamp 1704896540
transform 1 0 13708 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_149
timestamp 1704896540
transform 1 0 14812 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_161
timestamp 1704896540
transform 1 0 15916 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_167
timestamp 1704896540
transform 1 0 16468 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_169
timestamp 1704896540
transform 1 0 16652 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_181
timestamp 1704896540
transform 1 0 17756 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_193
timestamp 1704896540
transform 1 0 18860 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_205
timestamp 1704896540
transform 1 0 19964 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_217
timestamp 1704896540
transform 1 0 21068 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_223
timestamp 1704896540
transform 1 0 21620 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_225
timestamp 1704896540
transform 1 0 21804 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_237
timestamp 1704896540
transform 1 0 22908 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_249
timestamp 1704896540
transform 1 0 24012 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_261
timestamp 1704896540
transform 1 0 25116 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_273
timestamp 1704896540
transform 1 0 26220 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_279
timestamp 1704896540
transform 1 0 26772 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_281
timestamp 1704896540
transform 1 0 26956 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_99_293
timestamp 1704896540
transform 1 0 28060 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_99_299
timestamp 1704896540
transform 1 0 28612 0 -1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_307
timestamp 1704896540
transform 1 0 29348 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_319
timestamp 1704896540
transform 1 0 30452 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_99_331
timestamp 1704896540
transform 1 0 31556 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_335
timestamp 1704896540
transform 1 0 31924 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_337
timestamp 1704896540
transform 1 0 32108 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_99_349
timestamp 1704896540
transform 1 0 33212 0 -1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_357
timestamp 1704896540
transform 1 0 33948 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_369
timestamp 1704896540
transform 1 0 35052 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_99_381
timestamp 1704896540
transform 1 0 36156 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_99_389
timestamp 1704896540
transform 1 0 36892 0 -1 56576
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_416
timestamp 1704896540
transform 1 0 39376 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_428
timestamp 1704896540
transform 1 0 40480 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_3
timestamp 1704896540
transform 1 0 1380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_15
timestamp 1704896540
transform 1 0 2484 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_27
timestamp 1704896540
transform 1 0 3588 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_29
timestamp 1704896540
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_41
timestamp 1704896540
transform 1 0 4876 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_100_76
timestamp 1704896540
transform 1 0 8096 0 1 56576
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_85
timestamp 1704896540
transform 1 0 8924 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_97
timestamp 1704896540
transform 1 0 10028 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_109
timestamp 1704896540
transform 1 0 11132 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_121
timestamp 1704896540
transform 1 0 12236 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_133
timestamp 1704896540
transform 1 0 13340 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_139
timestamp 1704896540
transform 1 0 13892 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_141
timestamp 1704896540
transform 1 0 14076 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_153
timestamp 1704896540
transform 1 0 15180 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_165
timestamp 1704896540
transform 1 0 16284 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_177
timestamp 1704896540
transform 1 0 17388 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_189
timestamp 1704896540
transform 1 0 18492 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_195
timestamp 1704896540
transform 1 0 19044 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_197
timestamp 1704896540
transform 1 0 19228 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_209
timestamp 1704896540
transform 1 0 20332 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_221
timestamp 1704896540
transform 1 0 21436 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_233
timestamp 1704896540
transform 1 0 22540 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_245
timestamp 1704896540
transform 1 0 23644 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_251
timestamp 1704896540
transform 1 0 24196 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_253
timestamp 1704896540
transform 1 0 24380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_265
timestamp 1704896540
transform 1 0 25484 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_277
timestamp 1704896540
transform 1 0 26588 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_289
timestamp 1704896540
transform 1 0 27692 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_301
timestamp 1704896540
transform 1 0 28796 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_307
timestamp 1704896540
transform 1 0 29348 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_309
timestamp 1704896540
transform 1 0 29532 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_321
timestamp 1704896540
transform 1 0 30636 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_333
timestamp 1704896540
transform 1 0 31740 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_345
timestamp 1704896540
transform 1 0 32844 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_357
timestamp 1704896540
transform 1 0 33948 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_363
timestamp 1704896540
transform 1 0 34500 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_365
timestamp 1704896540
transform 1 0 34684 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_377
timestamp 1704896540
transform 1 0 35788 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_389
timestamp 1704896540
transform 1 0 36892 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_401
timestamp 1704896540
transform 1 0 37996 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_413
timestamp 1704896540
transform 1 0 39100 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_419
timestamp 1704896540
transform 1 0 39652 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_100_421
timestamp 1704896540
transform 1 0 39836 0 1 56576
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_3
timestamp 1704896540
transform 1 0 1380 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_101_15
timestamp 1704896540
transform 1 0 2484 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_55
timestamp 1704896540
transform 1 0 6164 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_57
timestamp 1704896540
transform 1 0 6348 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_69
timestamp 1704896540
transform 1 0 7452 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_81
timestamp 1704896540
transform 1 0 8556 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_93
timestamp 1704896540
transform 1 0 9660 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_105
timestamp 1704896540
transform 1 0 10764 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_111
timestamp 1704896540
transform 1 0 11316 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_113
timestamp 1704896540
transform 1 0 11500 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_125
timestamp 1704896540
transform 1 0 12604 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_137
timestamp 1704896540
transform 1 0 13708 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_149
timestamp 1704896540
transform 1 0 14812 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_161
timestamp 1704896540
transform 1 0 15916 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_167
timestamp 1704896540
transform 1 0 16468 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_169
timestamp 1704896540
transform 1 0 16652 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_181
timestamp 1704896540
transform 1 0 17756 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_193
timestamp 1704896540
transform 1 0 18860 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_205
timestamp 1704896540
transform 1 0 19964 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_217
timestamp 1704896540
transform 1 0 21068 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_223
timestamp 1704896540
transform 1 0 21620 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_225
timestamp 1704896540
transform 1 0 21804 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_237
timestamp 1704896540
transform 1 0 22908 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_249
timestamp 1704896540
transform 1 0 24012 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_261
timestamp 1704896540
transform 1 0 25116 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_273
timestamp 1704896540
transform 1 0 26220 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_279
timestamp 1704896540
transform 1 0 26772 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_281
timestamp 1704896540
transform 1 0 26956 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_293
timestamp 1704896540
transform 1 0 28060 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101_305
timestamp 1704896540
transform 1 0 29164 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_309
timestamp 1704896540
transform 1 0 29532 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_319
timestamp 1704896540
transform 1 0 30452 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101_331
timestamp 1704896540
transform 1 0 31556 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_335
timestamp 1704896540
transform 1 0 31924 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_337
timestamp 1704896540
transform 1 0 32108 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_101_349
timestamp 1704896540
transform 1 0 33212 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_101_357
timestamp 1704896540
transform 1 0 33948 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_385
timestamp 1704896540
transform 1 0 36524 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_391
timestamp 1704896540
transform 1 0 37076 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_393
timestamp 1704896540
transform 1 0 37260 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_405
timestamp 1704896540
transform 1 0 38364 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_417
timestamp 1704896540
transform 1 0 39468 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_3
timestamp 1704896540
transform 1 0 1380 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_15
timestamp 1704896540
transform 1 0 2484 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_27
timestamp 1704896540
transform 1 0 3588 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_29
timestamp 1704896540
transform 1 0 3772 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_41
timestamp 1704896540
transform 1 0 4876 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_53
timestamp 1704896540
transform 1 0 5980 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_65
timestamp 1704896540
transform 1 0 7084 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_102_77
timestamp 1704896540
transform 1 0 8188 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_83
timestamp 1704896540
transform 1 0 8740 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_85
timestamp 1704896540
transform 1 0 8924 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_97
timestamp 1704896540
transform 1 0 10028 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_109
timestamp 1704896540
transform 1 0 11132 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_121
timestamp 1704896540
transform 1 0 12236 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_102_133
timestamp 1704896540
transform 1 0 13340 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_139
timestamp 1704896540
transform 1 0 13892 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_141
timestamp 1704896540
transform 1 0 14076 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_153
timestamp 1704896540
transform 1 0 15180 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_165
timestamp 1704896540
transform 1 0 16284 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_177
timestamp 1704896540
transform 1 0 17388 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_102_189
timestamp 1704896540
transform 1 0 18492 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_195
timestamp 1704896540
transform 1 0 19044 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_197
timestamp 1704896540
transform 1 0 19228 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_209
timestamp 1704896540
transform 1 0 20332 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_221
timestamp 1704896540
transform 1 0 21436 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_233
timestamp 1704896540
transform 1 0 22540 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_102_245
timestamp 1704896540
transform 1 0 23644 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_251
timestamp 1704896540
transform 1 0 24196 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_253
timestamp 1704896540
transform 1 0 24380 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_265
timestamp 1704896540
transform 1 0 25484 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_277
timestamp 1704896540
transform 1 0 26588 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_289
timestamp 1704896540
transform 1 0 27692 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_102_301
timestamp 1704896540
transform 1 0 28796 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_307
timestamp 1704896540
transform 1 0 29348 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_309
timestamp 1704896540
transform 1 0 29532 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_321
timestamp 1704896540
transform 1 0 30636 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_333
timestamp 1704896540
transform 1 0 31740 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_345
timestamp 1704896540
transform 1 0 32844 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_102_357
timestamp 1704896540
transform 1 0 33948 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_363
timestamp 1704896540
transform 1 0 34500 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_365
timestamp 1704896540
transform 1 0 34684 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_377
timestamp 1704896540
transform 1 0 35788 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_389
timestamp 1704896540
transform 1 0 36892 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_401
timestamp 1704896540
transform 1 0 37996 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_102_413
timestamp 1704896540
transform 1 0 39100 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_419
timestamp 1704896540
transform 1 0 39652 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_102_425
timestamp 1704896540
transform 1 0 40204 0 1 57664
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_3
timestamp 1704896540
transform 1 0 1380 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_15
timestamp 1704896540
transform 1 0 2484 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_27
timestamp 1704896540
transform 1 0 3588 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_39
timestamp 1704896540
transform 1 0 4692 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_103_51
timestamp 1704896540
transform 1 0 5796 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_55
timestamp 1704896540
transform 1 0 6164 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_57
timestamp 1704896540
transform 1 0 6348 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_69
timestamp 1704896540
transform 1 0 7452 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_81
timestamp 1704896540
transform 1 0 8556 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_93
timestamp 1704896540
transform 1 0 9660 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_103_105
timestamp 1704896540
transform 1 0 10764 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_111
timestamp 1704896540
transform 1 0 11316 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_113
timestamp 1704896540
transform 1 0 11500 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_125
timestamp 1704896540
transform 1 0 12604 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_137
timestamp 1704896540
transform 1 0 13708 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_149
timestamp 1704896540
transform 1 0 14812 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_103_161
timestamp 1704896540
transform 1 0 15916 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_167
timestamp 1704896540
transform 1 0 16468 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_169
timestamp 1704896540
transform 1 0 16652 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_181
timestamp 1704896540
transform 1 0 17756 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_193
timestamp 1704896540
transform 1 0 18860 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_205
timestamp 1704896540
transform 1 0 19964 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_103_217
timestamp 1704896540
transform 1 0 21068 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_223
timestamp 1704896540
transform 1 0 21620 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_225
timestamp 1704896540
transform 1 0 21804 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_237
timestamp 1704896540
transform 1 0 22908 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_249
timestamp 1704896540
transform 1 0 24012 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_261
timestamp 1704896540
transform 1 0 25116 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_103_273
timestamp 1704896540
transform 1 0 26220 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_279
timestamp 1704896540
transform 1 0 26772 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_281
timestamp 1704896540
transform 1 0 26956 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_293
timestamp 1704896540
transform 1 0 28060 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_305
timestamp 1704896540
transform 1 0 29164 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_317
timestamp 1704896540
transform 1 0 30268 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_103_329
timestamp 1704896540
transform 1 0 31372 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_335
timestamp 1704896540
transform 1 0 31924 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_337
timestamp 1704896540
transform 1 0 32108 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_349
timestamp 1704896540
transform 1 0 33212 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_361
timestamp 1704896540
transform 1 0 34316 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_373
timestamp 1704896540
transform 1 0 35420 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_103_385
timestamp 1704896540
transform 1 0 36524 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_391
timestamp 1704896540
transform 1 0 37076 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_393
timestamp 1704896540
transform 1 0 37260 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_103_405
timestamp 1704896540
transform 1 0 38364 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_103_422
timestamp 1704896540
transform 1 0 39928 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_428
timestamp 1704896540
transform 1 0 40480 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_3
timestamp 1704896540
transform 1 0 1380 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_15
timestamp 1704896540
transform 1 0 2484 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_27
timestamp 1704896540
transform 1 0 3588 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_29
timestamp 1704896540
transform 1 0 3772 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_41
timestamp 1704896540
transform 1 0 4876 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_53
timestamp 1704896540
transform 1 0 5980 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_104_65
timestamp 1704896540
transform 1 0 7084 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_69
timestamp 1704896540
transform 1 0 7452 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_104_73
timestamp 1704896540
transform 1 0 7820 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_104_81
timestamp 1704896540
transform 1 0 8556 0 1 58752
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_85
timestamp 1704896540
transform 1 0 8924 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_97
timestamp 1704896540
transform 1 0 10028 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_109
timestamp 1704896540
transform 1 0 11132 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_121
timestamp 1704896540
transform 1 0 12236 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_104_133
timestamp 1704896540
transform 1 0 13340 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_139
timestamp 1704896540
transform 1 0 13892 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_141
timestamp 1704896540
transform 1 0 14076 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_153
timestamp 1704896540
transform 1 0 15180 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_165
timestamp 1704896540
transform 1 0 16284 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_177
timestamp 1704896540
transform 1 0 17388 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_104_189
timestamp 1704896540
transform 1 0 18492 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_195
timestamp 1704896540
transform 1 0 19044 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_197
timestamp 1704896540
transform 1 0 19228 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_209
timestamp 1704896540
transform 1 0 20332 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_221
timestamp 1704896540
transform 1 0 21436 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_233
timestamp 1704896540
transform 1 0 22540 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_104_245
timestamp 1704896540
transform 1 0 23644 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_251
timestamp 1704896540
transform 1 0 24196 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_253
timestamp 1704896540
transform 1 0 24380 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_265
timestamp 1704896540
transform 1 0 25484 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_277
timestamp 1704896540
transform 1 0 26588 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_289
timestamp 1704896540
transform 1 0 27692 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_104_301
timestamp 1704896540
transform 1 0 28796 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_307
timestamp 1704896540
transform 1 0 29348 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_309
timestamp 1704896540
transform 1 0 29532 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_321
timestamp 1704896540
transform 1 0 30636 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_333
timestamp 1704896540
transform 1 0 31740 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_345
timestamp 1704896540
transform 1 0 32844 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_104_357
timestamp 1704896540
transform 1 0 33948 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_363
timestamp 1704896540
transform 1 0 34500 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_365
timestamp 1704896540
transform 1 0 34684 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_377
timestamp 1704896540
transform 1 0 35788 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_389
timestamp 1704896540
transform 1 0 36892 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_401
timestamp 1704896540
transform 1 0 37996 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_104_413
timestamp 1704896540
transform 1 0 39100 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_419
timestamp 1704896540
transform 1 0 39652 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_104_421
timestamp 1704896540
transform 1 0 39836 0 1 58752
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_3
timestamp 1704896540
transform 1 0 1380 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_15
timestamp 1704896540
transform 1 0 2484 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_27
timestamp 1704896540
transform 1 0 3588 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_39
timestamp 1704896540
transform 1 0 4692 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_105_51
timestamp 1704896540
transform 1 0 5796 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_55
timestamp 1704896540
transform 1 0 6164 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_57
timestamp 1704896540
transform 1 0 6348 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_69
timestamp 1704896540
transform 1 0 7452 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_81
timestamp 1704896540
transform 1 0 8556 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_93
timestamp 1704896540
transform 1 0 9660 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105_105
timestamp 1704896540
transform 1 0 10764 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_111
timestamp 1704896540
transform 1 0 11316 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_113
timestamp 1704896540
transform 1 0 11500 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_125
timestamp 1704896540
transform 1 0 12604 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_137
timestamp 1704896540
transform 1 0 13708 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_149
timestamp 1704896540
transform 1 0 14812 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105_161
timestamp 1704896540
transform 1 0 15916 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_167
timestamp 1704896540
transform 1 0 16468 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_169
timestamp 1704896540
transform 1 0 16652 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_181
timestamp 1704896540
transform 1 0 17756 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_193
timestamp 1704896540
transform 1 0 18860 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_205
timestamp 1704896540
transform 1 0 19964 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105_217
timestamp 1704896540
transform 1 0 21068 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_223
timestamp 1704896540
transform 1 0 21620 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_225
timestamp 1704896540
transform 1 0 21804 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_237
timestamp 1704896540
transform 1 0 22908 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_249
timestamp 1704896540
transform 1 0 24012 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_261
timestamp 1704896540
transform 1 0 25116 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105_273
timestamp 1704896540
transform 1 0 26220 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_279
timestamp 1704896540
transform 1 0 26772 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_281
timestamp 1704896540
transform 1 0 26956 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_293
timestamp 1704896540
transform 1 0 28060 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_305
timestamp 1704896540
transform 1 0 29164 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_317
timestamp 1704896540
transform 1 0 30268 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105_329
timestamp 1704896540
transform 1 0 31372 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_335
timestamp 1704896540
transform 1 0 31924 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_337
timestamp 1704896540
transform 1 0 32108 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_349
timestamp 1704896540
transform 1 0 33212 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_361
timestamp 1704896540
transform 1 0 34316 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_373
timestamp 1704896540
transform 1 0 35420 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105_385
timestamp 1704896540
transform 1 0 36524 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_391
timestamp 1704896540
transform 1 0 37076 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_393
timestamp 1704896540
transform 1 0 37260 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_405
timestamp 1704896540
transform 1 0 38364 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_417
timestamp 1704896540
transform 1 0 39468 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_3
timestamp 1704896540
transform 1 0 1380 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_15
timestamp 1704896540
transform 1 0 2484 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_27
timestamp 1704896540
transform 1 0 3588 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_29
timestamp 1704896540
transform 1 0 3772 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_41
timestamp 1704896540
transform 1 0 4876 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_53
timestamp 1704896540
transform 1 0 5980 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_65
timestamp 1704896540
transform 1 0 7084 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106_77
timestamp 1704896540
transform 1 0 8188 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_83
timestamp 1704896540
transform 1 0 8740 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_85
timestamp 1704896540
transform 1 0 8924 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_97
timestamp 1704896540
transform 1 0 10028 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_109
timestamp 1704896540
transform 1 0 11132 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_121
timestamp 1704896540
transform 1 0 12236 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106_133
timestamp 1704896540
transform 1 0 13340 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_139
timestamp 1704896540
transform 1 0 13892 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_141
timestamp 1704896540
transform 1 0 14076 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_153
timestamp 1704896540
transform 1 0 15180 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_165
timestamp 1704896540
transform 1 0 16284 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_177
timestamp 1704896540
transform 1 0 17388 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106_189
timestamp 1704896540
transform 1 0 18492 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_195
timestamp 1704896540
transform 1 0 19044 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_197
timestamp 1704896540
transform 1 0 19228 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_209
timestamp 1704896540
transform 1 0 20332 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_221
timestamp 1704896540
transform 1 0 21436 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_233
timestamp 1704896540
transform 1 0 22540 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106_245
timestamp 1704896540
transform 1 0 23644 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_251
timestamp 1704896540
transform 1 0 24196 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_106_253
timestamp 1704896540
transform 1 0 24380 0 1 59840
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_259
timestamp 1704896540
transform 1 0 24932 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_271
timestamp 1704896540
transform 1 0 26036 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_283
timestamp 1704896540
transform 1 0 27140 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_295
timestamp 1704896540
transform 1 0 28244 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_307
timestamp 1704896540
transform 1 0 29348 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_309
timestamp 1704896540
transform 1 0 29532 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_321
timestamp 1704896540
transform 1 0 30636 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_333
timestamp 1704896540
transform 1 0 31740 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_345
timestamp 1704896540
transform 1 0 32844 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106_357
timestamp 1704896540
transform 1 0 33948 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_363
timestamp 1704896540
transform 1 0 34500 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_365
timestamp 1704896540
transform 1 0 34684 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_377
timestamp 1704896540
transform 1 0 35788 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_106_389
timestamp 1704896540
transform 1 0 36892 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_397
timestamp 1704896540
transform 1 0 37628 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_403
timestamp 1704896540
transform 1 0 38180 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_106_415
timestamp 1704896540
transform 1 0 39284 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_419
timestamp 1704896540
transform 1 0 39652 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_106_421
timestamp 1704896540
transform 1 0 39836 0 1 59840
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_3
timestamp 1704896540
transform 1 0 1380 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_15
timestamp 1704896540
transform 1 0 2484 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_27
timestamp 1704896540
transform 1 0 3588 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_39
timestamp 1704896540
transform 1 0 4692 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_107_51
timestamp 1704896540
transform 1 0 5796 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_55
timestamp 1704896540
transform 1 0 6164 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_57
timestamp 1704896540
transform 1 0 6348 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_69
timestamp 1704896540
transform 1 0 7452 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_81
timestamp 1704896540
transform 1 0 8556 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_93
timestamp 1704896540
transform 1 0 9660 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_107_105
timestamp 1704896540
transform 1 0 10764 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_111
timestamp 1704896540
transform 1 0 11316 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_113
timestamp 1704896540
transform 1 0 11500 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_125
timestamp 1704896540
transform 1 0 12604 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_137
timestamp 1704896540
transform 1 0 13708 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_149
timestamp 1704896540
transform 1 0 14812 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_107_161
timestamp 1704896540
transform 1 0 15916 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_167
timestamp 1704896540
transform 1 0 16468 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_169
timestamp 1704896540
transform 1 0 16652 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_181
timestamp 1704896540
transform 1 0 17756 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_193
timestamp 1704896540
transform 1 0 18860 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_205
timestamp 1704896540
transform 1 0 19964 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_107_217
timestamp 1704896540
transform 1 0 21068 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_223
timestamp 1704896540
transform 1 0 21620 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_225
timestamp 1704896540
transform 1 0 21804 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_237
timestamp 1704896540
transform 1 0 22908 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_249
timestamp 1704896540
transform 1 0 24012 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_261
timestamp 1704896540
transform 1 0 25116 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_107_273
timestamp 1704896540
transform 1 0 26220 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_279
timestamp 1704896540
transform 1 0 26772 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_281
timestamp 1704896540
transform 1 0 26956 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_293
timestamp 1704896540
transform 1 0 28060 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_305
timestamp 1704896540
transform 1 0 29164 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_317
timestamp 1704896540
transform 1 0 30268 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_107_329
timestamp 1704896540
transform 1 0 31372 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_335
timestamp 1704896540
transform 1 0 31924 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_337
timestamp 1704896540
transform 1 0 32108 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_349
timestamp 1704896540
transform 1 0 33212 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_361
timestamp 1704896540
transform 1 0 34316 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_373
timestamp 1704896540
transform 1 0 35420 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_107_385
timestamp 1704896540
transform 1 0 36524 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_391
timestamp 1704896540
transform 1 0 37076 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_393
timestamp 1704896540
transform 1 0 37260 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_405
timestamp 1704896540
transform 1 0 38364 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_417
timestamp 1704896540
transform 1 0 39468 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_3
timestamp 1704896540
transform 1 0 1380 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_15
timestamp 1704896540
transform 1 0 2484 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_27
timestamp 1704896540
transform 1 0 3588 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_29
timestamp 1704896540
transform 1 0 3772 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_41
timestamp 1704896540
transform 1 0 4876 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_53
timestamp 1704896540
transform 1 0 5980 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_65
timestamp 1704896540
transform 1 0 7084 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_108_77
timestamp 1704896540
transform 1 0 8188 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_83
timestamp 1704896540
transform 1 0 8740 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_85
timestamp 1704896540
transform 1 0 8924 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_97
timestamp 1704896540
transform 1 0 10028 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_109
timestamp 1704896540
transform 1 0 11132 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_121
timestamp 1704896540
transform 1 0 12236 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_108_133
timestamp 1704896540
transform 1 0 13340 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_139
timestamp 1704896540
transform 1 0 13892 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_141
timestamp 1704896540
transform 1 0 14076 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_153
timestamp 1704896540
transform 1 0 15180 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_165
timestamp 1704896540
transform 1 0 16284 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_177
timestamp 1704896540
transform 1 0 17388 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_108_189
timestamp 1704896540
transform 1 0 18492 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_195
timestamp 1704896540
transform 1 0 19044 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_197
timestamp 1704896540
transform 1 0 19228 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_209
timestamp 1704896540
transform 1 0 20332 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_221
timestamp 1704896540
transform 1 0 21436 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_233
timestamp 1704896540
transform 1 0 22540 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_108_245
timestamp 1704896540
transform 1 0 23644 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_251
timestamp 1704896540
transform 1 0 24196 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_253
timestamp 1704896540
transform 1 0 24380 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_265
timestamp 1704896540
transform 1 0 25484 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_277
timestamp 1704896540
transform 1 0 26588 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_289
timestamp 1704896540
transform 1 0 27692 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_108_301
timestamp 1704896540
transform 1 0 28796 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_307
timestamp 1704896540
transform 1 0 29348 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_309
timestamp 1704896540
transform 1 0 29532 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_321
timestamp 1704896540
transform 1 0 30636 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_333
timestamp 1704896540
transform 1 0 31740 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_345
timestamp 1704896540
transform 1 0 32844 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_108_357
timestamp 1704896540
transform 1 0 33948 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_363
timestamp 1704896540
transform 1 0 34500 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_365
timestamp 1704896540
transform 1 0 34684 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_377
timestamp 1704896540
transform 1 0 35788 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_389
timestamp 1704896540
transform 1 0 36892 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_401
timestamp 1704896540
transform 1 0 37996 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_108_413
timestamp 1704896540
transform 1 0 39100 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_419
timestamp 1704896540
transform 1 0 39652 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_108_421
timestamp 1704896540
transform 1 0 39836 0 1 60928
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_3
timestamp 1704896540
transform 1 0 1380 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_15
timestamp 1704896540
transform 1 0 2484 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_27
timestamp 1704896540
transform 1 0 3588 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_39
timestamp 1704896540
transform 1 0 4692 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_109_51
timestamp 1704896540
transform 1 0 5796 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109_55
timestamp 1704896540
transform 1 0 6164 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_57
timestamp 1704896540
transform 1 0 6348 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_69
timestamp 1704896540
transform 1 0 7452 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_81
timestamp 1704896540
transform 1 0 8556 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_93
timestamp 1704896540
transform 1 0 9660 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_109_105
timestamp 1704896540
transform 1 0 10764 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109_111
timestamp 1704896540
transform 1 0 11316 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_113
timestamp 1704896540
transform 1 0 11500 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_125
timestamp 1704896540
transform 1 0 12604 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_137
timestamp 1704896540
transform 1 0 13708 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_149
timestamp 1704896540
transform 1 0 14812 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_109_161
timestamp 1704896540
transform 1 0 15916 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109_167
timestamp 1704896540
transform 1 0 16468 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_169
timestamp 1704896540
transform 1 0 16652 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_181
timestamp 1704896540
transform 1 0 17756 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_193
timestamp 1704896540
transform 1 0 18860 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_205
timestamp 1704896540
transform 1 0 19964 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_109_217
timestamp 1704896540
transform 1 0 21068 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109_223
timestamp 1704896540
transform 1 0 21620 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_225
timestamp 1704896540
transform 1 0 21804 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_237
timestamp 1704896540
transform 1 0 22908 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_249
timestamp 1704896540
transform 1 0 24012 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_109_261
timestamp 1704896540
transform 1 0 25116 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_109_269
timestamp 1704896540
transform 1 0 25852 0 -1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_109_274
timestamp 1704896540
transform 1 0 26312 0 -1 62016
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_281
timestamp 1704896540
transform 1 0 26956 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_293
timestamp 1704896540
transform 1 0 28060 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_305
timestamp 1704896540
transform 1 0 29164 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_317
timestamp 1704896540
transform 1 0 30268 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_109_329
timestamp 1704896540
transform 1 0 31372 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109_335
timestamp 1704896540
transform 1 0 31924 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_337
timestamp 1704896540
transform 1 0 32108 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_349
timestamp 1704896540
transform 1 0 33212 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_361
timestamp 1704896540
transform 1 0 34316 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_373
timestamp 1704896540
transform 1 0 35420 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_109_385
timestamp 1704896540
transform 1 0 36524 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109_391
timestamp 1704896540
transform 1 0 37076 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_393
timestamp 1704896540
transform 1 0 37260 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_405
timestamp 1704896540
transform 1 0 38364 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_417
timestamp 1704896540
transform 1 0 39468 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_3
timestamp 1704896540
transform 1 0 1380 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_15
timestamp 1704896540
transform 1 0 2484 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_27
timestamp 1704896540
transform 1 0 3588 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_29
timestamp 1704896540
transform 1 0 3772 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_41
timestamp 1704896540
transform 1 0 4876 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_53
timestamp 1704896540
transform 1 0 5980 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_65
timestamp 1704896540
transform 1 0 7084 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_110_77
timestamp 1704896540
transform 1 0 8188 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_83
timestamp 1704896540
transform 1 0 8740 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_85
timestamp 1704896540
transform 1 0 8924 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_97
timestamp 1704896540
transform 1 0 10028 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_109
timestamp 1704896540
transform 1 0 11132 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_121
timestamp 1704896540
transform 1 0 12236 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_110_133
timestamp 1704896540
transform 1 0 13340 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_139
timestamp 1704896540
transform 1 0 13892 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_141
timestamp 1704896540
transform 1 0 14076 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_153
timestamp 1704896540
transform 1 0 15180 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_165
timestamp 1704896540
transform 1 0 16284 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_177
timestamp 1704896540
transform 1 0 17388 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_110_189
timestamp 1704896540
transform 1 0 18492 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_195
timestamp 1704896540
transform 1 0 19044 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_110_197
timestamp 1704896540
transform 1 0 19228 0 1 62016
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_208
timestamp 1704896540
transform 1 0 20240 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_220
timestamp 1704896540
transform 1 0 21344 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_232
timestamp 1704896540
transform 1 0 22448 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_110_244
timestamp 1704896540
transform 1 0 23552 0 1 62016
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_253
timestamp 1704896540
transform 1 0 24380 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_265
timestamp 1704896540
transform 1 0 25484 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_277
timestamp 1704896540
transform 1 0 26588 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_289
timestamp 1704896540
transform 1 0 27692 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_110_301
timestamp 1704896540
transform 1 0 28796 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_307
timestamp 1704896540
transform 1 0 29348 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_309
timestamp 1704896540
transform 1 0 29532 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_321
timestamp 1704896540
transform 1 0 30636 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_333
timestamp 1704896540
transform 1 0 31740 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_345
timestamp 1704896540
transform 1 0 32844 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_110_357
timestamp 1704896540
transform 1 0 33948 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_363
timestamp 1704896540
transform 1 0 34500 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_365
timestamp 1704896540
transform 1 0 34684 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_377
timestamp 1704896540
transform 1 0 35788 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_389
timestamp 1704896540
transform 1 0 36892 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_110_401
timestamp 1704896540
transform 1 0 37996 0 1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_419
timestamp 1704896540
transform 1 0 39652 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_110_421
timestamp 1704896540
transform 1 0 39836 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_425
timestamp 1704896540
transform 1 0 40204 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_3
timestamp 1704896540
transform 1 0 1380 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_15
timestamp 1704896540
transform 1 0 2484 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_27
timestamp 1704896540
transform 1 0 3588 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_39
timestamp 1704896540
transform 1 0 4692 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_111_51
timestamp 1704896540
transform 1 0 5796 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_55
timestamp 1704896540
transform 1 0 6164 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_57
timestamp 1704896540
transform 1 0 6348 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_69
timestamp 1704896540
transform 1 0 7452 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_81
timestamp 1704896540
transform 1 0 8556 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_93
timestamp 1704896540
transform 1 0 9660 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_111_105
timestamp 1704896540
transform 1 0 10764 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_111
timestamp 1704896540
transform 1 0 11316 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_113
timestamp 1704896540
transform 1 0 11500 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_125
timestamp 1704896540
transform 1 0 12604 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_137
timestamp 1704896540
transform 1 0 13708 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_149
timestamp 1704896540
transform 1 0 14812 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_111_161
timestamp 1704896540
transform 1 0 15916 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_167
timestamp 1704896540
transform 1 0 16468 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_169
timestamp 1704896540
transform 1 0 16652 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_181
timestamp 1704896540
transform 1 0 17756 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_193
timestamp 1704896540
transform 1 0 18860 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_208
timestamp 1704896540
transform 1 0 20240 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_111_220
timestamp 1704896540
transform 1 0 21344 0 -1 63104
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_225
timestamp 1704896540
transform 1 0 21804 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_237
timestamp 1704896540
transform 1 0 22908 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_249
timestamp 1704896540
transform 1 0 24012 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_261
timestamp 1704896540
transform 1 0 25116 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_111_273
timestamp 1704896540
transform 1 0 26220 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_279
timestamp 1704896540
transform 1 0 26772 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_281
timestamp 1704896540
transform 1 0 26956 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_293
timestamp 1704896540
transform 1 0 28060 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_305
timestamp 1704896540
transform 1 0 29164 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_317
timestamp 1704896540
transform 1 0 30268 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_111_329
timestamp 1704896540
transform 1 0 31372 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_335
timestamp 1704896540
transform 1 0 31924 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_337
timestamp 1704896540
transform 1 0 32108 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_349
timestamp 1704896540
transform 1 0 33212 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_361
timestamp 1704896540
transform 1 0 34316 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_373
timestamp 1704896540
transform 1 0 35420 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_111_385
timestamp 1704896540
transform 1 0 36524 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_391
timestamp 1704896540
transform 1 0 37076 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_393
timestamp 1704896540
transform 1 0 37260 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_405
timestamp 1704896540
transform 1 0 38364 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_417
timestamp 1704896540
transform 1 0 39468 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_3
timestamp 1704896540
transform 1 0 1380 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_15
timestamp 1704896540
transform 1 0 2484 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_27
timestamp 1704896540
transform 1 0 3588 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_34
timestamp 1704896540
transform 1 0 4232 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_46
timestamp 1704896540
transform 1 0 5336 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_58
timestamp 1704896540
transform 1 0 6440 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_70
timestamp 1704896540
transform 1 0 7544 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_112_82
timestamp 1704896540
transform 1 0 8648 0 1 63104
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_85
timestamp 1704896540
transform 1 0 8924 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_97
timestamp 1704896540
transform 1 0 10028 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_109
timestamp 1704896540
transform 1 0 11132 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_121
timestamp 1704896540
transform 1 0 12236 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_112_133
timestamp 1704896540
transform 1 0 13340 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_139
timestamp 1704896540
transform 1 0 13892 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_141
timestamp 1704896540
transform 1 0 14076 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_153
timestamp 1704896540
transform 1 0 15180 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_165
timestamp 1704896540
transform 1 0 16284 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_177
timestamp 1704896540
transform 1 0 17388 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_112_189
timestamp 1704896540
transform 1 0 18492 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_195
timestamp 1704896540
transform 1 0 19044 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_112_197
timestamp 1704896540
transform 1 0 19228 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_112_205
timestamp 1704896540
transform 1 0 19964 0 1 63104
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_212
timestamp 1704896540
transform 1 0 20608 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_224
timestamp 1704896540
transform 1 0 21712 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_236
timestamp 1704896540
transform 1 0 22816 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_112_248
timestamp 1704896540
transform 1 0 23920 0 1 63104
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_253
timestamp 1704896540
transform 1 0 24380 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_265
timestamp 1704896540
transform 1 0 25484 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_277
timestamp 1704896540
transform 1 0 26588 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_289
timestamp 1704896540
transform 1 0 27692 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_112_301
timestamp 1704896540
transform 1 0 28796 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_307
timestamp 1704896540
transform 1 0 29348 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_309
timestamp 1704896540
transform 1 0 29532 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_321
timestamp 1704896540
transform 1 0 30636 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_333
timestamp 1704896540
transform 1 0 31740 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_345
timestamp 1704896540
transform 1 0 32844 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_112_357
timestamp 1704896540
transform 1 0 33948 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_363
timestamp 1704896540
transform 1 0 34500 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_365
timestamp 1704896540
transform 1 0 34684 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_377
timestamp 1704896540
transform 1 0 35788 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_389
timestamp 1704896540
transform 1 0 36892 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_401
timestamp 1704896540
transform 1 0 37996 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_112_413
timestamp 1704896540
transform 1 0 39100 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_419
timestamp 1704896540
transform 1 0 39652 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_112_421
timestamp 1704896540
transform 1 0 39836 0 1 63104
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_3
timestamp 1704896540
transform 1 0 1380 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_15
timestamp 1704896540
transform 1 0 2484 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_27
timestamp 1704896540
transform 1 0 3588 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_39
timestamp 1704896540
transform 1 0 4692 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113_51
timestamp 1704896540
transform 1 0 5796 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_55
timestamp 1704896540
transform 1 0 6164 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_57
timestamp 1704896540
transform 1 0 6348 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_69
timestamp 1704896540
transform 1 0 7452 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_81
timestamp 1704896540
transform 1 0 8556 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_93
timestamp 1704896540
transform 1 0 9660 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113_105
timestamp 1704896540
transform 1 0 10764 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_111
timestamp 1704896540
transform 1 0 11316 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_113
timestamp 1704896540
transform 1 0 11500 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_125
timestamp 1704896540
transform 1 0 12604 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113_137
timestamp 1704896540
transform 1 0 13708 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113_148
timestamp 1704896540
transform 1 0 14720 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_152
timestamp 1704896540
transform 1 0 15088 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_113_157
timestamp 1704896540
transform 1 0 15548 0 -1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_113_165
timestamp 1704896540
transform 1 0 16284 0 -1 64192
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_169
timestamp 1704896540
transform 1 0 16652 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113_181
timestamp 1704896540
transform 1 0 17756 0 -1 64192
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_193
timestamp 1704896540
transform 1 0 18860 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_113_205
timestamp 1704896540
transform 1 0 19964 0 -1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_213
timestamp 1704896540
transform 1 0 20700 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113_217
timestamp 1704896540
transform 1 0 21068 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_223
timestamp 1704896540
transform 1 0 21620 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_225
timestamp 1704896540
transform 1 0 21804 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_237
timestamp 1704896540
transform 1 0 22908 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_249
timestamp 1704896540
transform 1 0 24012 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_261
timestamp 1704896540
transform 1 0 25116 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113_273
timestamp 1704896540
transform 1 0 26220 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_279
timestamp 1704896540
transform 1 0 26772 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_281
timestamp 1704896540
transform 1 0 26956 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_293
timestamp 1704896540
transform 1 0 28060 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_305
timestamp 1704896540
transform 1 0 29164 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_317
timestamp 1704896540
transform 1 0 30268 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113_329
timestamp 1704896540
transform 1 0 31372 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_335
timestamp 1704896540
transform 1 0 31924 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113_337
timestamp 1704896540
transform 1 0 32108 0 -1 64192
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_344
timestamp 1704896540
transform 1 0 32752 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_356
timestamp 1704896540
transform 1 0 33856 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_368
timestamp 1704896540
transform 1 0 34960 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_380
timestamp 1704896540
transform 1 0 36064 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_393
timestamp 1704896540
transform 1 0 37260 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_405
timestamp 1704896540
transform 1 0 38364 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_417
timestamp 1704896540
transform 1 0 39468 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_3
timestamp 1704896540
transform 1 0 1380 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_15
timestamp 1704896540
transform 1 0 2484 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_27
timestamp 1704896540
transform 1 0 3588 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_29
timestamp 1704896540
transform 1 0 3772 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_41
timestamp 1704896540
transform 1 0 4876 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_53
timestamp 1704896540
transform 1 0 5980 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_65
timestamp 1704896540
transform 1 0 7084 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_114_77
timestamp 1704896540
transform 1 0 8188 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_83
timestamp 1704896540
transform 1 0 8740 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_85
timestamp 1704896540
transform 1 0 8924 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_114_97
timestamp 1704896540
transform 1 0 10028 0 1 64192
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_118
timestamp 1704896540
transform 1 0 11960 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_114_130
timestamp 1704896540
transform 1 0 13064 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_114_138
timestamp 1704896540
transform 1 0 13800 0 1 64192
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_141
timestamp 1704896540
transform 1 0 14076 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_114_153
timestamp 1704896540
transform 1 0 15180 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_114_161
timestamp 1704896540
transform 1 0 15916 0 1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_114_165
timestamp 1704896540
transform 1 0 16284 0 1 64192
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_175
timestamp 1704896540
transform 1 0 17204 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_114_187
timestamp 1704896540
transform 1 0 18308 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_195
timestamp 1704896540
transform 1 0 19044 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_197
timestamp 1704896540
transform 1 0 19228 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_209
timestamp 1704896540
transform 1 0 20332 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_221
timestamp 1704896540
transform 1 0 21436 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_233
timestamp 1704896540
transform 1 0 22540 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_114_245
timestamp 1704896540
transform 1 0 23644 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_251
timestamp 1704896540
transform 1 0 24196 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_253
timestamp 1704896540
transform 1 0 24380 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_114_265
timestamp 1704896540
transform 1 0 25484 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_269
timestamp 1704896540
transform 1 0 25852 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_114_272
timestamp 1704896540
transform 1 0 26128 0 1 64192
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_281
timestamp 1704896540
transform 1 0 26956 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_293
timestamp 1704896540
transform 1 0 28060 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_114_305
timestamp 1704896540
transform 1 0 29164 0 1 64192
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_309
timestamp 1704896540
transform 1 0 29532 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_321
timestamp 1704896540
transform 1 0 30636 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_333
timestamp 1704896540
transform 1 0 31740 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_345
timestamp 1704896540
transform 1 0 32844 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_114_357
timestamp 1704896540
transform 1 0 33948 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_363
timestamp 1704896540
transform 1 0 34500 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_365
timestamp 1704896540
transform 1 0 34684 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_377
timestamp 1704896540
transform 1 0 35788 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_389
timestamp 1704896540
transform 1 0 36892 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_401
timestamp 1704896540
transform 1 0 37996 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_114_413
timestamp 1704896540
transform 1 0 39100 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_419
timestamp 1704896540
transform 1 0 39652 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_114_421
timestamp 1704896540
transform 1 0 39836 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_115_3
timestamp 1704896540
transform 1 0 1380 0 -1 65280
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_15
timestamp 1704896540
transform 1 0 2484 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_27
timestamp 1704896540
transform 1 0 3588 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_39
timestamp 1704896540
transform 1 0 4692 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_115_51
timestamp 1704896540
transform 1 0 5796 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_55
timestamp 1704896540
transform 1 0 6164 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_57
timestamp 1704896540
transform 1 0 6348 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_69
timestamp 1704896540
transform 1 0 7452 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_81
timestamp 1704896540
transform 1 0 8556 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_115_93
timestamp 1704896540
transform 1 0 9660 0 -1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_115_101
timestamp 1704896540
transform 1 0 10396 0 -1 65280
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_115_110
timestamp 1704896540
transform 1 0 11224 0 -1 65280
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_113
timestamp 1704896540
transform 1 0 11500 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_125
timestamp 1704896540
transform 1 0 12604 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_137
timestamp 1704896540
transform 1 0 13708 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_149
timestamp 1704896540
transform 1 0 14812 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_115_161
timestamp 1704896540
transform 1 0 15916 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_167
timestamp 1704896540
transform 1 0 16468 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_169
timestamp 1704896540
transform 1 0 16652 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_181
timestamp 1704896540
transform 1 0 17756 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_193
timestamp 1704896540
transform 1 0 18860 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_205
timestamp 1704896540
transform 1 0 19964 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_115_217
timestamp 1704896540
transform 1 0 21068 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_223
timestamp 1704896540
transform 1 0 21620 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_115_225
timestamp 1704896540
transform 1 0 21804 0 -1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_233
timestamp 1704896540
transform 1 0 22540 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_243
timestamp 1704896540
transform 1 0 23460 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_255
timestamp 1704896540
transform 1 0 24564 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_267
timestamp 1704896540
transform 1 0 25668 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_279
timestamp 1704896540
transform 1 0 26772 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_281
timestamp 1704896540
transform 1 0 26956 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_293
timestamp 1704896540
transform 1 0 28060 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_305
timestamp 1704896540
transform 1 0 29164 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_317
timestamp 1704896540
transform 1 0 30268 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_115_329
timestamp 1704896540
transform 1 0 31372 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_335
timestamp 1704896540
transform 1 0 31924 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_337
timestamp 1704896540
transform 1 0 32108 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_349
timestamp 1704896540
transform 1 0 33212 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_361
timestamp 1704896540
transform 1 0 34316 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_373
timestamp 1704896540
transform 1 0 35420 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_115_385
timestamp 1704896540
transform 1 0 36524 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_391
timestamp 1704896540
transform 1 0 37076 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_393
timestamp 1704896540
transform 1 0 37260 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_405
timestamp 1704896540
transform 1 0 38364 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_417
timestamp 1704896540
transform 1 0 39468 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_3
timestamp 1704896540
transform 1 0 1380 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_15
timestamp 1704896540
transform 1 0 2484 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_27
timestamp 1704896540
transform 1 0 3588 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_29
timestamp 1704896540
transform 1 0 3772 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_41
timestamp 1704896540
transform 1 0 4876 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_116_53
timestamp 1704896540
transform 1 0 5980 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_57
timestamp 1704896540
transform 1 0 6348 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_60
timestamp 1704896540
transform 1 0 6624 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_72
timestamp 1704896540
transform 1 0 7728 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_85
timestamp 1704896540
transform 1 0 8924 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_97
timestamp 1704896540
transform 1 0 10028 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_109
timestamp 1704896540
transform 1 0 11132 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_121
timestamp 1704896540
transform 1 0 12236 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_116_133
timestamp 1704896540
transform 1 0 13340 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_139
timestamp 1704896540
transform 1 0 13892 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_141
timestamp 1704896540
transform 1 0 14076 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_153
timestamp 1704896540
transform 1 0 15180 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_165
timestamp 1704896540
transform 1 0 16284 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_177
timestamp 1704896540
transform 1 0 17388 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_116_189
timestamp 1704896540
transform 1 0 18492 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_195
timestamp 1704896540
transform 1 0 19044 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_197
timestamp 1704896540
transform 1 0 19228 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_209
timestamp 1704896540
transform 1 0 20332 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_221
timestamp 1704896540
transform 1 0 21436 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_233
timestamp 1704896540
transform 1 0 22540 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_116_245
timestamp 1704896540
transform 1 0 23644 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_251
timestamp 1704896540
transform 1 0 24196 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_253
timestamp 1704896540
transform 1 0 24380 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_265
timestamp 1704896540
transform 1 0 25484 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_277
timestamp 1704896540
transform 1 0 26588 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_289
timestamp 1704896540
transform 1 0 27692 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_116_301
timestamp 1704896540
transform 1 0 28796 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_307
timestamp 1704896540
transform 1 0 29348 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_309
timestamp 1704896540
transform 1 0 29532 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_321
timestamp 1704896540
transform 1 0 30636 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_333
timestamp 1704896540
transform 1 0 31740 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_345
timestamp 1704896540
transform 1 0 32844 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_116_357
timestamp 1704896540
transform 1 0 33948 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_363
timestamp 1704896540
transform 1 0 34500 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_365
timestamp 1704896540
transform 1 0 34684 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_377
timestamp 1704896540
transform 1 0 35788 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_389
timestamp 1704896540
transform 1 0 36892 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_401
timestamp 1704896540
transform 1 0 37996 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_116_413
timestamp 1704896540
transform 1 0 39100 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_419
timestamp 1704896540
transform 1 0 39652 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_116_421
timestamp 1704896540
transform 1 0 39836 0 1 65280
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_3
timestamp 1704896540
transform 1 0 1380 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_15
timestamp 1704896540
transform 1 0 2484 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_27
timestamp 1704896540
transform 1 0 3588 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_39
timestamp 1704896540
transform 1 0 4692 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_117_51
timestamp 1704896540
transform 1 0 5796 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_55
timestamp 1704896540
transform 1 0 6164 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_57
timestamp 1704896540
transform 1 0 6348 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_69
timestamp 1704896540
transform 1 0 7452 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_81
timestamp 1704896540
transform 1 0 8556 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_93
timestamp 1704896540
transform 1 0 9660 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_117_105
timestamp 1704896540
transform 1 0 10764 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_111
timestamp 1704896540
transform 1 0 11316 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_113
timestamp 1704896540
transform 1 0 11500 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_125
timestamp 1704896540
transform 1 0 12604 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_137
timestamp 1704896540
transform 1 0 13708 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_149
timestamp 1704896540
transform 1 0 14812 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_117_161
timestamp 1704896540
transform 1 0 15916 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_167
timestamp 1704896540
transform 1 0 16468 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_169
timestamp 1704896540
transform 1 0 16652 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_181
timestamp 1704896540
transform 1 0 17756 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_193
timestamp 1704896540
transform 1 0 18860 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_205
timestamp 1704896540
transform 1 0 19964 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_117_217
timestamp 1704896540
transform 1 0 21068 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_223
timestamp 1704896540
transform 1 0 21620 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_225
timestamp 1704896540
transform 1 0 21804 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_237
timestamp 1704896540
transform 1 0 22908 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_117_240
timestamp 1704896540
transform 1 0 23184 0 -1 66368
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_247
timestamp 1704896540
transform 1 0 23828 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_259
timestamp 1704896540
transform 1 0 24932 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_117_271
timestamp 1704896540
transform 1 0 26036 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_279
timestamp 1704896540
transform 1 0 26772 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_281
timestamp 1704896540
transform 1 0 26956 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_293
timestamp 1704896540
transform 1 0 28060 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_305
timestamp 1704896540
transform 1 0 29164 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_317
timestamp 1704896540
transform 1 0 30268 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_117_329
timestamp 1704896540
transform 1 0 31372 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_335
timestamp 1704896540
transform 1 0 31924 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_337
timestamp 1704896540
transform 1 0 32108 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_349
timestamp 1704896540
transform 1 0 33212 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_361
timestamp 1704896540
transform 1 0 34316 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_373
timestamp 1704896540
transform 1 0 35420 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_117_385
timestamp 1704896540
transform 1 0 36524 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_391
timestamp 1704896540
transform 1 0 37076 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_393
timestamp 1704896540
transform 1 0 37260 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_405
timestamp 1704896540
transform 1 0 38364 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_417
timestamp 1704896540
transform 1 0 39468 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_3
timestamp 1704896540
transform 1 0 1380 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_15
timestamp 1704896540
transform 1 0 2484 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_27
timestamp 1704896540
transform 1 0 3588 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_29
timestamp 1704896540
transform 1 0 3772 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_41
timestamp 1704896540
transform 1 0 4876 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_118_53
timestamp 1704896540
transform 1 0 5980 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_57
timestamp 1704896540
transform 1 0 6348 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_62
timestamp 1704896540
transform 1 0 6808 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_118_74
timestamp 1704896540
transform 1 0 7912 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_118_82
timestamp 1704896540
transform 1 0 8648 0 1 66368
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_85
timestamp 1704896540
transform 1 0 8924 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_97
timestamp 1704896540
transform 1 0 10028 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_109
timestamp 1704896540
transform 1 0 11132 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_121
timestamp 1704896540
transform 1 0 12236 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118_133
timestamp 1704896540
transform 1 0 13340 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_139
timestamp 1704896540
transform 1 0 13892 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_141
timestamp 1704896540
transform 1 0 14076 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_153
timestamp 1704896540
transform 1 0 15180 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_165
timestamp 1704896540
transform 1 0 16284 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_177
timestamp 1704896540
transform 1 0 17388 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118_189
timestamp 1704896540
transform 1 0 18492 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_195
timestamp 1704896540
transform 1 0 19044 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_197
timestamp 1704896540
transform 1 0 19228 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_209
timestamp 1704896540
transform 1 0 20332 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_221
timestamp 1704896540
transform 1 0 21436 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_233
timestamp 1704896540
transform 1 0 22540 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118_245
timestamp 1704896540
transform 1 0 23644 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_251
timestamp 1704896540
transform 1 0 24196 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_253
timestamp 1704896540
transform 1 0 24380 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_265
timestamp 1704896540
transform 1 0 25484 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_277
timestamp 1704896540
transform 1 0 26588 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_289
timestamp 1704896540
transform 1 0 27692 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118_301
timestamp 1704896540
transform 1 0 28796 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_307
timestamp 1704896540
transform 1 0 29348 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_309
timestamp 1704896540
transform 1 0 29532 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_321
timestamp 1704896540
transform 1 0 30636 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_333
timestamp 1704896540
transform 1 0 31740 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_345
timestamp 1704896540
transform 1 0 32844 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118_357
timestamp 1704896540
transform 1 0 33948 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_363
timestamp 1704896540
transform 1 0 34500 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_365
timestamp 1704896540
transform 1 0 34684 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_377
timestamp 1704896540
transform 1 0 35788 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_389
timestamp 1704896540
transform 1 0 36892 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_401
timestamp 1704896540
transform 1 0 37996 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118_413
timestamp 1704896540
transform 1 0 39100 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_419
timestamp 1704896540
transform 1 0 39652 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_118_421
timestamp 1704896540
transform 1 0 39836 0 1 66368
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_3
timestamp 1704896540
transform 1 0 1380 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_15
timestamp 1704896540
transform 1 0 2484 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_27
timestamp 1704896540
transform 1 0 3588 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_39
timestamp 1704896540
transform 1 0 4692 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_119_51
timestamp 1704896540
transform 1 0 5796 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119_55
timestamp 1704896540
transform 1 0 6164 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_57
timestamp 1704896540
transform 1 0 6348 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_69
timestamp 1704896540
transform 1 0 7452 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_81
timestamp 1704896540
transform 1 0 8556 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_93
timestamp 1704896540
transform 1 0 9660 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_119_105
timestamp 1704896540
transform 1 0 10764 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119_111
timestamp 1704896540
transform 1 0 11316 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_113
timestamp 1704896540
transform 1 0 11500 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_125
timestamp 1704896540
transform 1 0 12604 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_119_137
timestamp 1704896540
transform 1 0 13708 0 -1 67456
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_154
timestamp 1704896540
transform 1 0 15272 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_119_166
timestamp 1704896540
transform 1 0 16376 0 -1 67456
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_169
timestamp 1704896540
transform 1 0 16652 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_181
timestamp 1704896540
transform 1 0 17756 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_193
timestamp 1704896540
transform 1 0 18860 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_205
timestamp 1704896540
transform 1 0 19964 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_119_217
timestamp 1704896540
transform 1 0 21068 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119_223
timestamp 1704896540
transform 1 0 21620 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_225
timestamp 1704896540
transform 1 0 21804 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_237
timestamp 1704896540
transform 1 0 22908 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_249
timestamp 1704896540
transform 1 0 24012 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_261
timestamp 1704896540
transform 1 0 25116 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_119_273
timestamp 1704896540
transform 1 0 26220 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119_279
timestamp 1704896540
transform 1 0 26772 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_281
timestamp 1704896540
transform 1 0 26956 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_293
timestamp 1704896540
transform 1 0 28060 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_305
timestamp 1704896540
transform 1 0 29164 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_317
timestamp 1704896540
transform 1 0 30268 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_119_329
timestamp 1704896540
transform 1 0 31372 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119_335
timestamp 1704896540
transform 1 0 31924 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_337
timestamp 1704896540
transform 1 0 32108 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_349
timestamp 1704896540
transform 1 0 33212 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_361
timestamp 1704896540
transform 1 0 34316 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_373
timestamp 1704896540
transform 1 0 35420 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_119_385
timestamp 1704896540
transform 1 0 36524 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119_391
timestamp 1704896540
transform 1 0 37076 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_393
timestamp 1704896540
transform 1 0 37260 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_405
timestamp 1704896540
transform 1 0 38364 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_417
timestamp 1704896540
transform 1 0 39468 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_120_3
timestamp 1704896540
transform 1 0 1380 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_120_9
timestamp 1704896540
transform 1 0 1932 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_13
timestamp 1704896540
transform 1 0 2300 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_120_25
timestamp 1704896540
transform 1 0 3404 0 1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_29
timestamp 1704896540
transform 1 0 3772 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_41
timestamp 1704896540
transform 1 0 4876 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_120_53
timestamp 1704896540
transform 1 0 5980 0 1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_59
timestamp 1704896540
transform 1 0 6532 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_71
timestamp 1704896540
transform 1 0 7636 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_120_83
timestamp 1704896540
transform 1 0 8740 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_85
timestamp 1704896540
transform 1 0 8924 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_97
timestamp 1704896540
transform 1 0 10028 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_109
timestamp 1704896540
transform 1 0 11132 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_121
timestamp 1704896540
transform 1 0 12236 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_120_133
timestamp 1704896540
transform 1 0 13340 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_120_139
timestamp 1704896540
transform 1 0 13892 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_141
timestamp 1704896540
transform 1 0 14076 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_153
timestamp 1704896540
transform 1 0 15180 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_165
timestamp 1704896540
transform 1 0 16284 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_177
timestamp 1704896540
transform 1 0 17388 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_120_189
timestamp 1704896540
transform 1 0 18492 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_120_195
timestamp 1704896540
transform 1 0 19044 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_197
timestamp 1704896540
transform 1 0 19228 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_209
timestamp 1704896540
transform 1 0 20332 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_221
timestamp 1704896540
transform 1 0 21436 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_233
timestamp 1704896540
transform 1 0 22540 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_120_245
timestamp 1704896540
transform 1 0 23644 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_120_251
timestamp 1704896540
transform 1 0 24196 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_120_253
timestamp 1704896540
transform 1 0 24380 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_120_257
timestamp 1704896540
transform 1 0 24748 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_263
timestamp 1704896540
transform 1 0 25300 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_275
timestamp 1704896540
transform 1 0 26404 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_287
timestamp 1704896540
transform 1 0 27508 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_120_299
timestamp 1704896540
transform 1 0 28612 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_120_307
timestamp 1704896540
transform 1 0 29348 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_309
timestamp 1704896540
transform 1 0 29532 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_321
timestamp 1704896540
transform 1 0 30636 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_333
timestamp 1704896540
transform 1 0 31740 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_345
timestamp 1704896540
transform 1 0 32844 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_120_357
timestamp 1704896540
transform 1 0 33948 0 1 67456
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_365
timestamp 1704896540
transform 1 0 34684 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_377
timestamp 1704896540
transform 1 0 35788 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_389
timestamp 1704896540
transform 1 0 36892 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_401
timestamp 1704896540
transform 1 0 37996 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_120_413
timestamp 1704896540
transform 1 0 39100 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_120_419
timestamp 1704896540
transform 1 0 39652 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_120_421
timestamp 1704896540
transform 1 0 39836 0 1 67456
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_3
timestamp 1704896540
transform 1 0 1380 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_15
timestamp 1704896540
transform 1 0 2484 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_27
timestamp 1704896540
transform 1 0 3588 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_39
timestamp 1704896540
transform 1 0 4692 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_121_51
timestamp 1704896540
transform 1 0 5796 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_121_55
timestamp 1704896540
transform 1 0 6164 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_121_57
timestamp 1704896540
transform 1 0 6348 0 -1 68544
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_70
timestamp 1704896540
transform 1 0 7544 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_121_82
timestamp 1704896540
transform 1 0 8648 0 -1 68544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_91
timestamp 1704896540
transform 1 0 9476 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_121_103
timestamp 1704896540
transform 1 0 10580 0 -1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_121_111
timestamp 1704896540
transform 1 0 11316 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_113
timestamp 1704896540
transform 1 0 11500 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_125
timestamp 1704896540
transform 1 0 12604 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_137
timestamp 1704896540
transform 1 0 13708 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_149
timestamp 1704896540
transform 1 0 14812 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_121_161
timestamp 1704896540
transform 1 0 15916 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_121_167
timestamp 1704896540
transform 1 0 16468 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_169
timestamp 1704896540
transform 1 0 16652 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_181
timestamp 1704896540
transform 1 0 17756 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_193
timestamp 1704896540
transform 1 0 18860 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_205
timestamp 1704896540
transform 1 0 19964 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_121_217
timestamp 1704896540
transform 1 0 21068 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_121_223
timestamp 1704896540
transform 1 0 21620 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_225
timestamp 1704896540
transform 1 0 21804 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_237
timestamp 1704896540
transform 1 0 22908 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_249
timestamp 1704896540
transform 1 0 24012 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_261
timestamp 1704896540
transform 1 0 25116 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_121_273
timestamp 1704896540
transform 1 0 26220 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_121_279
timestamp 1704896540
transform 1 0 26772 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_281
timestamp 1704896540
transform 1 0 26956 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_293
timestamp 1704896540
transform 1 0 28060 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_305
timestamp 1704896540
transform 1 0 29164 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_317
timestamp 1704896540
transform 1 0 30268 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_121_329
timestamp 1704896540
transform 1 0 31372 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_121_335
timestamp 1704896540
transform 1 0 31924 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_345
timestamp 1704896540
transform 1 0 32844 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_357
timestamp 1704896540
transform 1 0 33948 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_369
timestamp 1704896540
transform 1 0 35052 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_121_381
timestamp 1704896540
transform 1 0 36156 0 -1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_121_389
timestamp 1704896540
transform 1 0 36892 0 -1 68544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_393
timestamp 1704896540
transform 1 0 37260 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_405
timestamp 1704896540
transform 1 0 38364 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_417
timestamp 1704896540
transform 1 0 39468 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_3
timestamp 1704896540
transform 1 0 1380 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_15
timestamp 1704896540
transform 1 0 2484 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_122_27
timestamp 1704896540
transform 1 0 3588 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_29
timestamp 1704896540
transform 1 0 3772 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_41
timestamp 1704896540
transform 1 0 4876 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_53
timestamp 1704896540
transform 1 0 5980 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_65
timestamp 1704896540
transform 1 0 7084 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_122_77
timestamp 1704896540
transform 1 0 8188 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_122_83
timestamp 1704896540
transform 1 0 8740 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_85
timestamp 1704896540
transform 1 0 8924 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_97
timestamp 1704896540
transform 1 0 10028 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_109
timestamp 1704896540
transform 1 0 11132 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_121
timestamp 1704896540
transform 1 0 12236 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_122_133
timestamp 1704896540
transform 1 0 13340 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_122_139
timestamp 1704896540
transform 1 0 13892 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_141
timestamp 1704896540
transform 1 0 14076 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_153
timestamp 1704896540
transform 1 0 15180 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_165
timestamp 1704896540
transform 1 0 16284 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_177
timestamp 1704896540
transform 1 0 17388 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_122_189
timestamp 1704896540
transform 1 0 18492 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_122_195
timestamp 1704896540
transform 1 0 19044 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_197
timestamp 1704896540
transform 1 0 19228 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_209
timestamp 1704896540
transform 1 0 20332 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_221
timestamp 1704896540
transform 1 0 21436 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_233
timestamp 1704896540
transform 1 0 22540 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_122_245
timestamp 1704896540
transform 1 0 23644 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_122_251
timestamp 1704896540
transform 1 0 24196 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_253
timestamp 1704896540
transform 1 0 24380 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_265
timestamp 1704896540
transform 1 0 25484 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_277
timestamp 1704896540
transform 1 0 26588 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_289
timestamp 1704896540
transform 1 0 27692 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_122_301
timestamp 1704896540
transform 1 0 28796 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_122_307
timestamp 1704896540
transform 1 0 29348 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_309
timestamp 1704896540
transform 1 0 29532 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_321
timestamp 1704896540
transform 1 0 30636 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_333
timestamp 1704896540
transform 1 0 31740 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_345
timestamp 1704896540
transform 1 0 32844 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_122_357
timestamp 1704896540
transform 1 0 33948 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_122_363
timestamp 1704896540
transform 1 0 34500 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_122_365
timestamp 1704896540
transform 1 0 34684 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_122_373
timestamp 1704896540
transform 1 0 35420 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_122_377
timestamp 1704896540
transform 1 0 35788 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_122_388
timestamp 1704896540
transform 1 0 36800 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_122_392
timestamp 1704896540
transform 1 0 37168 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_122_398
timestamp 1704896540
transform 1 0 37720 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_402
timestamp 1704896540
transform 1 0 38088 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_122_414
timestamp 1704896540
transform 1 0 39192 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_122_421
timestamp 1704896540
transform 1 0 39836 0 1 68544
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_3
timestamp 1704896540
transform 1 0 1380 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_123_15
timestamp 1704896540
transform 1 0 2484 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_123_24
timestamp 1704896540
transform 1 0 3312 0 -1 69632
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_29
timestamp 1704896540
transform 1 0 3772 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_41
timestamp 1704896540
transform 1 0 4876 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_123_53
timestamp 1704896540
transform 1 0 5980 0 -1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_57
timestamp 1704896540
transform 1 0 6348 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_69
timestamp 1704896540
transform 1 0 7452 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_123_81
timestamp 1704896540
transform 1 0 8556 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_123_85
timestamp 1704896540
transform 1 0 8924 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_89
timestamp 1704896540
transform 1 0 9292 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_123_101
timestamp 1704896540
transform 1 0 10396 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_123_109
timestamp 1704896540
transform 1 0 11132 0 -1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_113
timestamp 1704896540
transform 1 0 11500 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_125
timestamp 1704896540
transform 1 0 12604 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_123_137
timestamp 1704896540
transform 1 0 13708 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_123_141
timestamp 1704896540
transform 1 0 14076 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_123_149
timestamp 1704896540
transform 1 0 14812 0 -1 69632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_154
timestamp 1704896540
transform 1 0 15272 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_123_166
timestamp 1704896540
transform 1 0 16376 0 -1 69632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_169
timestamp 1704896540
transform 1 0 16652 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_181
timestamp 1704896540
transform 1 0 17756 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_123_193
timestamp 1704896540
transform 1 0 18860 0 -1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_197
timestamp 1704896540
transform 1 0 19228 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_123_209
timestamp 1704896540
transform 1 0 20332 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_123_215
timestamp 1704896540
transform 1 0 20884 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_123_219
timestamp 1704896540
transform 1 0 21252 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_123_223
timestamp 1704896540
transform 1 0 21620 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_225
timestamp 1704896540
transform 1 0 21804 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_237
timestamp 1704896540
transform 1 0 22908 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_123_249
timestamp 1704896540
transform 1 0 24012 0 -1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_253
timestamp 1704896540
transform 1 0 24380 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_265
timestamp 1704896540
transform 1 0 25484 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_123_277
timestamp 1704896540
transform 1 0 26588 0 -1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_284
timestamp 1704896540
transform 1 0 27232 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_296
timestamp 1704896540
transform 1 0 28336 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_309
timestamp 1704896540
transform 1 0 29532 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_321
timestamp 1704896540
transform 1 0 30636 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_123_333
timestamp 1704896540
transform 1 0 31740 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_123_337
timestamp 1704896540
transform 1 0 32108 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_123_345
timestamp 1704896540
transform 1 0 32844 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_349
timestamp 1704896540
transform 1 0 33212 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_123_361
timestamp 1704896540
transform 1 0 34316 0 -1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_365
timestamp 1704896540
transform 1 0 34684 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_377
timestamp 1704896540
transform 1 0 35788 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_123_389
timestamp 1704896540
transform 1 0 36892 0 -1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_393
timestamp 1704896540
transform 1 0 37260 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_123_405
timestamp 1704896540
transform 1 0 38364 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_123_414
timestamp 1704896540
transform 1 0 39192 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_123_421
timestamp 1704896540
transform 1 0 39836 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 40572 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  output2
timestamp 1704896540
transform -1 0 39192 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output3
timestamp 1704896540
transform -1 0 33212 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output4
timestamp 1704896540
transform -1 0 27232 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output5
timestamp 1704896540
transform -1 0 21252 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output6
timestamp 1704896540
transform -1 0 15272 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output7
timestamp 1704896540
transform -1 0 9292 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output8
timestamp 1704896540
transform -1 0 3312 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_124
timestamp 1704896540
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1704896540
transform -1 0 40848 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_125
timestamp 1704896540
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1704896540
transform -1 0 40848 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_126
timestamp 1704896540
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1704896540
transform -1 0 40848 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_127
timestamp 1704896540
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1704896540
transform -1 0 40848 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_128
timestamp 1704896540
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1704896540
transform -1 0 40848 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_129
timestamp 1704896540
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1704896540
transform -1 0 40848 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_130
timestamp 1704896540
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1704896540
transform -1 0 40848 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_131
timestamp 1704896540
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1704896540
transform -1 0 40848 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_132
timestamp 1704896540
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1704896540
transform -1 0 40848 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_133
timestamp 1704896540
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1704896540
transform -1 0 40848 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_134
timestamp 1704896540
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1704896540
transform -1 0 40848 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_135
timestamp 1704896540
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1704896540
transform -1 0 40848 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_136
timestamp 1704896540
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1704896540
transform -1 0 40848 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_137
timestamp 1704896540
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1704896540
transform -1 0 40848 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_138
timestamp 1704896540
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1704896540
transform -1 0 40848 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_139
timestamp 1704896540
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1704896540
transform -1 0 40848 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_140
timestamp 1704896540
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1704896540
transform -1 0 40848 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_141
timestamp 1704896540
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1704896540
transform -1 0 40848 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_142
timestamp 1704896540
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1704896540
transform -1 0 40848 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_143
timestamp 1704896540
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1704896540
transform -1 0 40848 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_144
timestamp 1704896540
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1704896540
transform -1 0 40848 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_145
timestamp 1704896540
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1704896540
transform -1 0 40848 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_146
timestamp 1704896540
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1704896540
transform -1 0 40848 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_147
timestamp 1704896540
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1704896540
transform -1 0 40848 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_148
timestamp 1704896540
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1704896540
transform -1 0 40848 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_149
timestamp 1704896540
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1704896540
transform -1 0 40848 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_150
timestamp 1704896540
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1704896540
transform -1 0 40848 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_151
timestamp 1704896540
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1704896540
transform -1 0 40848 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_152
timestamp 1704896540
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1704896540
transform -1 0 40848 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_153
timestamp 1704896540
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1704896540
transform -1 0 40848 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_154
timestamp 1704896540
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1704896540
transform -1 0 40848 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_155
timestamp 1704896540
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1704896540
transform -1 0 40848 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_156
timestamp 1704896540
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1704896540
transform -1 0 40848 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_157
timestamp 1704896540
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1704896540
transform -1 0 40848 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_158
timestamp 1704896540
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1704896540
transform -1 0 40848 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_159
timestamp 1704896540
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1704896540
transform -1 0 40848 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_160
timestamp 1704896540
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 1704896540
transform -1 0 40848 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_161
timestamp 1704896540
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 1704896540
transform -1 0 40848 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_162
timestamp 1704896540
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 1704896540
transform -1 0 40848 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_163
timestamp 1704896540
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 1704896540
transform -1 0 40848 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_164
timestamp 1704896540
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 1704896540
transform -1 0 40848 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_165
timestamp 1704896540
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 1704896540
transform -1 0 40848 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_166
timestamp 1704896540
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp 1704896540
transform -1 0 40848 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_167
timestamp 1704896540
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp 1704896540
transform -1 0 40848 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_168
timestamp 1704896540
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp 1704896540
transform -1 0 40848 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_169
timestamp 1704896540
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp 1704896540
transform -1 0 40848 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_170
timestamp 1704896540
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp 1704896540
transform -1 0 40848 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_171
timestamp 1704896540
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp 1704896540
transform -1 0 40848 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Left_172
timestamp 1704896540
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Right_48
timestamp 1704896540
transform -1 0 40848 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Left_173
timestamp 1704896540
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Right_49
timestamp 1704896540
transform -1 0 40848 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Left_174
timestamp 1704896540
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Right_50
timestamp 1704896540
transform -1 0 40848 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Left_175
timestamp 1704896540
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Right_51
timestamp 1704896540
transform -1 0 40848 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Left_176
timestamp 1704896540
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Right_52
timestamp 1704896540
transform -1 0 40848 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Left_177
timestamp 1704896540
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Right_53
timestamp 1704896540
transform -1 0 40848 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Left_178
timestamp 1704896540
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Right_54
timestamp 1704896540
transform -1 0 40848 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Left_179
timestamp 1704896540
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Right_55
timestamp 1704896540
transform -1 0 40848 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Left_180
timestamp 1704896540
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Right_56
timestamp 1704896540
transform -1 0 40848 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Left_181
timestamp 1704896540
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Right_57
timestamp 1704896540
transform -1 0 40848 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Left_182
timestamp 1704896540
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Right_58
timestamp 1704896540
transform -1 0 40848 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Left_183
timestamp 1704896540
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Right_59
timestamp 1704896540
transform -1 0 40848 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Left_184
timestamp 1704896540
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Right_60
timestamp 1704896540
transform -1 0 40848 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Left_185
timestamp 1704896540
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Right_61
timestamp 1704896540
transform -1 0 40848 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Left_186
timestamp 1704896540
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Right_62
timestamp 1704896540
transform -1 0 40848 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Left_187
timestamp 1704896540
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Right_63
timestamp 1704896540
transform -1 0 40848 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Left_188
timestamp 1704896540
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Right_64
timestamp 1704896540
transform -1 0 40848 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_Left_189
timestamp 1704896540
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_Right_65
timestamp 1704896540
transform -1 0 40848 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_Left_190
timestamp 1704896540
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_Right_66
timestamp 1704896540
transform -1 0 40848 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_Left_191
timestamp 1704896540
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_Right_67
timestamp 1704896540
transform -1 0 40848 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_Left_192
timestamp 1704896540
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_Right_68
timestamp 1704896540
transform -1 0 40848 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_Left_193
timestamp 1704896540
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_Right_69
timestamp 1704896540
transform -1 0 40848 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_Left_194
timestamp 1704896540
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_Right_70
timestamp 1704896540
transform -1 0 40848 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_Left_195
timestamp 1704896540
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_Right_71
timestamp 1704896540
transform -1 0 40848 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_Left_196
timestamp 1704896540
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_Right_72
timestamp 1704896540
transform -1 0 40848 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_Left_197
timestamp 1704896540
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_Right_73
timestamp 1704896540
transform -1 0 40848 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_Left_198
timestamp 1704896540
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_Right_74
timestamp 1704896540
transform -1 0 40848 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_Left_199
timestamp 1704896540
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_Right_75
timestamp 1704896540
transform -1 0 40848 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_Left_200
timestamp 1704896540
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_Right_76
timestamp 1704896540
transform -1 0 40848 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_Left_201
timestamp 1704896540
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_Right_77
timestamp 1704896540
transform -1 0 40848 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_Left_202
timestamp 1704896540
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_Right_78
timestamp 1704896540
transform -1 0 40848 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_Left_203
timestamp 1704896540
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_Right_79
timestamp 1704896540
transform -1 0 40848 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_Left_204
timestamp 1704896540
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_Right_80
timestamp 1704896540
transform -1 0 40848 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_Left_205
timestamp 1704896540
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_Right_81
timestamp 1704896540
transform -1 0 40848 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_Left_206
timestamp 1704896540
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_Right_82
timestamp 1704896540
transform -1 0 40848 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_Left_207
timestamp 1704896540
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_Right_83
timestamp 1704896540
transform -1 0 40848 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_Left_208
timestamp 1704896540
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_Right_84
timestamp 1704896540
transform -1 0 40848 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_Left_209
timestamp 1704896540
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_Right_85
timestamp 1704896540
transform -1 0 40848 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_Left_210
timestamp 1704896540
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_Right_86
timestamp 1704896540
transform -1 0 40848 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_Left_211
timestamp 1704896540
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_Right_87
timestamp 1704896540
transform -1 0 40848 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_Left_212
timestamp 1704896540
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_Right_88
timestamp 1704896540
transform -1 0 40848 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_Left_213
timestamp 1704896540
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_Right_89
timestamp 1704896540
transform -1 0 40848 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_Left_214
timestamp 1704896540
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_Right_90
timestamp 1704896540
transform -1 0 40848 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_Left_215
timestamp 1704896540
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_Right_91
timestamp 1704896540
transform -1 0 40848 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_Left_216
timestamp 1704896540
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_Right_92
timestamp 1704896540
transform -1 0 40848 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_Left_217
timestamp 1704896540
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_Right_93
timestamp 1704896540
transform -1 0 40848 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_Left_218
timestamp 1704896540
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_Right_94
timestamp 1704896540
transform -1 0 40848 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_Left_219
timestamp 1704896540
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_Right_95
timestamp 1704896540
transform -1 0 40848 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_Left_220
timestamp 1704896540
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_Right_96
timestamp 1704896540
transform -1 0 40848 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_Left_221
timestamp 1704896540
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_Right_97
timestamp 1704896540
transform -1 0 40848 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_Left_222
timestamp 1704896540
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_Right_98
timestamp 1704896540
transform -1 0 40848 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_Left_223
timestamp 1704896540
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_Right_99
timestamp 1704896540
transform -1 0 40848 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_Left_224
timestamp 1704896540
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_Right_100
timestamp 1704896540
transform -1 0 40848 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_Left_225
timestamp 1704896540
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_Right_101
timestamp 1704896540
transform -1 0 40848 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_Left_226
timestamp 1704896540
transform 1 0 1104 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_Right_102
timestamp 1704896540
transform -1 0 40848 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_Left_227
timestamp 1704896540
transform 1 0 1104 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_Right_103
timestamp 1704896540
transform -1 0 40848 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_Left_228
timestamp 1704896540
transform 1 0 1104 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_Right_104
timestamp 1704896540
transform -1 0 40848 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_Left_229
timestamp 1704896540
transform 1 0 1104 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_Right_105
timestamp 1704896540
transform -1 0 40848 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_Left_230
timestamp 1704896540
transform 1 0 1104 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_Right_106
timestamp 1704896540
transform -1 0 40848 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_Left_231
timestamp 1704896540
transform 1 0 1104 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_Right_107
timestamp 1704896540
transform -1 0 40848 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_Left_232
timestamp 1704896540
transform 1 0 1104 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_Right_108
timestamp 1704896540
transform -1 0 40848 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_Left_233
timestamp 1704896540
transform 1 0 1104 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_Right_109
timestamp 1704896540
transform -1 0 40848 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_Left_234
timestamp 1704896540
transform 1 0 1104 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_Right_110
timestamp 1704896540
transform -1 0 40848 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_Left_235
timestamp 1704896540
transform 1 0 1104 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_Right_111
timestamp 1704896540
transform -1 0 40848 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_Left_236
timestamp 1704896540
transform 1 0 1104 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_Right_112
timestamp 1704896540
transform -1 0 40848 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_Left_237
timestamp 1704896540
transform 1 0 1104 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_Right_113
timestamp 1704896540
transform -1 0 40848 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_Left_238
timestamp 1704896540
transform 1 0 1104 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_Right_114
timestamp 1704896540
transform -1 0 40848 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_Left_239
timestamp 1704896540
transform 1 0 1104 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_Right_115
timestamp 1704896540
transform -1 0 40848 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_Left_240
timestamp 1704896540
transform 1 0 1104 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_Right_116
timestamp 1704896540
transform -1 0 40848 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_Left_241
timestamp 1704896540
transform 1 0 1104 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_Right_117
timestamp 1704896540
transform -1 0 40848 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_Left_242
timestamp 1704896540
transform 1 0 1104 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_Right_118
timestamp 1704896540
transform -1 0 40848 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_Left_243
timestamp 1704896540
transform 1 0 1104 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_Right_119
timestamp 1704896540
transform -1 0 40848 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_Left_244
timestamp 1704896540
transform 1 0 1104 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_Right_120
timestamp 1704896540
transform -1 0 40848 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_Left_245
timestamp 1704896540
transform 1 0 1104 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_Right_121
timestamp 1704896540
transform -1 0 40848 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_Left_246
timestamp 1704896540
transform 1 0 1104 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_Right_122
timestamp 1704896540
transform -1 0 40848 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_Left_247
timestamp 1704896540
transform 1 0 1104 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_Right_123
timestamp 1704896540
transform -1 0 40848 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_248 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_249
timestamp 1704896540
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_250
timestamp 1704896540
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_251
timestamp 1704896540
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_252
timestamp 1704896540
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_253
timestamp 1704896540
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_254
timestamp 1704896540
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_255
timestamp 1704896540
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_256
timestamp 1704896540
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_257
timestamp 1704896540
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_258
timestamp 1704896540
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_259
timestamp 1704896540
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_260
timestamp 1704896540
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_261
timestamp 1704896540
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_262
timestamp 1704896540
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_263
timestamp 1704896540
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_264
timestamp 1704896540
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_265
timestamp 1704896540
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_266
timestamp 1704896540
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_267
timestamp 1704896540
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_268
timestamp 1704896540
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_269
timestamp 1704896540
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_270
timestamp 1704896540
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_271
timestamp 1704896540
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_272
timestamp 1704896540
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_273
timestamp 1704896540
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_274
timestamp 1704896540
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_275
timestamp 1704896540
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_276
timestamp 1704896540
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_277
timestamp 1704896540
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_278
timestamp 1704896540
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_279
timestamp 1704896540
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_280
timestamp 1704896540
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_281
timestamp 1704896540
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_282
timestamp 1704896540
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_283
timestamp 1704896540
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_284
timestamp 1704896540
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_285
timestamp 1704896540
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_286
timestamp 1704896540
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_287
timestamp 1704896540
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_288
timestamp 1704896540
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_289
timestamp 1704896540
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_290
timestamp 1704896540
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_291
timestamp 1704896540
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_292
timestamp 1704896540
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_293
timestamp 1704896540
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_294
timestamp 1704896540
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_295
timestamp 1704896540
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_296
timestamp 1704896540
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_297
timestamp 1704896540
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_298
timestamp 1704896540
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_299
timestamp 1704896540
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_300
timestamp 1704896540
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_301
timestamp 1704896540
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_302
timestamp 1704896540
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_303
timestamp 1704896540
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_304
timestamp 1704896540
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_305
timestamp 1704896540
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_306
timestamp 1704896540
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_307
timestamp 1704896540
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_308
timestamp 1704896540
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_309
timestamp 1704896540
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_310
timestamp 1704896540
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_311
timestamp 1704896540
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_312
timestamp 1704896540
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_313
timestamp 1704896540
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_314
timestamp 1704896540
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_315
timestamp 1704896540
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_316
timestamp 1704896540
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_317
timestamp 1704896540
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_318
timestamp 1704896540
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_319
timestamp 1704896540
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_320
timestamp 1704896540
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_321
timestamp 1704896540
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_322
timestamp 1704896540
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_323
timestamp 1704896540
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_324
timestamp 1704896540
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_325
timestamp 1704896540
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_326
timestamp 1704896540
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_327
timestamp 1704896540
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_328
timestamp 1704896540
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_329
timestamp 1704896540
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_330
timestamp 1704896540
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_331
timestamp 1704896540
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_332
timestamp 1704896540
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_333
timestamp 1704896540
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_334
timestamp 1704896540
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_335
timestamp 1704896540
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_336
timestamp 1704896540
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_337
timestamp 1704896540
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_338
timestamp 1704896540
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_339
timestamp 1704896540
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_340
timestamp 1704896540
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_341
timestamp 1704896540
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_342
timestamp 1704896540
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_343
timestamp 1704896540
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_344
timestamp 1704896540
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_345
timestamp 1704896540
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_346
timestamp 1704896540
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_347
timestamp 1704896540
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_348
timestamp 1704896540
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_349
timestamp 1704896540
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_350
timestamp 1704896540
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_351
timestamp 1704896540
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_352
timestamp 1704896540
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_353
timestamp 1704896540
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_354
timestamp 1704896540
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_355
timestamp 1704896540
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_356
timestamp 1704896540
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_357
timestamp 1704896540
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_358
timestamp 1704896540
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_359
timestamp 1704896540
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_360
timestamp 1704896540
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_361
timestamp 1704896540
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_362
timestamp 1704896540
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_363
timestamp 1704896540
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_364
timestamp 1704896540
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_365
timestamp 1704896540
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_366
timestamp 1704896540
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_367
timestamp 1704896540
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_368
timestamp 1704896540
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_369
timestamp 1704896540
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_370
timestamp 1704896540
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_371
timestamp 1704896540
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_372
timestamp 1704896540
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_373
timestamp 1704896540
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_374
timestamp 1704896540
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_375
timestamp 1704896540
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_376
timestamp 1704896540
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_377
timestamp 1704896540
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_378
timestamp 1704896540
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_379
timestamp 1704896540
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_380
timestamp 1704896540
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_381
timestamp 1704896540
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_382
timestamp 1704896540
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_383
timestamp 1704896540
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_384
timestamp 1704896540
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_385
timestamp 1704896540
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_386
timestamp 1704896540
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_387
timestamp 1704896540
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_388
timestamp 1704896540
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_389
timestamp 1704896540
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_390
timestamp 1704896540
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_391
timestamp 1704896540
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_392
timestamp 1704896540
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_393
timestamp 1704896540
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_394
timestamp 1704896540
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_395
timestamp 1704896540
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_396
timestamp 1704896540
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_397
timestamp 1704896540
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_398
timestamp 1704896540
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_399
timestamp 1704896540
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_400
timestamp 1704896540
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_401
timestamp 1704896540
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_402
timestamp 1704896540
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_403
timestamp 1704896540
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_404
timestamp 1704896540
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_405
timestamp 1704896540
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_406
timestamp 1704896540
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_407
timestamp 1704896540
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_408
timestamp 1704896540
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_409
timestamp 1704896540
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_410
timestamp 1704896540
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_411
timestamp 1704896540
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_412
timestamp 1704896540
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_413
timestamp 1704896540
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_414
timestamp 1704896540
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_415
timestamp 1704896540
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_416
timestamp 1704896540
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_417
timestamp 1704896540
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_418
timestamp 1704896540
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_419
timestamp 1704896540
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_420
timestamp 1704896540
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_421
timestamp 1704896540
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_422
timestamp 1704896540
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_423
timestamp 1704896540
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_424
timestamp 1704896540
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_425
timestamp 1704896540
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_426
timestamp 1704896540
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_427
timestamp 1704896540
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_428
timestamp 1704896540
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_429
timestamp 1704896540
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_430
timestamp 1704896540
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_431
timestamp 1704896540
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_432
timestamp 1704896540
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_433
timestamp 1704896540
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_434
timestamp 1704896540
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_435
timestamp 1704896540
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_436
timestamp 1704896540
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_437
timestamp 1704896540
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_438
timestamp 1704896540
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_439
timestamp 1704896540
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_440
timestamp 1704896540
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_441
timestamp 1704896540
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_442
timestamp 1704896540
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_443
timestamp 1704896540
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_444
timestamp 1704896540
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_445
timestamp 1704896540
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_446
timestamp 1704896540
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_447
timestamp 1704896540
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_448
timestamp 1704896540
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_449
timestamp 1704896540
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_450
timestamp 1704896540
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_451
timestamp 1704896540
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_452
timestamp 1704896540
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_453
timestamp 1704896540
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_454
timestamp 1704896540
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_455
timestamp 1704896540
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_456
timestamp 1704896540
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_457
timestamp 1704896540
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_458
timestamp 1704896540
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_459
timestamp 1704896540
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_460
timestamp 1704896540
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_461
timestamp 1704896540
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_462
timestamp 1704896540
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_463
timestamp 1704896540
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_464
timestamp 1704896540
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_465
timestamp 1704896540
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_466
timestamp 1704896540
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_467
timestamp 1704896540
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_468
timestamp 1704896540
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_469
timestamp 1704896540
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_470
timestamp 1704896540
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_471
timestamp 1704896540
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_472
timestamp 1704896540
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_473
timestamp 1704896540
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_474
timestamp 1704896540
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_475
timestamp 1704896540
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_476
timestamp 1704896540
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_477
timestamp 1704896540
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_478
timestamp 1704896540
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_479
timestamp 1704896540
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_480
timestamp 1704896540
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_481
timestamp 1704896540
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_482
timestamp 1704896540
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_483
timestamp 1704896540
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_484
timestamp 1704896540
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_485
timestamp 1704896540
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_486
timestamp 1704896540
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_487
timestamp 1704896540
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_488
timestamp 1704896540
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_489
timestamp 1704896540
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_490
timestamp 1704896540
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_491
timestamp 1704896540
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_492
timestamp 1704896540
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_493
timestamp 1704896540
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_494
timestamp 1704896540
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_495
timestamp 1704896540
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_496
timestamp 1704896540
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_497
timestamp 1704896540
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_498
timestamp 1704896540
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_499
timestamp 1704896540
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_500
timestamp 1704896540
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_501
timestamp 1704896540
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_502
timestamp 1704896540
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_503
timestamp 1704896540
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_504
timestamp 1704896540
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_505
timestamp 1704896540
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_506
timestamp 1704896540
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_507
timestamp 1704896540
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_508
timestamp 1704896540
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_509
timestamp 1704896540
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_510
timestamp 1704896540
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_511
timestamp 1704896540
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_512
timestamp 1704896540
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_513
timestamp 1704896540
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_514
timestamp 1704896540
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_515
timestamp 1704896540
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_516
timestamp 1704896540
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_517
timestamp 1704896540
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_518
timestamp 1704896540
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_519
timestamp 1704896540
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_520
timestamp 1704896540
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_521
timestamp 1704896540
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_522
timestamp 1704896540
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_523
timestamp 1704896540
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_524
timestamp 1704896540
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_525
timestamp 1704896540
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_526
timestamp 1704896540
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_527
timestamp 1704896540
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_528
timestamp 1704896540
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_529
timestamp 1704896540
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_530
timestamp 1704896540
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_531
timestamp 1704896540
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_532
timestamp 1704896540
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_533
timestamp 1704896540
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_534
timestamp 1704896540
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_535
timestamp 1704896540
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_536
timestamp 1704896540
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_537
timestamp 1704896540
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_538
timestamp 1704896540
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_539
timestamp 1704896540
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_540
timestamp 1704896540
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_541
timestamp 1704896540
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_542
timestamp 1704896540
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_543
timestamp 1704896540
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_544
timestamp 1704896540
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_545
timestamp 1704896540
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_546
timestamp 1704896540
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_547
timestamp 1704896540
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_548
timestamp 1704896540
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_549
timestamp 1704896540
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_550
timestamp 1704896540
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_551
timestamp 1704896540
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_552
timestamp 1704896540
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_553
timestamp 1704896540
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_554
timestamp 1704896540
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_555
timestamp 1704896540
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_556
timestamp 1704896540
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_557
timestamp 1704896540
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_558
timestamp 1704896540
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_559
timestamp 1704896540
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_560
timestamp 1704896540
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_561
timestamp 1704896540
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_562
timestamp 1704896540
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_563
timestamp 1704896540
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_564
timestamp 1704896540
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_565
timestamp 1704896540
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_566
timestamp 1704896540
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_567
timestamp 1704896540
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_568
timestamp 1704896540
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_569
timestamp 1704896540
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_570
timestamp 1704896540
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_571
timestamp 1704896540
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_572
timestamp 1704896540
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_573
timestamp 1704896540
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_574
timestamp 1704896540
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_575
timestamp 1704896540
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_576
timestamp 1704896540
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_577
timestamp 1704896540
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_578
timestamp 1704896540
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_579
timestamp 1704896540
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_580
timestamp 1704896540
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_581
timestamp 1704896540
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_582
timestamp 1704896540
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_583
timestamp 1704896540
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_584
timestamp 1704896540
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_585
timestamp 1704896540
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_586
timestamp 1704896540
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_587
timestamp 1704896540
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_588
timestamp 1704896540
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_589
timestamp 1704896540
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_590
timestamp 1704896540
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_591
timestamp 1704896540
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_592
timestamp 1704896540
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_593
timestamp 1704896540
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_594
timestamp 1704896540
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_595
timestamp 1704896540
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_596
timestamp 1704896540
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_597
timestamp 1704896540
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_598
timestamp 1704896540
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_599
timestamp 1704896540
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_600
timestamp 1704896540
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_601
timestamp 1704896540
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_602
timestamp 1704896540
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_603
timestamp 1704896540
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_604
timestamp 1704896540
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_605
timestamp 1704896540
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_606
timestamp 1704896540
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_607
timestamp 1704896540
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_608
timestamp 1704896540
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_609
timestamp 1704896540
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_610
timestamp 1704896540
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_611
timestamp 1704896540
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_612
timestamp 1704896540
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_613
timestamp 1704896540
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_614
timestamp 1704896540
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_615
timestamp 1704896540
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_616
timestamp 1704896540
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_617
timestamp 1704896540
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_618
timestamp 1704896540
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_619
timestamp 1704896540
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_620
timestamp 1704896540
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_621
timestamp 1704896540
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_622
timestamp 1704896540
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_623
timestamp 1704896540
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_624
timestamp 1704896540
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_625
timestamp 1704896540
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_626
timestamp 1704896540
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_627
timestamp 1704896540
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_628
timestamp 1704896540
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_629
timestamp 1704896540
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_630
timestamp 1704896540
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_631
timestamp 1704896540
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_632
timestamp 1704896540
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_633
timestamp 1704896540
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_634
timestamp 1704896540
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_635
timestamp 1704896540
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_636
timestamp 1704896540
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_637
timestamp 1704896540
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_638
timestamp 1704896540
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_639
timestamp 1704896540
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_640
timestamp 1704896540
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_641
timestamp 1704896540
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_642
timestamp 1704896540
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_643
timestamp 1704896540
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_644
timestamp 1704896540
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_645
timestamp 1704896540
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_646
timestamp 1704896540
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_647
timestamp 1704896540
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_648
timestamp 1704896540
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_649
timestamp 1704896540
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_650
timestamp 1704896540
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_651
timestamp 1704896540
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_652
timestamp 1704896540
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_653
timestamp 1704896540
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_654
timestamp 1704896540
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_655
timestamp 1704896540
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_656
timestamp 1704896540
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_657
timestamp 1704896540
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_658
timestamp 1704896540
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_659
timestamp 1704896540
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_660
timestamp 1704896540
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_661
timestamp 1704896540
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_662
timestamp 1704896540
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_663
timestamp 1704896540
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_664
timestamp 1704896540
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_665
timestamp 1704896540
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_666
timestamp 1704896540
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_667
timestamp 1704896540
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_668
timestamp 1704896540
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_669
timestamp 1704896540
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_670
timestamp 1704896540
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_671
timestamp 1704896540
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_672
timestamp 1704896540
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_673
timestamp 1704896540
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_674
timestamp 1704896540
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_675
timestamp 1704896540
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_676
timestamp 1704896540
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_677
timestamp 1704896540
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_678
timestamp 1704896540
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_679
timestamp 1704896540
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_680
timestamp 1704896540
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_681
timestamp 1704896540
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_682
timestamp 1704896540
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_683
timestamp 1704896540
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_684
timestamp 1704896540
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_685
timestamp 1704896540
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_686
timestamp 1704896540
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_687
timestamp 1704896540
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_688
timestamp 1704896540
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_689
timestamp 1704896540
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_690
timestamp 1704896540
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_691
timestamp 1704896540
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_692
timestamp 1704896540
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_693
timestamp 1704896540
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_694
timestamp 1704896540
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_695
timestamp 1704896540
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_696
timestamp 1704896540
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_697
timestamp 1704896540
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_698
timestamp 1704896540
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_699
timestamp 1704896540
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_700
timestamp 1704896540
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_701
timestamp 1704896540
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_702
timestamp 1704896540
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_703
timestamp 1704896540
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_704
timestamp 1704896540
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_705
timestamp 1704896540
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_706
timestamp 1704896540
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_707
timestamp 1704896540
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_708
timestamp 1704896540
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_709
timestamp 1704896540
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_710
timestamp 1704896540
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_711
timestamp 1704896540
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_712
timestamp 1704896540
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_713
timestamp 1704896540
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_714
timestamp 1704896540
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_715
timestamp 1704896540
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_716
timestamp 1704896540
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_717
timestamp 1704896540
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_718
timestamp 1704896540
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_719
timestamp 1704896540
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_720
timestamp 1704896540
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_721
timestamp 1704896540
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_722
timestamp 1704896540
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_723
timestamp 1704896540
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_724
timestamp 1704896540
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_725
timestamp 1704896540
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_726
timestamp 1704896540
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_727
timestamp 1704896540
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_728
timestamp 1704896540
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_729
timestamp 1704896540
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_730
timestamp 1704896540
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_731
timestamp 1704896540
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_732
timestamp 1704896540
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_733
timestamp 1704896540
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_734
timestamp 1704896540
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_735
timestamp 1704896540
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_736
timestamp 1704896540
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_737
timestamp 1704896540
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_738
timestamp 1704896540
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_739
timestamp 1704896540
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_740
timestamp 1704896540
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_741
timestamp 1704896540
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_742
timestamp 1704896540
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_743
timestamp 1704896540
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_744
timestamp 1704896540
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_745
timestamp 1704896540
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_746
timestamp 1704896540
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_747
timestamp 1704896540
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_748
timestamp 1704896540
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_749
timestamp 1704896540
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_750
timestamp 1704896540
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_751
timestamp 1704896540
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_752
timestamp 1704896540
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_753
timestamp 1704896540
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_754
timestamp 1704896540
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_755
timestamp 1704896540
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_756
timestamp 1704896540
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_757
timestamp 1704896540
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_758
timestamp 1704896540
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_759
timestamp 1704896540
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_760
timestamp 1704896540
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_761
timestamp 1704896540
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_762
timestamp 1704896540
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_763
timestamp 1704896540
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_764
timestamp 1704896540
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_765
timestamp 1704896540
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_766
timestamp 1704896540
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_767
timestamp 1704896540
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_768
timestamp 1704896540
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_769
timestamp 1704896540
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_770
timestamp 1704896540
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_771
timestamp 1704896540
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_772
timestamp 1704896540
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_773
timestamp 1704896540
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_774
timestamp 1704896540
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_775
timestamp 1704896540
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_776
timestamp 1704896540
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_777
timestamp 1704896540
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_778
timestamp 1704896540
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_779
timestamp 1704896540
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_780
timestamp 1704896540
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_781
timestamp 1704896540
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_782
timestamp 1704896540
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_783
timestamp 1704896540
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_784
timestamp 1704896540
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_785
timestamp 1704896540
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_786
timestamp 1704896540
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_787
timestamp 1704896540
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_788
timestamp 1704896540
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_789
timestamp 1704896540
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_790
timestamp 1704896540
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_791
timestamp 1704896540
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_792
timestamp 1704896540
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_793
timestamp 1704896540
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_794
timestamp 1704896540
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_795
timestamp 1704896540
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_796
timestamp 1704896540
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_797
timestamp 1704896540
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_798
timestamp 1704896540
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_799
timestamp 1704896540
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_800
timestamp 1704896540
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_801
timestamp 1704896540
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_802
timestamp 1704896540
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_803
timestamp 1704896540
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_804
timestamp 1704896540
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_805
timestamp 1704896540
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_806
timestamp 1704896540
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_807
timestamp 1704896540
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_808
timestamp 1704896540
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_809
timestamp 1704896540
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_810
timestamp 1704896540
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_811
timestamp 1704896540
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_812
timestamp 1704896540
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_813
timestamp 1704896540
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_814
timestamp 1704896540
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_815
timestamp 1704896540
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_816
timestamp 1704896540
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_817
timestamp 1704896540
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_818
timestamp 1704896540
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_819
timestamp 1704896540
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_820
timestamp 1704896540
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_821
timestamp 1704896540
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_822
timestamp 1704896540
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_823
timestamp 1704896540
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_824
timestamp 1704896540
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_825
timestamp 1704896540
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_826
timestamp 1704896540
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_827
timestamp 1704896540
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_828
timestamp 1704896540
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_829
timestamp 1704896540
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_830
timestamp 1704896540
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_831
timestamp 1704896540
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_832
timestamp 1704896540
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_833
timestamp 1704896540
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_834
timestamp 1704896540
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_835
timestamp 1704896540
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_836
timestamp 1704896540
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_837
timestamp 1704896540
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_838
timestamp 1704896540
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_839
timestamp 1704896540
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_840
timestamp 1704896540
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_841
timestamp 1704896540
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_842
timestamp 1704896540
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_843
timestamp 1704896540
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_844
timestamp 1704896540
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_845
timestamp 1704896540
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_846
timestamp 1704896540
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_847
timestamp 1704896540
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_848
timestamp 1704896540
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_849
timestamp 1704896540
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_850
timestamp 1704896540
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_851
timestamp 1704896540
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_852
timestamp 1704896540
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_853
timestamp 1704896540
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_854
timestamp 1704896540
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_855
timestamp 1704896540
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_856
timestamp 1704896540
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_857
timestamp 1704896540
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_858
timestamp 1704896540
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_859
timestamp 1704896540
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_860
timestamp 1704896540
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_861
timestamp 1704896540
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_862
timestamp 1704896540
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_863
timestamp 1704896540
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_864
timestamp 1704896540
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_865
timestamp 1704896540
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_866
timestamp 1704896540
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_867
timestamp 1704896540
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_868
timestamp 1704896540
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_869
timestamp 1704896540
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_870
timestamp 1704896540
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_871
timestamp 1704896540
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_872
timestamp 1704896540
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_873
timestamp 1704896540
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_874
timestamp 1704896540
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_875
timestamp 1704896540
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_876
timestamp 1704896540
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_877
timestamp 1704896540
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_878
timestamp 1704896540
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_879
timestamp 1704896540
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_880
timestamp 1704896540
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_881
timestamp 1704896540
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_882
timestamp 1704896540
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_883
timestamp 1704896540
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_884
timestamp 1704896540
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_885
timestamp 1704896540
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_886
timestamp 1704896540
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_887
timestamp 1704896540
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_888
timestamp 1704896540
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_889
timestamp 1704896540
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_890
timestamp 1704896540
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_891
timestamp 1704896540
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_892
timestamp 1704896540
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_893
timestamp 1704896540
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_894
timestamp 1704896540
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_895
timestamp 1704896540
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_896
timestamp 1704896540
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_897
timestamp 1704896540
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_898
timestamp 1704896540
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_899
timestamp 1704896540
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_900
timestamp 1704896540
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_901
timestamp 1704896540
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_902
timestamp 1704896540
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_903
timestamp 1704896540
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_904
timestamp 1704896540
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_905
timestamp 1704896540
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_906
timestamp 1704896540
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_907
timestamp 1704896540
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_908
timestamp 1704896540
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_909
timestamp 1704896540
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_910
timestamp 1704896540
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_911
timestamp 1704896540
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_912
timestamp 1704896540
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_913
timestamp 1704896540
transform 1 0 32016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_914
timestamp 1704896540
transform 1 0 37168 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_915
timestamp 1704896540
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_916
timestamp 1704896540
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_917
timestamp 1704896540
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_918
timestamp 1704896540
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_919
timestamp 1704896540
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_920
timestamp 1704896540
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_921
timestamp 1704896540
transform 1 0 34592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_922
timestamp 1704896540
transform 1 0 39744 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_923
timestamp 1704896540
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_924
timestamp 1704896540
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_925
timestamp 1704896540
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_926
timestamp 1704896540
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_927
timestamp 1704896540
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_928
timestamp 1704896540
transform 1 0 32016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_929
timestamp 1704896540
transform 1 0 37168 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_930
timestamp 1704896540
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_931
timestamp 1704896540
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_932
timestamp 1704896540
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_933
timestamp 1704896540
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_934
timestamp 1704896540
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_935
timestamp 1704896540
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_936
timestamp 1704896540
transform 1 0 34592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_937
timestamp 1704896540
transform 1 0 39744 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_938
timestamp 1704896540
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_939
timestamp 1704896540
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_940
timestamp 1704896540
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_941
timestamp 1704896540
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_942
timestamp 1704896540
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_943
timestamp 1704896540
transform 1 0 32016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_944
timestamp 1704896540
transform 1 0 37168 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_945
timestamp 1704896540
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_946
timestamp 1704896540
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_947
timestamp 1704896540
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_948
timestamp 1704896540
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_949
timestamp 1704896540
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_950
timestamp 1704896540
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_951
timestamp 1704896540
transform 1 0 34592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_952
timestamp 1704896540
transform 1 0 39744 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_953
timestamp 1704896540
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_954
timestamp 1704896540
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_955
timestamp 1704896540
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_956
timestamp 1704896540
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_957
timestamp 1704896540
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_958
timestamp 1704896540
transform 1 0 32016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_959
timestamp 1704896540
transform 1 0 37168 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_960
timestamp 1704896540
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_961
timestamp 1704896540
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_962
timestamp 1704896540
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_963
timestamp 1704896540
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_964
timestamp 1704896540
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_965
timestamp 1704896540
transform 1 0 29440 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_966
timestamp 1704896540
transform 1 0 34592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_967
timestamp 1704896540
transform 1 0 39744 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_968
timestamp 1704896540
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_969
timestamp 1704896540
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_970
timestamp 1704896540
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_971
timestamp 1704896540
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_972
timestamp 1704896540
transform 1 0 26864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_973
timestamp 1704896540
transform 1 0 32016 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_974
timestamp 1704896540
transform 1 0 37168 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_975
timestamp 1704896540
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_976
timestamp 1704896540
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_977
timestamp 1704896540
transform 1 0 13984 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_978
timestamp 1704896540
transform 1 0 19136 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_979
timestamp 1704896540
transform 1 0 24288 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_980
timestamp 1704896540
transform 1 0 29440 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_981
timestamp 1704896540
transform 1 0 34592 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_982
timestamp 1704896540
transform 1 0 39744 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_983
timestamp 1704896540
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_984
timestamp 1704896540
transform 1 0 11408 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_985
timestamp 1704896540
transform 1 0 16560 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_986
timestamp 1704896540
transform 1 0 21712 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_987
timestamp 1704896540
transform 1 0 26864 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_988
timestamp 1704896540
transform 1 0 32016 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_989
timestamp 1704896540
transform 1 0 37168 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_990
timestamp 1704896540
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_991
timestamp 1704896540
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_992
timestamp 1704896540
transform 1 0 13984 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_993
timestamp 1704896540
transform 1 0 19136 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_994
timestamp 1704896540
transform 1 0 24288 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_995
timestamp 1704896540
transform 1 0 29440 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_996
timestamp 1704896540
transform 1 0 34592 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_997
timestamp 1704896540
transform 1 0 39744 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_998
timestamp 1704896540
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_999
timestamp 1704896540
transform 1 0 11408 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1000
timestamp 1704896540
transform 1 0 16560 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1001
timestamp 1704896540
transform 1 0 21712 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1002
timestamp 1704896540
transform 1 0 26864 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1003
timestamp 1704896540
transform 1 0 32016 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1004
timestamp 1704896540
transform 1 0 37168 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1005
timestamp 1704896540
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1006
timestamp 1704896540
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1007
timestamp 1704896540
transform 1 0 13984 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1008
timestamp 1704896540
transform 1 0 19136 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1009
timestamp 1704896540
transform 1 0 24288 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1010
timestamp 1704896540
transform 1 0 29440 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1011
timestamp 1704896540
transform 1 0 34592 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1012
timestamp 1704896540
transform 1 0 39744 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1013
timestamp 1704896540
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1014
timestamp 1704896540
transform 1 0 11408 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1015
timestamp 1704896540
transform 1 0 16560 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1016
timestamp 1704896540
transform 1 0 21712 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1017
timestamp 1704896540
transform 1 0 26864 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1018
timestamp 1704896540
transform 1 0 32016 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1019
timestamp 1704896540
transform 1 0 37168 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_1020
timestamp 1704896540
transform 1 0 3680 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_1021
timestamp 1704896540
transform 1 0 8832 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_1022
timestamp 1704896540
transform 1 0 13984 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_1023
timestamp 1704896540
transform 1 0 19136 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_1024
timestamp 1704896540
transform 1 0 24288 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_1025
timestamp 1704896540
transform 1 0 29440 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_1026
timestamp 1704896540
transform 1 0 34592 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_1027
timestamp 1704896540
transform 1 0 39744 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_103_1028
timestamp 1704896540
transform 1 0 6256 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_103_1029
timestamp 1704896540
transform 1 0 11408 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_103_1030
timestamp 1704896540
transform 1 0 16560 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_103_1031
timestamp 1704896540
transform 1 0 21712 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_103_1032
timestamp 1704896540
transform 1 0 26864 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_103_1033
timestamp 1704896540
transform 1 0 32016 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_103_1034
timestamp 1704896540
transform 1 0 37168 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_1035
timestamp 1704896540
transform 1 0 3680 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_1036
timestamp 1704896540
transform 1 0 8832 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_1037
timestamp 1704896540
transform 1 0 13984 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_1038
timestamp 1704896540
transform 1 0 19136 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_1039
timestamp 1704896540
transform 1 0 24288 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_1040
timestamp 1704896540
transform 1 0 29440 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_1041
timestamp 1704896540
transform 1 0 34592 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_1042
timestamp 1704896540
transform 1 0 39744 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_105_1043
timestamp 1704896540
transform 1 0 6256 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_105_1044
timestamp 1704896540
transform 1 0 11408 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_105_1045
timestamp 1704896540
transform 1 0 16560 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_105_1046
timestamp 1704896540
transform 1 0 21712 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_105_1047
timestamp 1704896540
transform 1 0 26864 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_105_1048
timestamp 1704896540
transform 1 0 32016 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_105_1049
timestamp 1704896540
transform 1 0 37168 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_1050
timestamp 1704896540
transform 1 0 3680 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_1051
timestamp 1704896540
transform 1 0 8832 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_1052
timestamp 1704896540
transform 1 0 13984 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_1053
timestamp 1704896540
transform 1 0 19136 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_1054
timestamp 1704896540
transform 1 0 24288 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_1055
timestamp 1704896540
transform 1 0 29440 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_1056
timestamp 1704896540
transform 1 0 34592 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_1057
timestamp 1704896540
transform 1 0 39744 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_1058
timestamp 1704896540
transform 1 0 6256 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_1059
timestamp 1704896540
transform 1 0 11408 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_1060
timestamp 1704896540
transform 1 0 16560 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_1061
timestamp 1704896540
transform 1 0 21712 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_1062
timestamp 1704896540
transform 1 0 26864 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_1063
timestamp 1704896540
transform 1 0 32016 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_1064
timestamp 1704896540
transform 1 0 37168 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_1065
timestamp 1704896540
transform 1 0 3680 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_1066
timestamp 1704896540
transform 1 0 8832 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_1067
timestamp 1704896540
transform 1 0 13984 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_1068
timestamp 1704896540
transform 1 0 19136 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_1069
timestamp 1704896540
transform 1 0 24288 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_1070
timestamp 1704896540
transform 1 0 29440 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_1071
timestamp 1704896540
transform 1 0 34592 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_1072
timestamp 1704896540
transform 1 0 39744 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_1073
timestamp 1704896540
transform 1 0 6256 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_1074
timestamp 1704896540
transform 1 0 11408 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_1075
timestamp 1704896540
transform 1 0 16560 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_1076
timestamp 1704896540
transform 1 0 21712 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_1077
timestamp 1704896540
transform 1 0 26864 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_1078
timestamp 1704896540
transform 1 0 32016 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_1079
timestamp 1704896540
transform 1 0 37168 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_1080
timestamp 1704896540
transform 1 0 3680 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_1081
timestamp 1704896540
transform 1 0 8832 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_1082
timestamp 1704896540
transform 1 0 13984 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_1083
timestamp 1704896540
transform 1 0 19136 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_1084
timestamp 1704896540
transform 1 0 24288 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_1085
timestamp 1704896540
transform 1 0 29440 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_1086
timestamp 1704896540
transform 1 0 34592 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_1087
timestamp 1704896540
transform 1 0 39744 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_1088
timestamp 1704896540
transform 1 0 6256 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_1089
timestamp 1704896540
transform 1 0 11408 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_1090
timestamp 1704896540
transform 1 0 16560 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_1091
timestamp 1704896540
transform 1 0 21712 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_1092
timestamp 1704896540
transform 1 0 26864 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_1093
timestamp 1704896540
transform 1 0 32016 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_1094
timestamp 1704896540
transform 1 0 37168 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_1095
timestamp 1704896540
transform 1 0 3680 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_1096
timestamp 1704896540
transform 1 0 8832 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_1097
timestamp 1704896540
transform 1 0 13984 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_1098
timestamp 1704896540
transform 1 0 19136 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_1099
timestamp 1704896540
transform 1 0 24288 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_1100
timestamp 1704896540
transform 1 0 29440 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_1101
timestamp 1704896540
transform 1 0 34592 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_1102
timestamp 1704896540
transform 1 0 39744 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_1103
timestamp 1704896540
transform 1 0 6256 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_1104
timestamp 1704896540
transform 1 0 11408 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_1105
timestamp 1704896540
transform 1 0 16560 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_1106
timestamp 1704896540
transform 1 0 21712 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_1107
timestamp 1704896540
transform 1 0 26864 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_1108
timestamp 1704896540
transform 1 0 32016 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_1109
timestamp 1704896540
transform 1 0 37168 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_1110
timestamp 1704896540
transform 1 0 3680 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_1111
timestamp 1704896540
transform 1 0 8832 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_1112
timestamp 1704896540
transform 1 0 13984 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_1113
timestamp 1704896540
transform 1 0 19136 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_1114
timestamp 1704896540
transform 1 0 24288 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_1115
timestamp 1704896540
transform 1 0 29440 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_1116
timestamp 1704896540
transform 1 0 34592 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_1117
timestamp 1704896540
transform 1 0 39744 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_1118
timestamp 1704896540
transform 1 0 6256 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_1119
timestamp 1704896540
transform 1 0 11408 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_1120
timestamp 1704896540
transform 1 0 16560 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_1121
timestamp 1704896540
transform 1 0 21712 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_1122
timestamp 1704896540
transform 1 0 26864 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_1123
timestamp 1704896540
transform 1 0 32016 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_1124
timestamp 1704896540
transform 1 0 37168 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_1125
timestamp 1704896540
transform 1 0 3680 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_1126
timestamp 1704896540
transform 1 0 8832 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_1127
timestamp 1704896540
transform 1 0 13984 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_1128
timestamp 1704896540
transform 1 0 19136 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_1129
timestamp 1704896540
transform 1 0 24288 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_1130
timestamp 1704896540
transform 1 0 29440 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_1131
timestamp 1704896540
transform 1 0 34592 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_1132
timestamp 1704896540
transform 1 0 39744 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1133
timestamp 1704896540
transform 1 0 6256 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1134
timestamp 1704896540
transform 1 0 11408 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1135
timestamp 1704896540
transform 1 0 16560 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1136
timestamp 1704896540
transform 1 0 21712 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1137
timestamp 1704896540
transform 1 0 26864 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1138
timestamp 1704896540
transform 1 0 32016 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1139
timestamp 1704896540
transform 1 0 37168 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1140
timestamp 1704896540
transform 1 0 3680 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1141
timestamp 1704896540
transform 1 0 8832 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1142
timestamp 1704896540
transform 1 0 13984 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1143
timestamp 1704896540
transform 1 0 19136 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1144
timestamp 1704896540
transform 1 0 24288 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1145
timestamp 1704896540
transform 1 0 29440 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1146
timestamp 1704896540
transform 1 0 34592 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1147
timestamp 1704896540
transform 1 0 39744 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1148
timestamp 1704896540
transform 1 0 6256 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1149
timestamp 1704896540
transform 1 0 11408 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1150
timestamp 1704896540
transform 1 0 16560 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1151
timestamp 1704896540
transform 1 0 21712 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1152
timestamp 1704896540
transform 1 0 26864 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1153
timestamp 1704896540
transform 1 0 32016 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1154
timestamp 1704896540
transform 1 0 37168 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1155
timestamp 1704896540
transform 1 0 3680 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1156
timestamp 1704896540
transform 1 0 8832 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1157
timestamp 1704896540
transform 1 0 13984 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1158
timestamp 1704896540
transform 1 0 19136 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1159
timestamp 1704896540
transform 1 0 24288 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1160
timestamp 1704896540
transform 1 0 29440 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1161
timestamp 1704896540
transform 1 0 34592 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1162
timestamp 1704896540
transform 1 0 39744 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1163
timestamp 1704896540
transform 1 0 6256 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1164
timestamp 1704896540
transform 1 0 11408 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1165
timestamp 1704896540
transform 1 0 16560 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1166
timestamp 1704896540
transform 1 0 21712 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1167
timestamp 1704896540
transform 1 0 26864 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1168
timestamp 1704896540
transform 1 0 32016 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1169
timestamp 1704896540
transform 1 0 37168 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1170
timestamp 1704896540
transform 1 0 3680 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1171
timestamp 1704896540
transform 1 0 8832 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1172
timestamp 1704896540
transform 1 0 13984 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1173
timestamp 1704896540
transform 1 0 19136 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1174
timestamp 1704896540
transform 1 0 24288 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1175
timestamp 1704896540
transform 1 0 29440 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1176
timestamp 1704896540
transform 1 0 34592 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1177
timestamp 1704896540
transform 1 0 39744 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1178
timestamp 1704896540
transform 1 0 3680 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1179
timestamp 1704896540
transform 1 0 6256 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1180
timestamp 1704896540
transform 1 0 8832 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1181
timestamp 1704896540
transform 1 0 11408 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1182
timestamp 1704896540
transform 1 0 13984 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1183
timestamp 1704896540
transform 1 0 16560 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1184
timestamp 1704896540
transform 1 0 19136 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1185
timestamp 1704896540
transform 1 0 21712 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1186
timestamp 1704896540
transform 1 0 24288 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1187
timestamp 1704896540
transform 1 0 26864 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1188
timestamp 1704896540
transform 1 0 29440 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1189
timestamp 1704896540
transform 1 0 32016 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1190
timestamp 1704896540
transform 1 0 34592 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1191
timestamp 1704896540
transform 1 0 37168 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1192
timestamp 1704896540
transform 1 0 39744 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  ZeroToFiveCounter_9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 2944 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ZeroToFiveCounter_10
timestamp 1704896540
transform 1 0 39836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ZeroToFiveCounter_11
timestamp 1704896540
transform 1 0 34132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ZeroToFiveCounter_12
timestamp 1704896540
transform 1 0 28888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ZeroToFiveCounter_13
timestamp 1704896540
transform 1 0 23644 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ZeroToFiveCounter_14
timestamp 1704896540
transform 1 0 18400 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ZeroToFiveCounter_15
timestamp 1704896540
transform 1 0 13156 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ZeroToFiveCounter_16
timestamp 1704896540
transform 1 0 7912 0 1 2176
box -38 -48 314 592
<< labels >>
flabel metal4 s 2604 2128 2924 69680 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 7604 2128 7924 69680 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 12604 2128 12924 69680 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17604 2128 17924 69680 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 22604 2128 22924 69680 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 27604 2128 27924 69680 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 32604 2128 32924 69680 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 37604 2128 37924 69680 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 3676 40896 3996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 8676 40896 8996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 13676 40896 13996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 18676 40896 18996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 23676 40896 23996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 28676 40896 28996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 33676 40896 33996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 38676 40896 38996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 43676 40896 43996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 48676 40896 48996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 53676 40896 53996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 58676 40896 58996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 63676 40896 63996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 68676 40896 68996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 1944 2128 2264 69680 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 6944 2128 7264 69680 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 11944 2128 12264 69680 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 16944 2128 17264 69680 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 21944 2128 22264 69680 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 26944 2128 27264 69680 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 31944 2128 32264 69680 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 36944 2128 37264 69680 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 3016 40896 3336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 8016 40896 8336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 13016 40896 13336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 18016 40896 18336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 23016 40896 23336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 28016 40896 28336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 33016 40896 33336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 38016 40896 38336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 43016 40896 43336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 48016 40896 48336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 53016 40896 53336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 58016 40896 58336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 63016 40896 63336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 68016 40896 68336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 39302 0 39358 800 0 FreeSans 224 90 0 0 an[0]
port 2 nsew signal output
flabel metal2 s 34058 0 34114 800 0 FreeSans 224 90 0 0 an[1]
port 3 nsew signal output
flabel metal2 s 28814 0 28870 800 0 FreeSans 224 90 0 0 an[2]
port 4 nsew signal output
flabel metal2 s 23570 0 23626 800 0 FreeSans 224 90 0 0 an[3]
port 5 nsew signal output
flabel metal2 s 18326 0 18382 800 0 FreeSans 224 90 0 0 an[4]
port 6 nsew signal output
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 an[5]
port 7 nsew signal output
flabel metal2 s 7838 0 7894 800 0 FreeSans 224 90 0 0 an[6]
port 8 nsew signal output
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 an[7]
port 9 nsew signal output
flabel metal3 s 0 35912 800 36032 0 FreeSans 480 0 0 0 clk
port 10 nsew signal input
flabel metal3 s 41200 35912 42000 36032 0 FreeSans 480 0 0 0 rst
port 11 nsew signal input
flabel metal2 s 38842 71200 38898 72000 0 FreeSans 224 90 0 0 seg[0]
port 12 nsew signal output
flabel metal2 s 32862 71200 32918 72000 0 FreeSans 224 90 0 0 seg[1]
port 13 nsew signal output
flabel metal2 s 26882 71200 26938 72000 0 FreeSans 224 90 0 0 seg[2]
port 14 nsew signal output
flabel metal2 s 20902 71200 20958 72000 0 FreeSans 224 90 0 0 seg[3]
port 15 nsew signal output
flabel metal2 s 14922 71200 14978 72000 0 FreeSans 224 90 0 0 seg[4]
port 16 nsew signal output
flabel metal2 s 8942 71200 8998 72000 0 FreeSans 224 90 0 0 seg[5]
port 17 nsew signal output
flabel metal2 s 2962 71200 3018 72000 0 FreeSans 224 90 0 0 seg[6]
port 18 nsew signal output
rlabel metal1 20976 69632 20976 69632 0 VGND
rlabel metal1 20976 69088 20976 69088 0 VPWR
rlabel metal1 28934 25194 28934 25194 0 _000_
rlabel metal1 37950 32334 37950 32334 0 _001_
rlabel metal2 3266 22882 3266 22882 0 _002_
rlabel metal1 14168 10506 14168 10506 0 _003_
rlabel metal1 22632 9146 22632 9146 0 _004_
rlabel metal1 31648 10506 31648 10506 0 _005_
rlabel metal1 4508 29070 4508 29070 0 _006_
rlabel metal2 6624 35880 6624 35880 0 _007_
rlabel metal2 5014 52938 5014 52938 0 _008_
rlabel metal1 18354 63750 18354 63750 0 _009_
rlabel metal1 21252 48518 21252 48518 0 _010_
rlabel metal1 28796 33286 28796 33286 0 _011_
rlabel metal2 1886 33082 1886 33082 0 _012_
rlabel metal1 32154 21386 32154 21386 0 _013_
rlabel metal1 23414 24718 23414 24718 0 _014_
rlabel metal2 22218 39202 22218 39202 0 _015_
rlabel metal1 8970 36686 8970 36686 0 _016_
rlabel metal2 3634 18496 3634 18496 0 _017_
rlabel metal1 36110 53448 36110 53448 0 _018_
rlabel metal1 4416 56746 4416 56746 0 _019_
rlabel via2 7590 9605 7590 9605 0 _020_
rlabel metal2 13570 47668 13570 47668 0 _021_
rlabel metal2 31602 53346 31602 53346 0 _022_
rlabel metal1 14214 29580 14214 29580 0 _023_
rlabel metal1 7222 30362 7222 30362 0 _024_
rlabel metal2 13662 10880 13662 10880 0 _025_
rlabel metal1 37812 56270 37812 56270 0 _026_
rlabel metal1 7452 3026 7452 3026 0 _027_
rlabel metal1 15325 25262 15325 25262 0 _028_
rlabel metal2 6394 60384 6394 60384 0 _029_
rlabel metal2 7406 56007 7406 56007 0 _030_
rlabel metal1 18400 16966 18400 16966 0 _031_
rlabel metal1 36593 37638 36593 37638 0 _032_
rlabel metal1 29111 53550 29111 53550 0 _033_
rlabel metal1 13616 4998 13616 4998 0 _034_
rlabel metal1 9292 8058 9292 8058 0 _035_
rlabel metal1 7866 58854 7866 58854 0 _036_
rlabel metal1 38831 56406 38831 56406 0 _037_
rlabel metal2 38686 27676 38686 27676 0 _038_
rlabel metal1 27876 37162 27876 37162 0 _039_
rlabel metal1 27784 13498 27784 13498 0 _040_
rlabel metal1 32568 63750 32568 63750 0 _041_
rlabel metal1 4347 4522 4347 4522 0 _042_
rlabel metal1 9798 41446 9798 41446 0 _043_
rlabel metal1 30452 11254 30452 11254 0 _044_
rlabel metal2 3910 56313 3910 56313 0 _045_
rlabel metal1 20838 63750 20838 63750 0 _046_
rlabel metal1 14069 19822 14069 19822 0 _047_
rlabel metal1 19511 19414 19511 19414 0 _048_
rlabel metal1 35979 57426 35979 57426 0 _049_
rlabel metal2 24242 24616 24242 24616 0 _050_
rlabel metal1 24012 59942 24012 59942 0 _051_
rlabel metal1 9844 33626 9844 33626 0 _052_
rlabel metal1 10166 18598 10166 18598 0 _053_
rlabel metal1 36195 53550 36195 53550 0 _054_
rlabel metal2 18722 31144 18722 31144 0 _055_
rlabel metal1 3542 20570 3542 20570 0 _056_
rlabel metal1 19182 14042 19182 14042 0 _057_
rlabel metal2 19642 27302 19642 27302 0 _058_
rlabel metal1 2070 45349 2070 45349 0 _059_
rlabel metal1 4830 20366 4830 20366 0 _060_
rlabel metal2 8694 44302 8694 44302 0 _061_
rlabel metal2 2438 48042 2438 48042 0 _062_
rlabel metal1 17664 10574 17664 10574 0 _063_
rlabel metal1 39606 58480 39606 58480 0 _064_
rlabel metal1 20240 63274 20240 63274 0 _065_
rlabel metal2 34914 18768 34914 18768 0 _066_
rlabel metal2 40158 57732 40158 57732 0 _067_
rlabel metal1 15364 16558 15364 16558 0 _068_
rlabel metal2 20378 49436 20378 49436 0 _069_
rlabel metal1 18814 63478 18814 63478 0 _070_
rlabel metal2 17434 44336 17434 44336 0 _071_
rlabel metal1 39839 57766 39839 57766 0 _072_
rlabel metal1 14490 44166 14490 44166 0 _073_
rlabel metal1 7314 41140 7314 41140 0 _074_
rlabel metal1 25024 63546 25024 63546 0 _075_
rlabel metal1 18584 30226 18584 30226 0 _076_
rlabel metal2 2898 3706 2898 3706 0 _077_
rlabel metal1 18492 64294 18492 64294 0 _078_
rlabel metal1 32384 51850 32384 51850 0 _079_
rlabel metal1 34546 26010 34546 26010 0 _080_
rlabel metal1 32246 25738 32246 25738 0 _081_
rlabel metal1 7222 41072 7222 41072 0 _082_
rlabel metal1 2944 17238 2944 17238 0 _083_
rlabel metal1 11178 41038 11178 41038 0 _084_
rlabel metal1 21298 64362 21298 64362 0 _085_
rlabel metal1 4952 3570 4952 3570 0 _086_
rlabel metal1 35742 14858 35742 14858 0 _087_
rlabel metal2 33212 12852 33212 12852 0 _088_
rlabel metal1 32430 33490 32430 33490 0 _089_
rlabel metal1 33626 23800 33626 23800 0 _090_
rlabel metal1 33350 23766 33350 23766 0 _091_
rlabel metal1 2208 67694 2208 67694 0 _092_
rlabel metal1 22770 64940 22770 64940 0 _093_
rlabel metal1 27232 64294 27232 64294 0 _094_
rlabel metal1 5612 17238 5612 17238 0 _095_
rlabel metal1 38226 60282 38226 60282 0 _096_
rlabel metal1 37704 60010 37704 60010 0 _097_
rlabel metal1 38042 59942 38042 59942 0 _098_
rlabel metal1 13524 38794 13524 38794 0 _099_
rlabel metal1 25622 4760 25622 4760 0 _100_
rlabel metal2 4554 16864 4554 16864 0 _101_
rlabel metal1 2806 16966 2806 16966 0 _102_
rlabel metal1 10028 17034 10028 17034 0 _103_
rlabel metal1 2254 3468 2254 3468 0 _104_
rlabel via2 38962 14365 38962 14365 0 _105_
rlabel metal1 17434 29240 17434 29240 0 _106_
rlabel via2 18906 7837 18906 7837 0 _107_
rlabel metal2 12098 31756 12098 31756 0 _108_
rlabel metal1 19872 17238 19872 17238 0 _109_
rlabel metal1 28750 55590 28750 55590 0 _110_
rlabel metal1 25576 28186 25576 28186 0 _111_
rlabel metal1 29946 3026 29946 3026 0 _112_
rlabel metal2 19366 25568 19366 25568 0 _113_
rlabel metal1 2852 40494 2852 40494 0 _114_
rlabel metal2 29578 39338 29578 39338 0 _115_
rlabel metal2 33994 33728 33994 33728 0 _116_
rlabel metal1 5612 10642 5612 10642 0 _117_
rlabel metal2 9568 35880 9568 35880 0 _118_
rlabel metal1 3726 63342 3726 63342 0 _119_
rlabel metal1 16146 8942 16146 8942 0 _120_
rlabel metal1 23920 66130 23920 66130 0 _121_
rlabel metal1 4002 63546 4002 63546 0 _122_
rlabel metal1 24656 65994 24656 65994 0 _123_
rlabel metal1 36616 52462 36616 52462 0 _124_
rlabel metal1 29854 32470 29854 32470 0 _125_
rlabel metal1 22586 62118 22586 62118 0 _126_
rlabel metal1 3036 44914 3036 44914 0 _127_
rlabel metal1 39560 30906 39560 30906 0 _128_
rlabel metal2 18998 36958 18998 36958 0 _129_
rlabel metal2 6486 66164 6486 66164 0 _130_
rlabel metal1 9476 36346 9476 36346 0 _131_
rlabel metal1 18446 63920 18446 63920 0 _132_
rlabel metal2 18630 49980 18630 49980 0 _133_
rlabel metal1 2622 44778 2622 44778 0 _134_
rlabel metal2 6118 52666 6118 52666 0 _135_
rlabel metal2 18630 7344 18630 7344 0 _136_
rlabel metal2 4738 7616 4738 7616 0 _137_
rlabel metal1 18354 2822 18354 2822 0 _138_
rlabel metal1 36432 18054 36432 18054 0 _139_
rlabel metal1 36754 2618 36754 2618 0 _140_
rlabel metal2 1702 32538 1702 32538 0 _141_
rlabel metal1 37674 68646 37674 68646 0 _142_
rlabel metal1 32614 21379 32614 21379 0 _143_
rlabel metal1 28520 14790 28520 14790 0 _144_
rlabel metal2 8924 45540 8924 45540 0 _145_
rlabel metal1 23138 19822 23138 19822 0 _146_
rlabel metal1 19205 3026 19205 3026 0 _147_
rlabel metal2 8510 3366 8510 3366 0 _148_
rlabel metal2 30590 28713 30590 28713 0 _149_
rlabel metal2 20562 55454 20562 55454 0 _150_
rlabel metal2 34592 55200 34592 55200 0 _151_
rlabel metal1 21850 55046 21850 55046 0 _152_
rlabel metal1 3450 18768 3450 18768 0 _153_
rlabel metal2 16606 41242 16606 41242 0 _154_
rlabel metal2 36846 60010 36846 60010 0 _155_
rlabel metal1 39606 62254 39606 62254 0 _156_
rlabel metal1 39008 2346 39008 2346 0 _157_
rlabel metal2 6394 35428 6394 35428 0 _158_
rlabel metal1 20608 5202 20608 5202 0 _159_
rlabel metal1 1886 4624 1886 4624 0 _160_
rlabel metal2 24886 61472 24886 61472 0 _161_
rlabel metal3 1579 35972 1579 35972 0 clk
rlabel via2 24610 22661 24610 22661 0 clknet_0_clk
rlabel metal2 6670 19856 6670 19856 0 clknet_2_0__leaf_clk
rlabel metal1 25300 22406 25300 22406 0 clknet_2_1__leaf_clk
rlabel metal1 5658 56882 5658 56882 0 clknet_2_2__leaf_clk
rlabel metal2 37306 56814 37306 56814 0 clknet_2_3__leaf_clk
rlabel metal1 3220 20502 3220 20502 0 decoder.digit\[0\]
rlabel metal1 17342 54196 17342 54196 0 decoder.digit\[1\]
rlabel metal1 39054 58514 39054 58514 0 decoder.digit\[2\]
rlabel metal2 1426 45220 1426 45220 0 decoder.digit\[3\]
rlabel metal1 40296 29138 40296 29138 0 net1
rlabel metal2 39330 1588 39330 1588 0 net10
rlabel metal2 34086 1520 34086 1520 0 net11
rlabel metal2 28842 1520 28842 1520 0 net12
rlabel metal2 23598 1520 23598 1520 0 net13
rlabel metal2 18354 1520 18354 1520 0 net14
rlabel metal2 13110 1520 13110 1520 0 net15
rlabel metal2 7866 959 7866 959 0 net16
rlabel metal2 39146 50031 39146 50031 0 net2
rlabel metal1 28658 52598 28658 52598 0 net3
rlabel metal1 31188 24310 31188 24310 0 net4
rlabel metal2 21206 50116 21206 50116 0 net5
rlabel metal1 27324 2550 27324 2550 0 net6
rlabel metal1 7682 38386 7682 38386 0 net7
rlabel metal1 3312 69394 3312 69394 0 net8
rlabel metal2 2622 1027 2622 1027 0 net9
rlabel metal1 37812 8942 37812 8942 0 one_second_counter\[0\]
rlabel metal1 26082 27982 26082 27982 0 one_second_counter\[10\]
rlabel metal2 19642 56746 19642 56746 0 one_second_counter\[11\]
rlabel metal2 17480 31892 17480 31892 0 one_second_counter\[12\]
rlabel metal1 3082 40460 3082 40460 0 one_second_counter\[13\]
rlabel metal2 16606 64192 16606 64192 0 one_second_counter\[14\]
rlabel metal1 36754 68714 36754 68714 0 one_second_counter\[15\]
rlabel metal1 3174 44846 3174 44846 0 one_second_counter\[16\]
rlabel via1 5474 44795 5474 44795 0 one_second_counter\[17\]
rlabel metal1 4462 44914 4462 44914 0 one_second_counter\[18\]
rlabel metal1 4140 44982 4140 44982 0 one_second_counter\[19\]
rlabel metal1 23138 53006 23138 53006 0 one_second_counter\[1\]
rlabel metal2 3358 17442 3358 17442 0 one_second_counter\[20\]
rlabel metal1 4876 17170 4876 17170 0 one_second_counter\[21\]
rlabel metal1 4600 17102 4600 17102 0 one_second_counter\[22\]
rlabel metal1 3634 17272 3634 17272 0 one_second_counter\[23\]
rlabel metal1 8096 41106 8096 41106 0 one_second_counter\[24\]
rlabel metal1 17112 44166 17112 44166 0 one_second_counter\[25\]
rlabel metal1 17158 51374 17158 51374 0 one_second_counter\[26\]
rlabel metal1 11960 3366 11960 3366 0 one_second_counter\[2\]
rlabel metal1 20562 34034 20562 34034 0 one_second_counter\[3\]
rlabel metal1 24840 4522 24840 4522 0 one_second_counter\[4\]
rlabel metal2 22034 39236 22034 39236 0 one_second_counter\[5\]
rlabel metal1 5842 52326 5842 52326 0 one_second_counter\[6\]
rlabel metal1 5980 30566 5980 30566 0 one_second_counter\[7\]
rlabel metal1 18584 17306 18584 17306 0 one_second_counter\[8\]
rlabel metal2 18538 17408 18538 17408 0 one_second_counter\[9\]
rlabel metal1 39652 57902 39652 57902 0 one_second_enable
rlabel metal2 40526 36057 40526 36057 0 rst
rlabel metal2 38962 70431 38962 70431 0 seg[0]
rlabel metal2 32982 70431 32982 70431 0 seg[1]
rlabel metal2 27002 70431 27002 70431 0 seg[2]
rlabel metal2 21022 70431 21022 70431 0 seg[3]
rlabel metal2 15042 70431 15042 70431 0 seg[4]
rlabel metal1 9016 69530 9016 69530 0 seg[5]
rlabel metal2 3082 70431 3082 70431 0 seg[6]
<< properties >>
string FIXED_BBOX 0 0 42000 72000
<< end >>
